//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(KEYINPUT81), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G162gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n212), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n209), .B(new_n215), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n214), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(new_n225), .A3(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(G127gat), .A2(G134gat), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT72), .B(G127gat), .Z(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G113gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(G120gat), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(G113gat), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT73), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT74), .ZN(new_n245));
  NAND2_X1  g044(.A1(G127gat), .A2(G134gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G127gat), .A2(G134gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(G127gat), .A2(G134gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT74), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT1), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n244), .A2(new_n251), .A3(KEYINPUT75), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT75), .B1(new_n244), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n236), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT82), .B1(new_n228), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n244), .A2(new_n251), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT75), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n251), .A3(KEYINPUT75), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n235), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT82), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n260), .A2(new_n227), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n203), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n221), .A2(new_n222), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n236), .C1(new_n252), .C2(new_n253), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n259), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n236), .A4(new_n264), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT84), .B1(new_n263), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n203), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n228), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n261), .B1(new_n260), .B2(new_n227), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n271), .A4(new_n272), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n223), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n282), .A2(new_n265), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT5), .B1(new_n283), .B2(new_n203), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G1gat), .B(G29gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT0), .ZN(new_n288));
  XNOR2_X1  g087(.A(G57gat), .B(G85gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n269), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n278), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n290), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n284), .B1(new_n274), .B2(new_n280), .ZN(new_n296));
  INV_X1    g095(.A(new_n293), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G8gat), .B(G36gat), .Z(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT80), .ZN(new_n302));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT23), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n308), .B(KEYINPUT25), .C1(G176gat), .C2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT67), .B(KEYINPUT24), .ZN(new_n312));
  AND2_X1   g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT68), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT67), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n314), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n311), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n314), .A2(new_n322), .A3(KEYINPUT69), .A4(new_n325), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  AND2_X1   g129(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n310), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(KEYINPUT23), .B2(new_n306), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT66), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n310), .ZN(new_n337));
  INV_X1    g136(.A(new_n332), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n308), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n323), .A2(new_n343), .B1(new_n321), .B2(new_n315), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n324), .A2(G190gat), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n344), .B(new_n345), .C1(new_n343), .C2(new_n323), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n336), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(new_n313), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT71), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n306), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n348), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G226gat), .ZN(new_n362));
  INV_X1    g161(.A(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n313), .B1(new_n316), .B2(new_n318), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n325), .B1(new_n365), .B2(new_n320), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n312), .A2(KEYINPUT68), .A3(new_n313), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n327), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n311), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n329), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n330), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n361), .A2(new_n364), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  XNOR2_X1  g176(.A(G197gat), .B(G204gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT22), .ZN(new_n379));
  INV_X1    g178(.A(G211gat), .ZN(new_n380));
  INV_X1    g179(.A(G218gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n364), .A2(KEYINPUT29), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n348), .B2(new_n360), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n376), .A2(new_n377), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n376), .A2(new_n385), .A3(new_n387), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT79), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n360), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n364), .A3(new_n374), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n388), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT37), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n305), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n361), .A2(new_n375), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n386), .ZN(new_n401));
  INV_X1    g200(.A(new_n384), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n383), .B(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n376), .A2(new_n403), .A3(new_n387), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n405), .A2(KEYINPUT37), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT38), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT6), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n396), .A2(new_n305), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n300), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT38), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT79), .B(new_n389), .C1(new_n401), .C2(new_n385), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT37), .A3(new_n388), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT89), .B(new_n412), .C1(new_n398), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n397), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n304), .A3(new_n414), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(KEYINPUT38), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n411), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n304), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n413), .A2(new_n304), .A3(new_n388), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT30), .B1(new_n396), .B2(new_n305), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n422), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(KEYINPUT88), .A3(new_n425), .A4(new_n424), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n292), .B1(new_n255), .B2(new_n262), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n275), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n283), .A2(new_n203), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(KEYINPUT39), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n435), .A3(new_n275), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n290), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT40), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n434), .A2(KEYINPUT40), .A3(new_n290), .A4(new_n436), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n439), .A2(new_n298), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n428), .A2(new_n430), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT3), .B1(new_n403), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n445), .B2(new_n264), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n225), .B1(new_n385), .B2(KEYINPUT29), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n223), .ZN(new_n448));
  INV_X1    g247(.A(G228gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(new_n363), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n226), .A2(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n385), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n446), .A2(new_n448), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT86), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n452), .A2(new_n450), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n448), .A4(new_n446), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(new_n223), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n450), .B1(new_n459), .B2(new_n452), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(KEYINPUT87), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n458), .B2(new_n461), .ZN(new_n468));
  AOI211_X1 g267(.A(G22gat), .B(new_n460), .C1(new_n454), .C2(new_n457), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT31), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G50gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n466), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n467), .B(new_n473), .C1(new_n468), .C2(new_n469), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n442), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n420), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n260), .B1(new_n348), .B2(new_n360), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n372), .A2(new_n374), .A3(new_n254), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(new_n363), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n487), .A2(KEYINPUT34), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(KEYINPUT34), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT32), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT76), .A4(new_n485), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT33), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  XOR2_X1   g297(.A(G15gat), .B(G43gat), .Z(new_n499));
  XNOR2_X1  g298(.A(G71gat), .B(G99gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  AOI221_X4 g302(.A(new_n492), .B1(KEYINPUT33), .B2(new_n501), .C1(new_n495), .C2(new_n496), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n491), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n495), .A2(new_n496), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n497), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n504), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n490), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n480), .B1(new_n505), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT77), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n505), .A2(new_n514), .A3(new_n512), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT77), .B(new_n491), .C1(new_n503), .C2(new_n504), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n513), .B1(new_n517), .B2(new_n480), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n300), .A2(new_n409), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n426), .A2(new_n427), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n475), .A2(new_n476), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n479), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n477), .A2(new_n505), .A3(new_n512), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT35), .B1(new_n526), .B2(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n428), .A2(new_n430), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n517), .A3(new_n529), .A4(new_n519), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n202), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n531), .B(KEYINPUT90), .C1(new_n479), .C2(new_n524), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT12), .Z(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT14), .B(G29gat), .Z(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(G36gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546));
  XNOR2_X1  g345(.A(G43gat), .B(G50gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n545), .A2(new_n546), .B1(KEYINPUT15), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(KEYINPUT15), .B2(new_n547), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT17), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552));
  AOI21_X1  g351(.A(G1gat), .B1(new_n552), .B2(KEYINPUT93), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n552), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT16), .ZN(new_n555));
  AOI211_X1 g354(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n552), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT94), .B1(new_n552), .B2(G1gat), .ZN(new_n557));
  INV_X1    g356(.A(G8gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n556), .B(new_n559), .ZN(new_n560));
  MUX2_X1   g359(.A(new_n550), .B(new_n551), .S(new_n560), .Z(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n560), .B(new_n550), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n562), .B(KEYINPUT13), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n541), .B1(new_n567), .B2(KEYINPUT95), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT18), .B1(new_n561), .B2(new_n562), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n535), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n300), .A2(new_n409), .ZN(new_n574));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  NAND2_X1  g376(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(G85gat), .A3(G92gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT100), .ZN(new_n580));
  NOR2_X1   g379(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G99gat), .B(G106gat), .Z(new_n583));
  INV_X1    g382(.A(G99gat), .ZN(new_n584));
  INV_X1    g383(.A(G106gat), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT8), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT101), .B(G85gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(G92gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT102), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n582), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n583), .B1(new_n582), .B2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  OR2_X1    g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G78gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT96), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n594), .A2(new_n600), .B1(new_n598), .B2(new_n599), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n597), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT98), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n592), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT105), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n602), .B(KEYINPUT104), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  MUX2_X1   g408(.A(new_n607), .B(new_n609), .S(new_n592), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n604), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n610), .A2(new_n613), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n577), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n616), .A3(new_n577), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n592), .A2(new_n550), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n622));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n590), .A2(new_n591), .ZN(new_n624));
  OAI221_X1 g423(.A(new_n621), .B1(new_n622), .B2(new_n623), .C1(new_n551), .C2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT103), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G134gat), .B(G162gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n622), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n628), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n602), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT97), .Z(new_n637));
  XOR2_X1   g436(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n560), .B1(new_n603), .B2(new_n635), .ZN(new_n642));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n642), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n620), .A2(new_n634), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT106), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n573), .A2(new_n574), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n573), .A2(new_n653), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n528), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND4_X1  g458(.A1(new_n657), .A2(KEYINPUT42), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(KEYINPUT107), .A3(new_n658), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n656), .B2(new_n528), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(G8gat), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n659), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n661), .B2(new_n663), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n660), .B(new_n664), .C1(new_n666), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n656), .B2(new_n518), .ZN(new_n668));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n669), .A3(new_n517), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n572), .B2(new_n670), .ZN(G1326gat));
  OR3_X1    g470(.A1(new_n656), .A2(KEYINPUT108), .A3(new_n477), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT108), .B1(new_n656), .B2(new_n477), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1327gat));
  NOR2_X1   g478(.A1(new_n620), .A2(new_n650), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n634), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n535), .A2(new_n571), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n519), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT45), .Z(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT109), .B1(new_n479), .B2(new_n524), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n418), .A2(KEYINPUT38), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n418), .A2(new_n416), .A3(KEYINPUT38), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n408), .A2(new_n410), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n574), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n477), .A3(new_n442), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n477), .B1(new_n519), .B2(new_n520), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT36), .B1(new_n515), .B2(new_n516), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n695), .A2(new_n696), .A3(new_n513), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n532), .B1(new_n688), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n687), .B1(new_n700), .B2(new_n682), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n682), .A2(new_n687), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n533), .A2(new_n534), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n571), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n519), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n708), .ZN(G1328gat));
  AOI21_X1  g508(.A(G36gat), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n658), .A2(new_n710), .ZN(new_n711));
  OR4_X1    g510(.A1(KEYINPUT110), .A2(new_n684), .A3(KEYINPUT46), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n707), .B2(new_n528), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n684), .A2(new_n711), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  OAI21_X1  g514(.A(G43gat), .B1(new_n707), .B2(new_n518), .ZN(new_n716));
  INV_X1    g515(.A(new_n517), .ZN(new_n717));
  OR3_X1    g516(.A1(new_n684), .A2(G43gat), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1330gat));
  INV_X1    g520(.A(new_n684), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n477), .A2(G50gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n701), .A2(new_n522), .A3(new_n703), .A4(new_n706), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G50gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(KEYINPUT48), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n726), .A2(new_n729), .B1(new_n722), .B2(new_n723), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n728), .B(KEYINPUT48), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n729), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n731), .A3(new_n724), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT112), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n727), .B1(new_n732), .B2(new_n736), .ZN(G1331gat));
  NAND2_X1  g536(.A1(new_n688), .A2(new_n699), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n531), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n634), .A2(new_n651), .ZN(new_n740));
  AND4_X1   g539(.A1(new_n705), .A2(new_n739), .A3(new_n740), .A4(new_n620), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n574), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n658), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT49), .B(G64gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(G1333gat));
  INV_X1    g546(.A(new_n518), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n598), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n717), .A2(G71gat), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n741), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n741), .A2(new_n522), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT114), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT113), .B(G78gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1335gat));
  INV_X1    g555(.A(new_n620), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(new_n571), .A3(new_n650), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n704), .A2(new_n574), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n587), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n571), .A2(new_n650), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n739), .A2(new_n634), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n739), .A2(KEYINPUT51), .A3(new_n634), .A4(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n757), .A2(new_n519), .A3(new_n587), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n760), .A2(new_n768), .ZN(G1336gat));
  NOR3_X1   g568(.A1(new_n757), .A2(G92gat), .A3(new_n528), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n701), .A2(new_n658), .A3(new_n703), .A4(new_n758), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n764), .A2(KEYINPUT115), .A3(new_n765), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n778), .A3(new_n763), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n779), .A3(new_n770), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n774), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n776), .B1(new_n781), .B2(KEYINPUT52), .ZN(new_n782));
  AOI211_X1 g581(.A(KEYINPUT116), .B(new_n772), .C1(new_n780), .C2(new_n774), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n775), .B1(new_n782), .B2(new_n783), .ZN(G1337gat));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n584), .A3(new_n517), .A4(new_n620), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n704), .A2(new_n748), .A3(new_n758), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n584), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n704), .A2(new_n522), .A3(new_n758), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n757), .A2(G106gat), .A3(new_n477), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT117), .Z(new_n791));
  NAND3_X1  g590(.A1(new_n777), .A2(new_n779), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT53), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT53), .B1(new_n766), .B2(new_n790), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n652), .A2(new_n705), .ZN(new_n798));
  INV_X1    g597(.A(new_n613), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n606), .A2(new_n611), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n614), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n577), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n612), .A2(new_n803), .A3(new_n613), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n541), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n561), .A2(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n570), .A2(new_n809), .B1(new_n810), .B2(new_n540), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n634), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n802), .A4(new_n804), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n619), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n808), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n807), .A2(new_n571), .A3(new_n619), .A4(new_n813), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n620), .A2(new_n811), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n634), .B1(new_n818), .B2(KEYINPUT118), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n815), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n798), .B1(new_n822), .B2(new_n650), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n574), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n658), .A2(new_n526), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n571), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n823), .A2(new_n477), .A3(new_n517), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n658), .A2(new_n519), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n239), .A3(new_n705), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n828), .A2(new_n832), .ZN(G1340gat));
  AOI21_X1  g632(.A(G120gat), .B1(new_n827), .B2(new_n620), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n831), .A2(new_n241), .A3(new_n757), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(G1341gat));
  INV_X1    g635(.A(new_n230), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n831), .B2(new_n651), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n824), .A2(new_n230), .A3(new_n650), .A4(new_n825), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT119), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1342gat));
  NOR3_X1   g643(.A1(new_n826), .A2(G134gat), .A3(new_n682), .ZN(new_n845));
  XOR2_X1   g644(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n831), .B2(new_n682), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n823), .A2(new_n851), .A3(new_n522), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n830), .A2(new_n518), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n818), .A2(new_n682), .ZN(new_n854));
  INV_X1    g653(.A(new_n815), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n650), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n798), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n522), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n853), .B1(new_n858), .B2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G141gat), .B1(new_n860), .B2(new_n705), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n748), .A2(new_n477), .A3(new_n658), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n824), .A2(new_n204), .A3(new_n571), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT58), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n861), .B(new_n865), .C1(new_n862), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1344gat));
  AND2_X1   g669(.A1(new_n824), .A2(new_n864), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n205), .A3(new_n620), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n851), .B1(new_n823), .B2(new_n522), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n856), .B1(new_n653), .B2(new_n705), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n522), .A2(new_n851), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n757), .B1(new_n853), .B2(KEYINPUT122), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n878), .B(new_n879), .C1(KEYINPUT122), .C2(new_n853), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n860), .A2(new_n757), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(KEYINPUT59), .A3(new_n205), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n872), .B1(new_n881), .B2(new_n883), .ZN(G1345gat));
  NAND3_X1  g683(.A1(new_n871), .A2(new_n212), .A3(new_n650), .ZN(new_n885));
  OAI21_X1  g684(.A(G155gat), .B1(new_n860), .B2(new_n651), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1346gat));
  NAND2_X1  g686(.A1(new_n216), .A2(new_n218), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n682), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n824), .A2(new_n864), .A3(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT123), .Z(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n860), .B2(new_n682), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n528), .A2(new_n574), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n823), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n526), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n571), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n894), .B(KEYINPUT124), .Z(new_n900));
  NAND2_X1  g699(.A1(new_n829), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n309), .A3(new_n705), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n899), .A2(new_n902), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n898), .B2(new_n620), .ZN(new_n904));
  INV_X1    g703(.A(new_n901), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n757), .B1(new_n338), .B2(new_n339), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(G1349gat));
  OAI21_X1  g706(.A(G183gat), .B1(new_n901), .B2(new_n651), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n895), .A2(new_n351), .A3(new_n896), .A4(new_n650), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT60), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n350), .A3(new_n634), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n829), .A2(new_n634), .A3(new_n900), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G190gat), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(KEYINPUT61), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(KEYINPUT61), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n748), .A2(new_n477), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n705), .A2(G197gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n895), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT125), .Z(new_n924));
  INV_X1    g723(.A(G197gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n900), .A2(new_n518), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n874), .A2(new_n877), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(new_n571), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n925), .B2(new_n928), .ZN(G1352gat));
  NOR2_X1   g728(.A1(new_n757), .A2(G204gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n895), .A2(new_n921), .A3(new_n930), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT62), .Z(new_n932));
  NAND2_X1  g731(.A1(new_n927), .A2(new_n620), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G204gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  NOR4_X1   g734(.A1(new_n874), .A2(new_n877), .A3(new_n651), .A4(new_n926), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n936), .A2(KEYINPUT63), .A3(new_n380), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(new_n380), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n895), .A2(new_n380), .A3(new_n650), .A4(new_n921), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(G1354gat));
  NAND4_X1  g740(.A1(new_n895), .A2(new_n381), .A3(new_n634), .A4(new_n921), .ZN(new_n942));
  NOR4_X1   g741(.A1(new_n874), .A2(new_n877), .A3(new_n682), .A4(new_n926), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n381), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n942), .B(KEYINPUT127), .C1(new_n943), .C2(new_n381), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1355gat));
endmodule


