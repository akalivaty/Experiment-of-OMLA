//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n912,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT82), .B(G22gat), .Z(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G228gat), .A2(G233gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n216), .A2(new_n218), .B1(KEYINPUT2), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n212), .B(new_n214), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n217), .A2(G141gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n215), .A2(G148gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT76), .B1(new_n226), .B2(KEYINPUT75), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n213), .B1(new_n220), .B2(new_n212), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n222), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT78), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231));
  INV_X1    g030(.A(G211gat), .ZN(new_n232));
  INV_X1    g031(.A(G218gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n235), .A2(G204gat), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(G204gat), .B1(new_n235), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G211gat), .B(G218gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(new_n234), .C1(new_n237), .C2(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G141gat), .B(G148gat), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT76), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n216), .A2(new_n218), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n221), .B1(new_n251), .B2(new_n223), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n250), .B(new_n213), .C1(new_n252), .C2(KEYINPUT76), .ZN(new_n253));
  AOI211_X1 g052(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n253), .C2(new_n222), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n229), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n245), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n244), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT81), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n247), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(KEYINPUT81), .A3(new_n259), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n211), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n211), .B1(new_n246), .B2(new_n229), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(new_n259), .B2(new_n258), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n209), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n229), .A2(new_n256), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT77), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n229), .A2(new_n255), .A3(new_n256), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT29), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n261), .B1(new_n271), .B2(new_n244), .ZN(new_n272));
  INV_X1    g071(.A(new_n247), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n263), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n210), .ZN(new_n275));
  INV_X1    g074(.A(new_n266), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n208), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n207), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(G22gat), .B1(new_n264), .B2(new_n266), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n277), .A3(new_n207), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n266), .B1(new_n274), .B2(new_n210), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n206), .B1(new_n283), .B2(new_n208), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(KEYINPUT83), .A3(new_n279), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n278), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G8gat), .B(G36gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT74), .ZN(new_n288));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(G226gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT64), .B(G169gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(G176gat), .ZN(new_n297));
  AOI211_X1 g096(.A(KEYINPUT25), .B(new_n294), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(KEYINPUT24), .ZN(new_n300));
  XNOR2_X1  g099(.A(G183gat), .B(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n302), .B2(KEYINPUT24), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT65), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n298), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT28), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(KEYINPUT26), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n294), .B1(new_n312), .B2(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n299), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n306), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n301), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT66), .B1(new_n322), .B2(new_n300), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n294), .B1(KEYINPUT23), .B2(new_n311), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n320), .A2(new_n323), .A3(new_n305), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT25), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n293), .B1(new_n327), .B2(new_n245), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n317), .B1(KEYINPUT25), .B2(new_n325), .ZN(new_n329));
  INV_X1    g128(.A(new_n293), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT72), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT72), .B1(new_n327), .B2(new_n293), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n244), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n330), .B1(new_n329), .B2(KEYINPUT29), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT73), .B1(new_n327), .B2(new_n293), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n338));
  AOI211_X1 g137(.A(new_n338), .B(new_n330), .C1(new_n318), .C2(new_n326), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n336), .B(new_n244), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n290), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n290), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n293), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n333), .B1(new_n345), .B2(KEYINPUT72), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n340), .B(new_n343), .C1(new_n346), .C2(new_n244), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(KEYINPUT30), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n335), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n340), .A4(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT0), .ZN(new_n354));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  XNOR2_X1  g157(.A(G127gat), .B(G134gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n362), .A2(G134gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364));
  OAI221_X1 g163(.A(new_n361), .B1(new_n360), .B2(new_n363), .C1(KEYINPUT1), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  OR3_X1    g167(.A1(new_n368), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n366), .A2(new_n367), .A3(new_n359), .A4(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n229), .ZN(new_n372));
  INV_X1    g171(.A(new_n229), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n358), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(KEYINPUT79), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n372), .B2(KEYINPUT4), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n229), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT69), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n365), .A2(KEYINPUT69), .A3(new_n370), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n383), .B(new_n385), .C1(new_n392), .C2(new_n382), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n269), .A2(new_n270), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n371), .B1(KEYINPUT3), .B2(new_n373), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n378), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n380), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n390), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT69), .B1(new_n365), .B2(new_n370), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n230), .A2(new_n400), .A3(new_n382), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n358), .A3(new_n396), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n357), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n383), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n382), .B1(new_n230), .B2(new_n400), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n395), .B1(new_n257), .B2(new_n254), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n377), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n379), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n356), .A3(new_n404), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n406), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n356), .B1(new_n413), .B2(new_n404), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT6), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n352), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n327), .A2(new_n391), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n329), .A2(new_n400), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G227gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n292), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT70), .ZN(new_n432));
  INV_X1    g231(.A(new_n427), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n423), .B2(new_n424), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT32), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n428), .B(KEYINPUT32), .C1(new_n429), .C2(new_n422), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n433), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n440), .B(KEYINPUT34), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(new_n441), .A3(new_n438), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n286), .A2(new_n419), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT35), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT87), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n278), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n284), .A2(KEYINPUT83), .A3(new_n279), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT83), .B1(new_n284), .B2(new_n279), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n351), .A2(new_n348), .B1(new_n415), .B2(new_n417), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n443), .A2(new_n444), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT35), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n454), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n414), .A2(new_n407), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n356), .B(KEYINPUT84), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n397), .B2(new_n405), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n417), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n352), .A3(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n457), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n286), .A2(new_n419), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n445), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n349), .A2(new_n471), .A3(new_n340), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n290), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n349), .B2(new_n340), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT38), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n459), .A2(new_n461), .B1(KEYINPUT6), .B2(new_n416), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n336), .B(new_n259), .C1(new_n337), .C2(new_n339), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT37), .B(new_n477), .C1(new_n346), .C2(new_n259), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(new_n478), .A3(new_n479), .A4(new_n290), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n476), .A3(new_n347), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n352), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n401), .A2(new_n402), .B1(new_n394), .B2(new_n395), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n377), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT39), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n460), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n372), .A2(new_n375), .A3(new_n377), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT39), .B(new_n487), .C1(new_n483), .C2(new_n377), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(KEYINPUT40), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n461), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT40), .B1(new_n486), .B2(new_n488), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n482), .A2(new_n492), .A3(KEYINPUT85), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n488), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n461), .A3(new_n489), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n494), .B1(new_n498), .B2(new_n352), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n468), .B(new_n470), .C1(new_n500), .C2(new_n286), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  NOR3_X1   g303(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(KEYINPUT89), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(KEYINPUT89), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n510), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n504), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n506), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n503), .A2(KEYINPUT15), .B1(new_n517), .B2(new_n505), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n512), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT17), .B1(new_n511), .B2(new_n519), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  AOI21_X1  g324(.A(G1gat), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(KEYINPUT91), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(KEYINPUT91), .C1(new_n525), .C2(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n523), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n511), .A2(new_n519), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n536), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OR3_X1    g344(.A1(new_n537), .A2(KEYINPUT93), .A3(new_n540), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n539), .B(KEYINPUT13), .Z(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n535), .A3(new_n532), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(KEYINPUT93), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n539), .A4(new_n542), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  INV_X1    g352(.A(G197gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT11), .B(G169gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT12), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n552), .B2(KEYINPUT88), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G190gat), .B(G218gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT100), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT101), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570));
  OAI211_X1 g369(.A(G85gat), .B(G92gat), .C1(new_n570), .C2(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(KEYINPUT96), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT97), .B(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n574), .A2(new_n575), .B1(KEYINPUT8), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n573), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n584), .B(new_n573), .C1(new_n579), .C2(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n523), .A3(KEYINPUT99), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT99), .B1(new_n586), .B2(new_n523), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n586), .B2(new_n540), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n567), .B(new_n569), .C1(new_n590), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n586), .A2(new_n523), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n597), .B2(new_n587), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n568), .B1(new_n598), .B2(new_n566), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n564), .A2(new_n565), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  AND3_X1   g401(.A1(new_n594), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n594), .B2(new_n599), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n607), .A2(G57gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(G57gat), .ZN(new_n609));
  INV_X1    g408(.A(G71gat), .ZN(new_n610));
  INV_X1    g409(.A(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI22_X1  g411(.A1(new_n608), .A2(new_n609), .B1(new_n612), .B2(KEYINPUT9), .ZN(new_n613));
  NOR2_X1   g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n616));
  OAI22_X1  g415(.A1(new_n612), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n613), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G127gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n537), .B1(new_n619), .B2(new_n618), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT95), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G155gat), .ZN(new_n628));
  XOR2_X1   g427(.A(G183gat), .B(G211gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n625), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n606), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n618), .B1(new_n585), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n586), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n583), .B(new_n585), .C1(new_n634), .C2(new_n618), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT10), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n586), .A2(new_n639), .A3(new_n618), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n633), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n633), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT103), .ZN(new_n645));
  XOR2_X1   g444(.A(G176gat), .B(G204gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n643), .A2(new_n647), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n632), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n502), .A2(new_n561), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n418), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n482), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G8gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(KEYINPUT42), .B2(new_n659), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n652), .A2(new_n662), .A3(new_n454), .ZN(new_n663));
  INV_X1    g462(.A(new_n470), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n665), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n652), .A2(new_n286), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n603), .B2(new_n604), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n594), .A2(new_n599), .ZN(new_n672));
  INV_X1    g471(.A(new_n602), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n594), .A2(new_n599), .A3(new_n602), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(KEYINPUT106), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n467), .B2(new_n501), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT35), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n456), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n458), .A2(new_n465), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n501), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n605), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n680), .B1(new_n686), .B2(KEYINPUT44), .ZN(new_n687));
  INV_X1    g486(.A(new_n561), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n650), .A2(new_n631), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT105), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT107), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n502), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n606), .B1(new_n467), .B2(new_n501), .ZN(new_n694));
  OAI22_X1  g493(.A1(new_n693), .A2(new_n679), .B1(new_n694), .B2(new_n678), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n690), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n692), .A2(new_n653), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n692), .A2(new_n697), .A3(new_n700), .A4(new_n653), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(G29gat), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n694), .A2(new_n689), .ZN(new_n703));
  INV_X1    g502(.A(G29gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n653), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(G1328gat));
  INV_X1    g506(.A(G36gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n708), .A3(new_n482), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  AND3_X1   g509(.A1(new_n692), .A2(new_n482), .A3(new_n697), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n708), .B2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n703), .A2(new_n713), .A3(new_n454), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n687), .A2(new_n470), .A3(new_n691), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT47), .B(new_n714), .C1(new_n715), .C2(new_n713), .ZN(new_n716));
  INV_X1    g515(.A(new_n714), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n692), .A2(new_n664), .A3(new_n697), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n203), .A3(new_n286), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n687), .A2(new_n452), .A3(new_n691), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT48), .B(new_n721), .C1(new_n722), .C2(new_n203), .ZN(new_n723));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n692), .A2(new_n286), .A3(new_n697), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(G50gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g526(.A(new_n650), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n632), .A2(new_n728), .A3(new_n561), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n502), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n418), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT109), .B(G57gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n352), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n730), .B2(new_n470), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n454), .A2(new_n610), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n730), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g541(.A1(new_n730), .A2(new_n452), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n611), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n631), .A2(new_n561), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n650), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n695), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n418), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n502), .A2(new_n605), .A3(new_n745), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n653), .A2(new_n574), .A3(new_n650), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n749), .A2(new_n574), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  NOR3_X1   g554(.A1(new_n728), .A2(new_n352), .A3(G92gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n748), .A2(new_n352), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(new_n575), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n757), .B(new_n761), .C1(new_n758), .C2(new_n575), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1337gat));
  AOI21_X1  g562(.A(new_n678), .B1(new_n502), .B2(new_n605), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n664), .B(new_n747), .C1(new_n764), .C2(new_n680), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n695), .A2(new_n767), .A3(new_n664), .A4(new_n747), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(G99gat), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n728), .A2(new_n445), .A3(G99gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1338gat));
  NOR2_X1   g575(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G106gat), .B1(new_n748), .B2(new_n452), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n452), .A2(new_n728), .A3(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n752), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n782));
  AND4_X1   g581(.A1(new_n778), .A2(new_n779), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n752), .A2(new_n780), .B1(KEYINPUT112), .B2(KEYINPUT53), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n778), .B1(new_n784), .B2(new_n779), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n783), .A2(new_n785), .ZN(G1339gat));
  INV_X1    g585(.A(new_n631), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n547), .B1(new_n546), .B2(new_n549), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n539), .B1(new_n538), .B2(new_n542), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n557), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n545), .A2(new_n550), .A3(new_n551), .A4(new_n558), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n648), .B2(new_n649), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n642), .A2(new_n639), .ZN(new_n795));
  INV_X1    g594(.A(new_n640), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n795), .A2(G230gat), .A3(G233gat), .A4(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n797), .A2(KEYINPUT54), .A3(new_n641), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(new_n633), .C1(new_n638), .C2(new_n640), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n647), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n794), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n649), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n797), .A2(KEYINPUT54), .A3(new_n641), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n647), .A4(new_n800), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n802), .A2(new_n561), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n677), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n802), .A2(new_n803), .A3(new_n792), .A4(new_n805), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n676), .B2(new_n671), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n787), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n632), .A2(new_n561), .A3(new_n650), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n458), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n482), .A2(new_n418), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n688), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n688), .A2(G113gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT113), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n815), .B2(new_n818), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n815), .B2(new_n728), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n650), .A2(new_n368), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT114), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n815), .B2(new_n822), .ZN(G1341gat));
  NOR2_X1   g622(.A1(new_n815), .A2(new_n787), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(new_n362), .ZN(G1342gat));
  NAND2_X1  g624(.A1(new_n352), .A2(new_n605), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT115), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(G134gat), .A3(new_n418), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT116), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT117), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n815), .B2(new_n606), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n832), .B(new_n833), .C1(KEYINPUT56), .C2(new_n830), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n810), .A2(new_n812), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT119), .A3(new_n653), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n664), .A2(new_n452), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT119), .B1(new_n835), .B2(new_n653), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n838), .A2(KEYINPUT121), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n688), .A2(G141gat), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT121), .B1(new_n838), .B2(new_n839), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n840), .A2(new_n352), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n470), .A2(new_n814), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n835), .B2(new_n286), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n286), .A2(KEYINPUT57), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n605), .B1(new_n806), .B2(new_n793), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n787), .B1(new_n809), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(new_n812), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n846), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n852), .A2(KEYINPUT122), .A3(new_n688), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT122), .B1(new_n852), .B2(new_n688), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G141gat), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n843), .B(new_n844), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n806), .A2(new_n793), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n671), .A2(new_n676), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n677), .A3(new_n792), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n631), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n286), .B1(new_n862), .B2(new_n811), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT118), .B1(new_n865), .B2(new_n845), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n846), .C1(new_n847), .C2(new_n851), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n868), .A3(new_n561), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G141gat), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n838), .A2(new_n839), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n352), .A3(new_n841), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT120), .B1(new_n873), .B2(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n875), .B(new_n844), .C1(new_n870), .C2(new_n872), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n856), .B1(new_n874), .B2(new_n876), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n866), .A2(new_n868), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n728), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(KEYINPUT59), .A3(new_n217), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n808), .A2(new_n606), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n787), .B1(new_n849), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n452), .B1(new_n812), .B2(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n884), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n835), .A2(KEYINPUT57), .A3(new_n286), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n884), .B2(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n650), .A3(new_n846), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n881), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n840), .A2(new_n842), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n352), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n650), .A2(new_n217), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n880), .A2(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n878), .B2(new_n787), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n787), .A2(G155gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(G1346gat));
  NOR2_X1   g696(.A1(new_n827), .A2(G162gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n840), .A2(new_n842), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(KEYINPUT124), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(KEYINPUT124), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n866), .A2(new_n868), .A3(new_n677), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G162gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n900), .A2(new_n901), .B1(new_n905), .B2(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n653), .A2(new_n352), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n813), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n688), .ZN(new_n910));
  MUX2_X1   g709(.A(G169gat), .B(new_n295), .S(new_n910), .Z(G1348gat));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n728), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g712(.A1(new_n909), .A2(new_n787), .ZN(new_n914));
  MUX2_X1   g713(.A(G183gat), .B(new_n307), .S(new_n914), .Z(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n909), .B2(new_n606), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n677), .A2(new_n308), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n909), .B2(new_n919), .ZN(G1351gat));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n888), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n470), .A2(new_n908), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n888), .A2(new_n921), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n554), .A3(new_n688), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n835), .A2(new_n837), .A3(new_n908), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n561), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n926), .A2(new_n929), .ZN(G1352gat));
  XNOR2_X1  g729(.A(KEYINPUT127), .B(G204gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n925), .B2(new_n728), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n927), .A2(new_n728), .A3(new_n931), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n232), .A3(new_n631), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n888), .A2(new_n631), .A3(new_n923), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1354gat));
  NOR3_X1   g739(.A1(new_n925), .A2(new_n233), .A3(new_n606), .ZN(new_n941));
  AOI21_X1  g740(.A(G218gat), .B1(new_n928), .B2(new_n677), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1355gat));
endmodule


