//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G143), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n189), .A2(G143), .ZN(new_n194));
  OAI22_X1  g008(.A1(new_n190), .A2(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n189), .A3(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT64), .B1(new_n192), .B2(G146), .ZN(new_n198));
  OAI211_X1 g012(.A(G128), .B(new_n197), .C1(new_n198), .C2(new_n193), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G137), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n207), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(new_n197), .C1(new_n198), .C2(new_n193), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n216), .B(new_n219), .C1(new_n193), .C2(new_n194), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n218), .B2(new_n220), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n212), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT30), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(KEYINPUT67), .A3(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(new_n220), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n215), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n215), .A3(KEYINPUT68), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(KEYINPUT30), .A3(new_n212), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n225), .A2(new_n247), .A3(new_n226), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n228), .A2(new_n239), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n215), .A3(new_n222), .ZN(new_n252));
  AOI211_X1 g066(.A(KEYINPUT66), .B(KEYINPUT30), .C1(new_n252), .C2(new_n212), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n247), .B1(new_n225), .B2(new_n226), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n239), .A4(new_n246), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT70), .A2(G237), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT70), .A2(G237), .ZN(new_n260));
  AOI21_X1  g074(.A(G953), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n244), .A2(new_n245), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n238), .A3(new_n212), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n250), .A2(new_n257), .A3(new_n265), .A4(new_n267), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n273));
  INV_X1    g087(.A(new_n267), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n238), .B1(new_n252), .B2(new_n212), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n212), .A2(new_n238), .A3(new_n242), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(KEYINPUT28), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT72), .B1(new_n272), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n283), .B(new_n280), .C1(new_n268), .C2(new_n271), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT32), .B(new_n187), .C1(new_n282), .C2(new_n284), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n238), .B1(new_n266), .B2(new_n212), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n274), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n278), .B1(new_n290), .B2(KEYINPUT28), .ZN(new_n291));
  INV_X1    g105(.A(new_n265), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n250), .A2(new_n257), .A3(new_n267), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n298), .B2(new_n265), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(KEYINPUT73), .A3(new_n292), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n293), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n276), .A2(new_n265), .A3(new_n279), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G472), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n287), .A2(new_n288), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  XNOR2_X1  g120(.A(G125), .B(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n309), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(G146), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n307), .B(KEYINPUT77), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n189), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n191), .A2(G119), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT74), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT24), .B(G110), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT76), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  MUX2_X1   g137(.A(new_n323), .B(new_n322), .S(new_n315), .Z(new_n324));
  INV_X1    g138(.A(G110), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n311), .B(new_n313), .C1(new_n321), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n308), .A2(new_n310), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n189), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n311), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n324), .B(KEYINPUT75), .Z(new_n332));
  OAI221_X1 g146(.A(new_n331), .B1(new_n318), .B2(new_n319), .C1(new_n332), .C2(new_n325), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n328), .A2(KEYINPUT78), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT78), .B1(new_n328), .B2(new_n333), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT22), .B(G137), .Z(new_n336));
  INV_X1    g150(.A(G221), .ZN(new_n337));
  INV_X1    g151(.A(G234), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n337), .A2(new_n338), .A3(G953), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n336), .B(new_n339), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n334), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  AOI211_X1 g156(.A(KEYINPUT78), .B(new_n342), .C1(new_n328), .C2(new_n333), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n306), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT25), .B(new_n306), .C1(new_n341), .C2(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n306), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n341), .A2(new_n343), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(G902), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G469), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n306), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT80), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n362), .B(G101), .C1(new_n365), .C2(new_n361), .ZN(new_n366));
  OR3_X1    g180(.A1(new_n360), .A2(KEYINPUT3), .A3(G107), .ZN(new_n367));
  INV_X1    g181(.A(G101), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n363), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n366), .A2(new_n370), .A3(KEYINPUT81), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n200), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n197), .B1(new_n198), .B2(new_n193), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n191), .B2(new_n190), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n371), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n215), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n359), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n378), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n370), .A3(new_n366), .ZN(new_n384));
  INV_X1    g198(.A(new_n374), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT81), .B1(new_n366), .B2(new_n370), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(new_n200), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n215), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n381), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n367), .A2(new_n363), .A3(new_n369), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n396), .B2(KEYINPUT4), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n398), .A4(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n370), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n241), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n215), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n373), .A2(KEYINPUT10), .A3(new_n200), .A4(new_n374), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n393), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  INV_X1    g220(.A(G953), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(G227), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n406), .B(new_n408), .Z(new_n409));
  AND2_X1   g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n391), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n393), .A2(new_n402), .A3(new_n404), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n215), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n405), .ZN(new_n414));
  INV_X1    g228(.A(new_n409), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n358), .B1(new_n417), .B2(new_n357), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n391), .A2(new_n405), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n413), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G469), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT9), .B(G234), .Z(new_n424));
  AOI21_X1  g238(.A(new_n337), .B1(new_n424), .B2(new_n306), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n239), .A2(new_n400), .A3(new_n401), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n314), .A3(G116), .ZN(new_n430));
  OAI211_X1 g244(.A(G113), .B(new_n430), .C1(new_n230), .C2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n234), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n385), .A2(new_n432), .A3(new_n386), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(G110), .B(G122), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n428), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n200), .A2(new_n309), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n309), .B2(new_n240), .ZN(new_n442));
  INV_X1    g256(.A(G224), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n442), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n447), .A3(new_n436), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n440), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n442), .B1(new_n450), .B2(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT7), .B(new_n445), .C1(new_n442), .C2(new_n450), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n436), .B(KEYINPUT8), .Z(new_n455));
  AND2_X1   g269(.A1(new_n432), .A2(new_n371), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n433), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .A4(new_n439), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n449), .A2(new_n306), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n449), .A2(new_n306), .A3(new_n460), .A4(new_n458), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n427), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n360), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n259), .A2(new_n260), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(G214), .A3(new_n407), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n192), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT18), .B(G131), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(KEYINPUT84), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT18), .A4(G131), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n313), .B1(new_n189), .B2(new_n307), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(G131), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n472), .A2(new_n206), .A3(new_n473), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT19), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n307), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n307), .A2(new_n486), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n312), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n487), .B1(new_n489), .B2(new_n485), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n311), .B(new_n484), .C1(new_n490), .C2(G146), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n469), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n494), .A3(new_n483), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n206), .B1(new_n472), .B2(new_n473), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n331), .B1(KEYINPUT17), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n494), .A4(new_n483), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n481), .A3(new_n469), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT20), .ZN(new_n504));
  INV_X1    g318(.A(G475), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n306), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n501), .A2(new_n481), .A3(new_n469), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n505), .B(new_n306), .C1(new_n507), .C2(new_n492), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n469), .B1(new_n501), .B2(new_n481), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n306), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT87), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(new_n306), .C1(new_n507), .C2(new_n511), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(G475), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(G234), .A2(G237), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n518), .A2(G952), .A3(new_n407), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(G902), .A3(G953), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n520), .B(KEYINPUT92), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT21), .B(G898), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n519), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G116), .B(G122), .ZN(new_n526));
  INV_X1    g340(.A(G107), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G128), .B(G143), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n202), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT89), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(KEYINPUT13), .ZN(new_n532));
  OR3_X1    g346(.A1(new_n191), .A2(KEYINPUT13), .A3(G143), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(G134), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n528), .B(new_n531), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT14), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n526), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G116), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT14), .A3(G122), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(G107), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n526), .A2(new_n527), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n529), .B(new_n202), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n424), .A2(G217), .A3(new_n407), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n553));
  INV_X1    g367(.A(new_n551), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n538), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(KEYINPUT91), .A3(new_n551), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n306), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G478), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n558), .B(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n517), .A2(new_n525), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n467), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n305), .A2(new_n356), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  AND2_X1   g379(.A1(new_n269), .A2(new_n270), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n269), .A2(new_n270), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n281), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n283), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n272), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n285), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n556), .A2(new_n574), .A3(new_n557), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT93), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n556), .A2(new_n577), .A3(new_n574), .A4(new_n557), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n552), .A2(KEYINPUT33), .A3(new_n555), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n559), .A2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n558), .A2(new_n559), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n517), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n525), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n464), .A2(new_n465), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR4_X1   g402(.A1(new_n573), .A2(new_n355), .A3(new_n427), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  OAI21_X1  g405(.A(new_n306), .B1(new_n282), .B2(new_n284), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n569), .A2(new_n570), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n592), .A2(G472), .B1(new_n593), .B2(new_n187), .ZN(new_n594));
  INV_X1    g408(.A(new_n427), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n510), .A2(KEYINPUT94), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n510), .A2(KEYINPUT94), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n516), .B(new_n561), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n587), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n594), .A2(new_n356), .A3(new_n595), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT95), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  NAND2_X1  g417(.A1(new_n328), .A2(new_n333), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n348), .A2(new_n350), .B1(new_n353), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n594), .A2(new_n563), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT37), .B(G110), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G12));
  AND2_X1   g425(.A1(new_n305), .A2(new_n608), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT96), .B(G900), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n522), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n519), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n598), .A2(new_n466), .A3(new_n427), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  XOR2_X1   g434(.A(new_n616), .B(KEYINPUT39), .Z(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n595), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n623), .A2(KEYINPUT40), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n607), .B1(new_n623), .B2(KEYINPUT40), .ZN(new_n625));
  INV_X1    g439(.A(new_n465), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n290), .A2(new_n292), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n269), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n306), .B1(new_n629), .B2(KEYINPUT97), .ZN(new_n631));
  OAI21_X1  g445(.A(G472), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n287), .A2(new_n288), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n464), .B(KEYINPUT38), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n517), .A2(new_n561), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n627), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  NAND3_X1  g453(.A1(new_n517), .A2(new_n584), .A3(new_n616), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n517), .A2(new_n584), .A3(KEYINPUT98), .A4(new_n616), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n467), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n612), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G146), .ZN(G48));
  AND2_X1   g460(.A1(new_n305), .A2(new_n356), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n417), .A2(new_n357), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n417), .A2(new_n357), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n426), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n588), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT41), .B(G113), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G15));
  NOR3_X1   g468(.A1(new_n598), .A2(new_n587), .A3(new_n650), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G116), .ZN(G18));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n466), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n305), .A2(new_n562), .A3(new_n608), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G119), .ZN(G21));
  NOR4_X1   g474(.A1(new_n636), .A2(new_n650), .A3(new_n466), .A4(new_n525), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n272), .B1(new_n265), .B2(new_n291), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n187), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT99), .B(G472), .Z(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n571), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n666), .A2(new_n667), .A3(new_n355), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n592), .A2(new_n664), .B1(new_n187), .B2(new_n662), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT100), .B1(new_n669), .B2(new_n356), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n661), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  NAND2_X1  g486(.A1(new_n642), .A2(new_n643), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n669), .A3(new_n608), .A4(new_n658), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G125), .ZN(G27));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n422), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n419), .A2(new_n415), .B1(new_n410), .B2(new_n413), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(KEYINPUT101), .A3(G469), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n418), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n425), .A2(new_n626), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n462), .A2(new_n463), .A3(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT102), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT102), .B1(new_n681), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n673), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n288), .A2(KEYINPUT104), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(new_n287), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n285), .A2(KEYINPUT104), .A3(new_n286), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n304), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n688), .B(new_n356), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n691), .A2(new_n304), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n287), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n355), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n688), .ZN(new_n699));
  INV_X1    g513(.A(new_n686), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n647), .A2(new_n674), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n694), .A2(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n206), .ZN(G33));
  NOR2_X1   g518(.A1(new_n598), .A2(new_n617), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n305), .A2(new_n700), .A3(new_n356), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  INV_X1    g521(.A(new_n584), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n517), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n708), .B2(new_n517), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n573), .A4(new_n608), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n462), .A2(new_n465), .A3(new_n463), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(KEYINPUT45), .A2(G469), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n422), .A2(KEYINPUT106), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n722), .B(G469), .C1(new_n679), .C2(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n679), .A2(KEYINPUT45), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n358), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n649), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT46), .B1(new_n725), .B2(new_n726), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n426), .A3(new_n622), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n713), .A2(new_n573), .A3(new_n608), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n714), .A2(KEYINPUT107), .A3(new_n716), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n719), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT108), .B(G137), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G39));
  OAI21_X1  g552(.A(new_n426), .B1(new_n728), .B2(new_n729), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n742), .B1(new_n739), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n305), .A2(new_n356), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n674), .A3(new_n716), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  OR2_X1    g563(.A1(new_n668), .A2(new_n670), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n713), .A2(new_n519), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n658), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n650), .A2(new_n715), .A3(new_n615), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n713), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n697), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT48), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(G952), .A3(new_n407), .ZN(new_n760));
  INV_X1    g574(.A(new_n756), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n633), .A2(new_n355), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(new_n585), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n755), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n746), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n648), .A2(new_n649), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT115), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n425), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n715), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n634), .A2(new_n465), .A3(new_n650), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(KEYINPUT50), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n752), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n752), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT50), .B1(new_n773), .B2(new_n770), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n762), .A2(new_n517), .A3(new_n584), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n757), .A2(new_n608), .A3(new_n669), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT51), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n777), .A3(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(KEYINPUT51), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n772), .A2(new_n774), .A3(new_n782), .A4(new_n779), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n764), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n305), .B(new_n608), .C1(new_n618), .C2(new_n644), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n607), .A2(new_n616), .A3(new_n681), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n636), .A2(new_n466), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n633), .A2(new_n786), .A3(new_n426), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n788), .A3(new_n675), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n788), .A3(KEYINPUT52), .A4(new_n675), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n794), .B1(new_n789), .B2(new_n790), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n510), .A2(new_n516), .A3(new_n561), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n587), .B1(new_n585), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n594), .A2(new_n356), .A3(new_n595), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n564), .A2(new_n609), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n305), .B(new_n356), .C1(new_n655), .C2(new_n651), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n659), .A3(new_n671), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n700), .A2(new_n608), .A3(new_n674), .A4(new_n669), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n706), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n427), .A2(new_n617), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n516), .B1(new_n596), .B2(new_n597), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n561), .A3(new_n715), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n305), .A2(new_n608), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n808), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n703), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n798), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n701), .A2(new_n702), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n698), .B1(new_n697), .B2(new_n688), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n671), .A2(new_n804), .A3(new_n659), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n802), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n812), .A2(new_n813), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n812), .A2(new_n813), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n807), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n823), .A2(new_n825), .A3(new_n793), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n818), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n796), .B1(new_n793), .B2(new_n794), .ZN(new_n834));
  AND4_X1   g648(.A1(KEYINPUT53), .A2(new_n564), .A3(new_n609), .A4(new_n801), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n808), .C1(new_n814), .C2(new_n815), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n671), .A2(new_n804), .A3(new_n839), .A4(new_n659), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n841), .A3(new_n823), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n784), .A2(new_n831), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(G952), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n407), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n356), .A2(new_n682), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT110), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(KEYINPUT110), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n709), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(KEYINPUT111), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n633), .B1(new_n852), .B2(KEYINPUT111), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n766), .B(KEYINPUT49), .Z(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n635), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n847), .A2(new_n856), .ZN(G75));
  NAND2_X1  g671(.A1(new_n845), .A2(G953), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT118), .Z(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n832), .B1(new_n834), .B2(new_n842), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(G902), .ZN(new_n863));
  INV_X1    g677(.A(G210), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n440), .A2(new_n448), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(new_n446), .Z(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n868), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n861), .B(new_n870), .C1(new_n863), .C2(new_n864), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n860), .B1(new_n869), .B2(new_n871), .ZN(G51));
  XNOR2_X1  g686(.A(new_n358), .B(KEYINPUT57), .ZN(new_n873));
  INV_X1    g687(.A(new_n843), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n836), .B1(new_n838), .B2(new_n840), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n798), .A2(new_n875), .A3(new_n823), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n833), .B1(new_n876), .B2(new_n832), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n411), .A2(new_n416), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT119), .Z(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n863), .A2(new_n725), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n860), .B1(new_n881), .B2(new_n882), .ZN(G54));
  AOI21_X1  g697(.A(new_n306), .B1(new_n876), .B2(new_n832), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n503), .ZN(new_n886));
  INV_X1    g700(.A(new_n503), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n860), .B1(new_n886), .B2(new_n888), .ZN(G60));
  AND2_X1   g703(.A1(new_n579), .A2(new_n580), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n831), .A2(new_n843), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT59), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n893), .ZN(new_n895));
  INV_X1    g709(.A(new_n877), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n896), .B2(new_n843), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n894), .A2(new_n897), .A3(new_n860), .ZN(G63));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT60), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n842), .A2(new_n834), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n817), .B2(new_n793), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n606), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n859), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n352), .B1(new_n862), .B2(new_n901), .ZN(new_n906));
  XNOR2_X1  g720(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n900), .B1(new_n876), .B2(new_n832), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n860), .B1(new_n910), .B2(new_n606), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n862), .A2(new_n901), .ZN(new_n912));
  INV_X1    g726(.A(new_n352), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n907), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n909), .A2(new_n915), .ZN(G66));
  OAI21_X1  g730(.A(G953), .B1(new_n524), .B2(new_n443), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n825), .B2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n866), .B1(G898), .B2(new_n407), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G69));
  AOI21_X1  g734(.A(new_n407), .B1(G227), .B2(G900), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT124), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n785), .A2(new_n675), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n638), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n623), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n585), .A2(new_n799), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n647), .A2(new_n926), .A3(new_n716), .A4(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n736), .A2(new_n925), .A3(new_n748), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n638), .ZN(new_n930));
  OR2_X1    g744(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n407), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n255), .A2(new_n246), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n490), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(G900), .A2(G953), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n697), .A2(new_n787), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n706), .B1(new_n944), .B2(new_n731), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n703), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n736), .A2(new_n923), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT123), .B1(new_n736), .B2(new_n923), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n748), .B(new_n946), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n936), .B(new_n943), .C1(new_n951), .C2(G953), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n922), .B1(new_n942), .B2(new_n952), .ZN(new_n953));
  AND4_X1   g767(.A1(new_n922), .A2(new_n952), .A3(new_n939), .A4(new_n941), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  NAND3_X1  g771(.A1(new_n299), .A2(new_n269), .A3(new_n300), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n819), .A2(new_n830), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n297), .B(KEYINPUT125), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n265), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n736), .A2(new_n928), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n925), .A2(new_n748), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n825), .A4(new_n932), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(new_n957), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n967), .B(new_n961), .C1(new_n964), .C2(new_n957), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n859), .B(new_n959), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n947), .B(new_n948), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n748), .A3(new_n825), .A4(new_n946), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n972), .B2(new_n957), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n970), .B(new_n957), .C1(new_n951), .C2(new_n805), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n960), .A2(new_n265), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(G57));
endmodule


