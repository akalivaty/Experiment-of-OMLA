

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768;

  NOR2_X1 U376 ( .A1(G953), .A2(G237), .ZN(n496) );
  XNOR2_X2 U377 ( .A(n392), .B(KEYINPUT39), .ZN(n527) );
  NOR2_X1 U378 ( .A1(n598), .A2(n530), .ZN(n370) );
  XNOR2_X1 U379 ( .A(n380), .B(n379), .ZN(n766) );
  NAND2_X1 U380 ( .A1(n536), .A2(n684), .ZN(n605) );
  XNOR2_X1 U381 ( .A(n602), .B(KEYINPUT42), .ZN(n768) );
  NAND2_X1 U382 ( .A1(n416), .A2(n415), .ZN(n419) );
  XNOR2_X1 U383 ( .A(n406), .B(KEYINPUT19), .ZN(n606) );
  AND2_X1 U384 ( .A1(n595), .A2(n532), .ZN(n360) );
  XNOR2_X1 U385 ( .A(n370), .B(n365), .ZN(n521) );
  INV_X2 U386 ( .A(n596), .ZN(n464) );
  XNOR2_X1 U387 ( .A(n550), .B(n519), .ZN(n701) );
  XNOR2_X1 U388 ( .A(n578), .B(KEYINPUT101), .ZN(n598) );
  OR2_X1 U389 ( .A1(n657), .A2(G902), .ZN(n481) );
  XNOR2_X1 U390 ( .A(n412), .B(G125), .ZN(n489) );
  INV_X1 U391 ( .A(KEYINPUT64), .ZN(n451) );
  XNOR2_X1 U392 ( .A(n535), .B(n534), .ZN(n536) );
  NAND2_X1 U393 ( .A1(n419), .A2(n413), .ZN(n535) );
  BUF_X1 U394 ( .A(n486), .Z(n355) );
  BUF_X1 U395 ( .A(n640), .Z(n356) );
  XNOR2_X1 U396 ( .A(n625), .B(KEYINPUT85), .ZN(n640) );
  NOR2_X1 U397 ( .A1(n565), .A2(n464), .ZN(n669) );
  AND2_X2 U398 ( .A1(n642), .A2(n722), .ZN(n357) );
  XNOR2_X1 U399 ( .A(n754), .B(n430), .ZN(n358) );
  XNOR2_X1 U400 ( .A(n754), .B(n430), .ZN(n479) );
  XNOR2_X2 U401 ( .A(n592), .B(n591), .ZN(n636) );
  XNOR2_X2 U402 ( .A(n486), .B(n429), .ZN(n754) );
  XNOR2_X2 U403 ( .A(n511), .B(n404), .ZN(n486) );
  XNOR2_X1 U404 ( .A(n489), .B(n444), .ZN(n495) );
  XNOR2_X1 U405 ( .A(KEYINPUT10), .B(KEYINPUT71), .ZN(n444) );
  NAND2_X1 U406 ( .A1(n550), .A2(n700), .ZN(n406) );
  NAND2_X1 U407 ( .A1(n399), .A2(n397), .ZN(n403) );
  NOR2_X1 U408 ( .A1(n705), .A2(n398), .ZN(n397) );
  INV_X1 U409 ( .A(KEYINPUT47), .ZN(n402) );
  NOR2_X1 U410 ( .A1(n669), .A2(n764), .ZN(n572) );
  XNOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT97), .ZN(n411) );
  XNOR2_X1 U412 ( .A(KEYINPUT5), .B(G137), .ZN(n431) );
  XNOR2_X1 U413 ( .A(n435), .B(KEYINPUT3), .ZN(n437) );
  INV_X1 U414 ( .A(KEYINPUT75), .ZN(n435) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n428) );
  NAND2_X1 U416 ( .A1(n389), .A2(KEYINPUT41), .ZN(n388) );
  OR2_X1 U417 ( .A1(n701), .A2(n593), .ZN(n391) );
  XNOR2_X1 U418 ( .A(n452), .B(n396), .ZN(n507) );
  INV_X1 U419 ( .A(KEYINPUT8), .ZN(n396) );
  XNOR2_X1 U420 ( .A(G119), .B(G110), .ZN(n448) );
  XNOR2_X1 U421 ( .A(n495), .B(n409), .ZN(n504) );
  XOR2_X1 U422 ( .A(G137), .B(G140), .Z(n472) );
  XNOR2_X1 U423 ( .A(n422), .B(n382), .ZN(n651) );
  NAND2_X1 U424 ( .A1(n521), .A2(n522), .ZN(n392) );
  AND2_X1 U425 ( .A1(n606), .A2(n362), .ZN(n551) );
  BUF_X1 U426 ( .A(n618), .Z(n381) );
  XNOR2_X1 U427 ( .A(n403), .B(n402), .ZN(n612) );
  INV_X1 U428 ( .A(G146), .ZN(n412) );
  XNOR2_X1 U429 ( .A(KEYINPUT73), .B(KEYINPUT48), .ZN(n616) );
  INV_X1 U430 ( .A(G237), .ZN(n441) );
  XOR2_X1 U431 ( .A(G122), .B(G104), .Z(n498) );
  XOR2_X1 U432 ( .A(G116), .B(G107), .Z(n510) );
  XOR2_X1 U433 ( .A(KEYINPUT96), .B(G131), .Z(n500) );
  XNOR2_X1 U434 ( .A(G113), .B(G143), .ZN(n499) );
  XNOR2_X1 U435 ( .A(n410), .B(n497), .ZN(n409) );
  XNOR2_X1 U436 ( .A(n494), .B(n411), .ZN(n410) );
  XNOR2_X1 U437 ( .A(G140), .B(KEYINPUT11), .ZN(n494) );
  XNOR2_X1 U438 ( .A(n421), .B(G101), .ZN(n487) );
  INV_X1 U439 ( .A(KEYINPUT69), .ZN(n421) );
  XNOR2_X1 U440 ( .A(n424), .B(n407), .ZN(n423) );
  XNOR2_X1 U441 ( .A(n487), .B(n408), .ZN(n407) );
  XNOR2_X1 U442 ( .A(n489), .B(KEYINPUT18), .ZN(n424) );
  XNOR2_X1 U443 ( .A(KEYINPUT17), .B(KEYINPUT81), .ZN(n408) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n465) );
  XNOR2_X1 U445 ( .A(n594), .B(KEYINPUT1), .ZN(n618) );
  XNOR2_X1 U446 ( .A(n479), .B(n439), .ZN(n643) );
  XOR2_X1 U447 ( .A(G122), .B(KEYINPUT9), .Z(n509) );
  XNOR2_X1 U448 ( .A(KEYINPUT80), .B(G107), .ZN(n474) );
  XNOR2_X1 U449 ( .A(G104), .B(G110), .ZN(n473) );
  NAND2_X1 U450 ( .A1(n387), .A2(n384), .ZN(n698) );
  AND2_X1 U451 ( .A1(n391), .A2(n388), .ZN(n387) );
  NOR2_X1 U452 ( .A1(n663), .A2(n414), .ZN(n413) );
  NAND2_X1 U453 ( .A1(n620), .A2(n700), .ZN(n414) );
  AND2_X1 U454 ( .A1(n687), .A2(n533), .ZN(n420) );
  NAND2_X1 U455 ( .A1(n606), .A2(n401), .ZN(n398) );
  INV_X1 U456 ( .A(n600), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n453), .B(n395), .ZN(n454) );
  AND2_X1 U458 ( .A1(n507), .A2(G221), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n527), .A2(n526), .ZN(n405) );
  INV_X1 U460 ( .A(KEYINPUT35), .ZN(n379) );
  NAND2_X1 U461 ( .A1(n555), .A2(n554), .ZN(n380) );
  XNOR2_X1 U462 ( .A(n553), .B(n552), .ZN(n555) );
  XNOR2_X1 U463 ( .A(n426), .B(n425), .ZN(n677) );
  XNOR2_X1 U464 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n425) );
  NAND2_X1 U465 ( .A1(n399), .A2(n400), .ZN(n673) );
  INV_X1 U466 ( .A(n398), .ZN(n400) );
  NAND2_X1 U467 ( .A1(n573), .A2(n563), .ZN(n564) );
  INV_X1 U468 ( .A(KEYINPUT60), .ZN(n373) );
  INV_X1 U469 ( .A(KEYINPUT56), .ZN(n375) );
  AND2_X1 U470 ( .A1(n492), .A2(G210), .ZN(n359) );
  XNOR2_X1 U471 ( .A(G110), .B(KEYINPUT16), .ZN(n361) );
  OR2_X1 U472 ( .A1(n549), .A2(n548), .ZN(n362) );
  AND2_X1 U473 ( .A1(n720), .A2(n630), .ZN(n363) );
  AND2_X1 U474 ( .A1(n419), .A2(n418), .ZN(n364) );
  XNOR2_X1 U475 ( .A(n582), .B(KEYINPUT102), .ZN(n663) );
  XOR2_X1 U476 ( .A(n443), .B(KEYINPUT106), .Z(n365) );
  XOR2_X1 U477 ( .A(n653), .B(n654), .Z(n366) );
  XOR2_X1 U478 ( .A(n651), .B(n650), .Z(n367) );
  AND2_X1 U479 ( .A1(n635), .A2(n371), .ZN(n368) );
  OR2_X1 U480 ( .A1(n484), .A2(G952), .ZN(n660) );
  AND2_X1 U481 ( .A1(KEYINPUT2), .A2(KEYINPUT68), .ZN(n369) );
  NAND2_X1 U482 ( .A1(n629), .A2(n363), .ZN(n372) );
  NAND2_X1 U483 ( .A1(n372), .A2(n368), .ZN(n642) );
  NAND2_X1 U484 ( .A1(n630), .A2(n369), .ZN(n371) );
  BUF_X2 U485 ( .A(n732), .Z(n733) );
  XNOR2_X1 U486 ( .A(n374), .B(n373), .ZN(G60) );
  NAND2_X1 U487 ( .A1(n377), .A2(n660), .ZN(n374) );
  XNOR2_X1 U488 ( .A(n376), .B(n375), .ZN(G51) );
  NAND2_X1 U489 ( .A1(n378), .A2(n660), .ZN(n376) );
  XNOR2_X1 U490 ( .A(n655), .B(n366), .ZN(n377) );
  XNOR2_X1 U491 ( .A(n652), .B(n367), .ZN(n378) );
  NOR2_X2 U492 ( .A1(n589), .A2(n588), .ZN(n592) );
  XNOR2_X2 U493 ( .A(n440), .B(G472), .ZN(n578) );
  INV_X1 U494 ( .A(n739), .ZN(n382) );
  XNOR2_X1 U495 ( .A(n383), .B(n491), .ZN(n739) );
  XNOR2_X1 U496 ( .A(n490), .B(n361), .ZN(n383) );
  NAND2_X1 U497 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U498 ( .A1(n701), .A2(n385), .ZN(n384) );
  NOR2_X1 U499 ( .A1(n703), .A2(n386), .ZN(n385) );
  NAND2_X1 U500 ( .A1(n700), .A2(n593), .ZN(n386) );
  NAND2_X1 U501 ( .A1(n390), .A2(n700), .ZN(n389) );
  INV_X1 U502 ( .A(n703), .ZN(n390) );
  NAND2_X1 U503 ( .A1(n393), .A2(n615), .ZN(n617) );
  XNOR2_X1 U504 ( .A(n394), .B(n604), .ZN(n393) );
  NAND2_X1 U505 ( .A1(n603), .A2(n768), .ZN(n394) );
  XNOR2_X2 U506 ( .A(n405), .B(n529), .ZN(n603) );
  NOR2_X1 U507 ( .A1(n600), .A2(n601), .ZN(n607) );
  INV_X1 U508 ( .A(n601), .ZN(n401) );
  XNOR2_X2 U509 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n404) );
  XNOR2_X2 U510 ( .A(G143), .B(G128), .ZN(n511) );
  XNOR2_X1 U511 ( .A(n423), .B(n488), .ZN(n422) );
  NAND2_X1 U512 ( .A1(n420), .A2(n360), .ZN(n415) );
  NAND2_X1 U513 ( .A1(n417), .A2(KEYINPUT105), .ZN(n416) );
  NAND2_X1 U514 ( .A1(n360), .A2(n687), .ZN(n417) );
  NOR2_X1 U515 ( .A1(n663), .A2(n530), .ZN(n418) );
  INV_X1 U516 ( .A(n527), .ZN(n524) );
  NAND2_X1 U517 ( .A1(n696), .A2(n580), .ZN(n426) );
  XNOR2_X2 U518 ( .A(n551), .B(KEYINPUT0), .ZN(n580) );
  BUF_X1 U519 ( .A(n550), .Z(n620) );
  AND2_X2 U520 ( .A1(n642), .A2(n722), .ZN(n732) );
  XOR2_X1 U521 ( .A(n468), .B(KEYINPUT104), .Z(n427) );
  INV_X1 U522 ( .A(n618), .ZN(n539) );
  INV_X1 U523 ( .A(KEYINPUT76), .ZN(n447) );
  XNOR2_X1 U524 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U525 ( .A(n450), .B(n449), .ZN(n453) );
  INV_X1 U526 ( .A(KEYINPUT22), .ZN(n560) );
  INV_X1 U527 ( .A(KEYINPUT41), .ZN(n593) );
  INV_X1 U528 ( .A(KEYINPUT36), .ZN(n534) );
  XNOR2_X1 U529 ( .A(n734), .B(KEYINPUT118), .ZN(n735) );
  XNOR2_X1 U530 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U531 ( .A(n428), .B(KEYINPUT72), .ZN(n429) );
  XNOR2_X1 U532 ( .A(n487), .B(G146), .ZN(n430) );
  NAND2_X1 U533 ( .A1(n496), .A2(G210), .ZN(n432) );
  XNOR2_X1 U534 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U535 ( .A(G116), .B(KEYINPUT94), .ZN(n433) );
  XNOR2_X1 U536 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U537 ( .A(G119), .B(G113), .ZN(n436) );
  XNOR2_X1 U538 ( .A(n437), .B(n436), .ZN(n490) );
  XNOR2_X1 U539 ( .A(n438), .B(n490), .ZN(n439) );
  OR2_X2 U540 ( .A1(n643), .A2(G902), .ZN(n440) );
  INV_X1 U541 ( .A(G902), .ZN(n442) );
  NAND2_X1 U542 ( .A1(n442), .A2(n441), .ZN(n492) );
  NAND2_X1 U543 ( .A1(n492), .A2(G214), .ZN(n700) );
  INV_X1 U544 ( .A(n700), .ZN(n530) );
  XNOR2_X1 U545 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n443) );
  XOR2_X1 U546 ( .A(n495), .B(n472), .Z(n756) );
  XOR2_X1 U547 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n446) );
  XNOR2_X1 U548 ( .A(G128), .B(KEYINPUT23), .ZN(n445) );
  XNOR2_X1 U549 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X2 U550 ( .A(n451), .B(G953), .ZN(n484) );
  NAND2_X1 U551 ( .A1(n484), .A2(G234), .ZN(n452) );
  XNOR2_X1 U552 ( .A(n756), .B(n454), .ZN(n734) );
  NOR2_X1 U553 ( .A1(n734), .A2(G902), .ZN(n459) );
  XOR2_X1 U554 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n457) );
  XNOR2_X1 U555 ( .A(G902), .B(KEYINPUT15), .ZN(n632) );
  NAND2_X1 U556 ( .A1(n632), .A2(G234), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n455), .B(KEYINPUT20), .ZN(n460) );
  NAND2_X1 U558 ( .A1(n460), .A2(G217), .ZN(n456) );
  XNOR2_X1 U559 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U560 ( .A(n459), .B(n458), .ZN(n596) );
  NAND2_X1 U561 ( .A1(n460), .A2(G221), .ZN(n462) );
  XOR2_X1 U562 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n461) );
  XNOR2_X1 U563 ( .A(n462), .B(n461), .ZN(n688) );
  INV_X1 U564 ( .A(n688), .ZN(n463) );
  NAND2_X1 U565 ( .A1(n464), .A2(n463), .ZN(n538) );
  XNOR2_X1 U566 ( .A(n465), .B(KEYINPUT14), .ZN(n469) );
  NAND2_X1 U567 ( .A1(G902), .A2(n469), .ZN(n544) );
  NOR2_X1 U568 ( .A1(n484), .A2(n544), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n466), .B(KEYINPUT103), .ZN(n467) );
  NOR2_X1 U570 ( .A1(G900), .A2(n467), .ZN(n468) );
  NAND2_X1 U571 ( .A1(G952), .A2(n469), .ZN(n716) );
  NOR2_X1 U572 ( .A1(G953), .A2(n716), .ZN(n549) );
  INV_X1 U573 ( .A(n549), .ZN(n470) );
  NAND2_X1 U574 ( .A1(n427), .A2(n470), .ZN(n531) );
  INV_X1 U575 ( .A(n531), .ZN(n471) );
  NOR2_X1 U576 ( .A1(n538), .A2(n471), .ZN(n483) );
  XNOR2_X1 U577 ( .A(n473), .B(n472), .ZN(n477) );
  NAND2_X1 U578 ( .A1(n484), .A2(G227), .ZN(n475) );
  XNOR2_X1 U579 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U580 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U581 ( .A(n358), .B(n478), .ZN(n657) );
  XOR2_X1 U582 ( .A(KEYINPUT74), .B(G469), .Z(n480) );
  XNOR2_X2 U583 ( .A(n481), .B(n480), .ZN(n594) );
  INV_X1 U584 ( .A(n594), .ZN(n482) );
  AND2_X1 U585 ( .A1(n483), .A2(n482), .ZN(n520) );
  AND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n518) );
  NAND2_X1 U587 ( .A1(n484), .A2(G224), .ZN(n485) );
  XNOR2_X1 U588 ( .A(n355), .B(n485), .ZN(n488) );
  XNOR2_X1 U589 ( .A(n498), .B(n510), .ZN(n491) );
  NAND2_X1 U590 ( .A1(n651), .A2(n632), .ZN(n493) );
  XNOR2_X2 U591 ( .A(n493), .B(n359), .ZN(n550) );
  NAND2_X1 U592 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n498), .B(KEYINPUT98), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U595 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n504), .B(n503), .ZN(n653) );
  NOR2_X1 U597 ( .A1(n653), .A2(G902), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n505), .B(G475), .ZN(n506) );
  XNOR2_X1 U599 ( .A(n506), .B(KEYINPUT13), .ZN(n525) );
  INV_X1 U600 ( .A(n525), .ZN(n557) );
  NAND2_X1 U601 ( .A1(G217), .A2(n507), .ZN(n508) );
  XNOR2_X1 U602 ( .A(n509), .B(n508), .ZN(n515) );
  XOR2_X1 U603 ( .A(KEYINPUT7), .B(n510), .Z(n513) );
  XOR2_X1 U604 ( .A(n511), .B(G134), .Z(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n729) );
  NOR2_X1 U607 ( .A1(n729), .A2(G902), .ZN(n516) );
  XNOR2_X1 U608 ( .A(G478), .B(n516), .ZN(n556) );
  NOR2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n554) );
  AND2_X1 U610 ( .A1(n620), .A2(n554), .ZN(n517) );
  NAND2_X1 U611 ( .A1(n518), .A2(n517), .ZN(n610) );
  XNOR2_X1 U612 ( .A(n610), .B(G143), .ZN(G45) );
  INV_X1 U613 ( .A(KEYINPUT38), .ZN(n519) );
  AND2_X1 U614 ( .A1(n520), .A2(n701), .ZN(n522) );
  INV_X1 U615 ( .A(n556), .ZN(n523) );
  NAND2_X1 U616 ( .A1(n557), .A2(n523), .ZN(n678) );
  OR2_X1 U617 ( .A1(n524), .A2(n678), .ZN(n637) );
  XNOR2_X1 U618 ( .A(n637), .B(G134), .ZN(G36) );
  NAND2_X1 U619 ( .A1(n525), .A2(n556), .ZN(n582) );
  INV_X1 U620 ( .A(n582), .ZN(n526) );
  INV_X1 U621 ( .A(KEYINPUT109), .ZN(n528) );
  XNOR2_X1 U622 ( .A(n528), .B(KEYINPUT40), .ZN(n529) );
  XNOR2_X1 U623 ( .A(n603), .B(G131), .ZN(G33) );
  INV_X1 U624 ( .A(n464), .ZN(n687) );
  AND2_X1 U625 ( .A1(n531), .A2(n463), .ZN(n595) );
  XNOR2_X1 U626 ( .A(n578), .B(KEYINPUT6), .ZN(n541) );
  INV_X1 U627 ( .A(n541), .ZN(n532) );
  INV_X1 U628 ( .A(KEYINPUT105), .ZN(n533) );
  INV_X1 U629 ( .A(n381), .ZN(n684) );
  XOR2_X1 U630 ( .A(G125), .B(KEYINPUT37), .Z(n537) );
  XNOR2_X1 U631 ( .A(n605), .B(n537), .ZN(G27) );
  INV_X1 U632 ( .A(n538), .ZN(n685) );
  NAND2_X1 U633 ( .A1(n539), .A2(n685), .ZN(n540) );
  XNOR2_X1 U634 ( .A(n540), .B(KEYINPUT78), .ZN(n577) );
  NOR2_X1 U635 ( .A1(n577), .A2(n541), .ZN(n543) );
  INV_X1 U636 ( .A(KEYINPUT33), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n543), .B(n542), .ZN(n682) );
  INV_X1 U638 ( .A(n544), .ZN(n546) );
  INV_X1 U639 ( .A(G953), .ZN(n545) );
  NOR2_X1 U640 ( .A1(G898), .A2(n545), .ZN(n742) );
  NAND2_X1 U641 ( .A1(n546), .A2(n742), .ZN(n547) );
  XOR2_X1 U642 ( .A(KEYINPUT90), .B(n547), .Z(n548) );
  NAND2_X1 U643 ( .A1(n682), .A2(n580), .ZN(n553) );
  XNOR2_X1 U644 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n552) );
  AND2_X1 U645 ( .A1(n766), .A2(KEYINPUT70), .ZN(n569) );
  NAND2_X1 U646 ( .A1(n557), .A2(n556), .ZN(n703) );
  NOR2_X1 U647 ( .A1(n688), .A2(n703), .ZN(n558) );
  XNOR2_X1 U648 ( .A(KEYINPUT100), .B(n558), .ZN(n559) );
  NAND2_X1 U649 ( .A1(n559), .A2(n580), .ZN(n561) );
  XNOR2_X2 U650 ( .A(n561), .B(n560), .ZN(n573) );
  INV_X1 U651 ( .A(n598), .ZN(n562) );
  NOR2_X1 U652 ( .A1(n684), .A2(n562), .ZN(n563) );
  XOR2_X1 U653 ( .A(n564), .B(KEYINPUT67), .Z(n565) );
  AND2_X1 U654 ( .A1(n541), .A2(n687), .ZN(n566) );
  NAND2_X1 U655 ( .A1(n573), .A2(n566), .ZN(n567) );
  NOR2_X1 U656 ( .A1(n567), .A2(n381), .ZN(n568) );
  XNOR2_X1 U657 ( .A(n568), .B(KEYINPUT32), .ZN(n764) );
  NAND2_X1 U658 ( .A1(n569), .A2(n572), .ZN(n570) );
  XNOR2_X1 U659 ( .A(n570), .B(KEYINPUT44), .ZN(n589) );
  NOR2_X1 U660 ( .A1(KEYINPUT70), .A2(n766), .ZN(n571) );
  NAND2_X1 U661 ( .A1(n572), .A2(n571), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n573), .A2(n541), .ZN(n574) );
  XOR2_X1 U663 ( .A(KEYINPUT87), .B(n574), .Z(n575) );
  NOR2_X1 U664 ( .A1(n687), .A2(n575), .ZN(n576) );
  NAND2_X1 U665 ( .A1(n381), .A2(n576), .ZN(n662) );
  INV_X1 U666 ( .A(n578), .ZN(n690) );
  NOR2_X1 U667 ( .A1(n577), .A2(n690), .ZN(n696) );
  NOR2_X1 U668 ( .A1(n594), .A2(n578), .ZN(n579) );
  AND2_X1 U669 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U670 ( .A1(n685), .A2(n581), .ZN(n665) );
  NAND2_X1 U671 ( .A1(n677), .A2(n665), .ZN(n583) );
  NAND2_X1 U672 ( .A1(n582), .A2(n678), .ZN(n608) );
  NAND2_X1 U673 ( .A1(n583), .A2(n608), .ZN(n584) );
  XOR2_X1 U674 ( .A(n584), .B(KEYINPUT99), .Z(n585) );
  AND2_X1 U675 ( .A1(n662), .A2(n585), .ZN(n586) );
  NAND2_X1 U676 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U677 ( .A(KEYINPUT65), .ZN(n590) );
  XNOR2_X1 U678 ( .A(n590), .B(KEYINPUT45), .ZN(n591) );
  INV_X1 U679 ( .A(n636), .ZN(n720) );
  XNOR2_X1 U680 ( .A(n594), .B(KEYINPUT108), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n596), .A2(n595), .ZN(n597) );
  OR2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U683 ( .A(n599), .B(KEYINPUT28), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n698), .A2(n607), .ZN(n602) );
  INV_X1 U685 ( .A(KEYINPUT46), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT86), .ZN(n614) );
  INV_X1 U687 ( .A(n608), .ZN(n705) );
  INV_X1 U688 ( .A(KEYINPUT83), .ZN(n609) );
  XNOR2_X1 U689 ( .A(n610), .B(n609), .ZN(n611) );
  AND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  AND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n364), .A2(n381), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT43), .ZN(n622) );
  INV_X1 U695 ( .A(n620), .ZN(n621) );
  AND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n681) );
  INV_X1 U697 ( .A(n681), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n640), .A2(n637), .ZN(n627) );
  INV_X1 U700 ( .A(KEYINPUT84), .ZN(n626) );
  XNOR2_X2 U701 ( .A(n627), .B(n626), .ZN(n719) );
  INV_X1 U702 ( .A(KEYINPUT79), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n719), .B(n628), .ZN(n629) );
  INV_X1 U704 ( .A(n632), .ZN(n630) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n631) );
  OR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n634) );
  INV_X1 U707 ( .A(KEYINPUT68), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n637), .A2(KEYINPUT2), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT82), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n636), .A2(n639), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n641), .A2(n356), .ZN(n722) );
  NAND2_X1 U713 ( .A1(n357), .A2(G472), .ZN(n645) );
  XOR2_X1 U714 ( .A(KEYINPUT62), .B(n643), .Z(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n646), .A2(n660), .ZN(n648) );
  XNOR2_X1 U717 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(G57) );
  NAND2_X1 U719 ( .A1(n732), .A2(G210), .ZN(n652) );
  XOR2_X1 U720 ( .A(KEYINPUT89), .B(KEYINPUT54), .Z(n649) );
  XNOR2_X1 U721 ( .A(n649), .B(KEYINPUT55), .ZN(n650) );
  INV_X1 U722 ( .A(n660), .ZN(n738) );
  NAND2_X1 U723 ( .A1(n357), .A2(G475), .ZN(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT117), .B(KEYINPUT59), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n733), .A2(G469), .ZN(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n661) );
  AND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(G54) );
  XNOR2_X1 U730 ( .A(G101), .B(n662), .ZN(G3) );
  NOR2_X1 U731 ( .A1(n663), .A2(n665), .ZN(n664) );
  XOR2_X1 U732 ( .A(G104), .B(n664), .Z(G6) );
  NOR2_X1 U733 ( .A1(n678), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(G107), .B(n668), .ZN(G9) );
  XOR2_X1 U737 ( .A(n669), .B(G110), .Z(G12) );
  NOR2_X1 U738 ( .A1(n678), .A2(n673), .ZN(n671) );
  XNOR2_X1 U739 ( .A(KEYINPUT29), .B(KEYINPUT110), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(G128), .B(n672), .ZN(G30) );
  NOR2_X1 U742 ( .A1(n663), .A2(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(G146), .B(KEYINPUT111), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(G48) );
  NOR2_X1 U745 ( .A1(n663), .A2(n677), .ZN(n676) );
  XOR2_X1 U746 ( .A(G113), .B(n676), .Z(G15) );
  NOR2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U748 ( .A(KEYINPUT112), .B(n679), .Z(n680) );
  XNOR2_X1 U749 ( .A(G116), .B(n680), .ZN(G18) );
  XOR2_X1 U750 ( .A(G140), .B(n681), .Z(G42) );
  BUF_X1 U751 ( .A(n682), .Z(n708) );
  NAND2_X1 U752 ( .A1(n698), .A2(n708), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n683), .B(KEYINPUT115), .ZN(n718) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT50), .ZN(n694) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U757 ( .A(KEYINPUT49), .B(n689), .Z(n691) );
  NAND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U759 ( .A(n692), .B(KEYINPUT113), .Z(n693) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(KEYINPUT51), .B(n697), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n713) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n710) );
  INV_X1 U768 ( .A(n708), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U770 ( .A(KEYINPUT114), .B(n711), .Z(n712) );
  NAND2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U772 ( .A(KEYINPUT52), .B(n714), .Z(n715) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U776 ( .A1(n721), .A2(n631), .ZN(n723) );
  NAND2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U779 ( .A(KEYINPUT116), .B(n726), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n727), .A2(G953), .ZN(n728) );
  XNOR2_X1 U781 ( .A(n728), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U782 ( .A1(n733), .A2(G478), .ZN(n730) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n738), .A2(n731), .ZN(G63) );
  NAND2_X1 U785 ( .A1(n733), .A2(G217), .ZN(n736) );
  NOR2_X1 U786 ( .A1(n738), .A2(n737), .ZN(G66) );
  BUF_X1 U787 ( .A(n739), .Z(n740) );
  XNOR2_X1 U788 ( .A(G101), .B(n740), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n741), .B(KEYINPUT122), .ZN(n743) );
  NOR2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n752) );
  XOR2_X1 U791 ( .A(KEYINPUT120), .B(KEYINPUT61), .Z(n745) );
  NAND2_X1 U792 ( .A1(G224), .A2(G953), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U794 ( .A(KEYINPUT119), .B(n746), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G898), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n748), .B(KEYINPUT121), .ZN(n750) );
  NOR2_X1 U797 ( .A1(n636), .A2(G953), .ZN(n749) );
  NOR2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U800 ( .A(KEYINPUT123), .B(n753), .ZN(G69) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT124), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n756), .B(n755), .ZN(n758) );
  XNOR2_X1 U803 ( .A(n719), .B(n758), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(n484), .ZN(n762) );
  XOR2_X1 U805 ( .A(G227), .B(n758), .Z(n759) );
  NAND2_X1 U806 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U807 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U809 ( .A(KEYINPUT125), .B(n763), .Z(G72) );
  XNOR2_X1 U810 ( .A(G119), .B(KEYINPUT127), .ZN(n765) );
  XNOR2_X1 U811 ( .A(n765), .B(n764), .ZN(G21) );
  XNOR2_X1 U812 ( .A(G122), .B(KEYINPUT126), .ZN(n767) );
  XNOR2_X1 U813 ( .A(n767), .B(n766), .ZN(G24) );
  XNOR2_X1 U814 ( .A(G137), .B(n768), .ZN(G39) );
endmodule

