//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n203));
  AND2_X1   g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR3_X1   g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT22), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT22), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT76), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n203), .B(new_n206), .C1(new_n210), .C2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n202), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n204), .A2(new_n205), .ZN(new_n219));
  OR2_X1    g018(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(G218gat), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n202), .A2(new_n217), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n203), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT80), .B1(new_n218), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n206), .B1(new_n210), .B2(new_n215), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n225), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT79), .B1(new_n224), .B2(new_n203), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n228), .B(new_n231), .C1(new_n232), .C2(new_n202), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G226gat), .ZN(new_n236));
  INV_X1    g035(.A(G233gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G176gat), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT24), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT24), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(G183gat), .A3(G190gat), .ZN(new_n251));
  AND3_X1   g050(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n249), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n239), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n258));
  OAI211_X1 g057(.A(G183gat), .B(G190gat), .C1(new_n258), .C2(KEYINPUT24), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n246), .A2(KEYINPUT68), .A3(new_n250), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT69), .B(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n259), .B(new_n260), .C1(new_n262), .C2(G190gat), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n252), .A2(new_n253), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n249), .A2(KEYINPUT25), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT67), .B(new_n239), .C1(new_n248), .C2(new_n254), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n257), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OR3_X1    g070(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n272), .B(new_n273), .C1(new_n253), .C2(new_n252), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  AND2_X1   g074(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT28), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT70), .ZN(new_n279));
  INV_X1    g078(.A(new_n277), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT27), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n280), .B1(new_n261), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT28), .B1(new_n282), .B2(new_n275), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n246), .B(new_n274), .C1(new_n279), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n238), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n238), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n271), .B2(new_n284), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n235), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n285), .A2(new_n286), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  AOI211_X1 g099(.A(KEYINPUT82), .B(new_n288), .C1(new_n271), .C2(new_n284), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n298), .B(new_n234), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT81), .B(new_n235), .C1(new_n287), .C2(new_n289), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n292), .A2(new_n296), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT83), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT30), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n292), .A2(new_n302), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n295), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(KEYINPUT83), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G134gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G127gat), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G134gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n318), .B(new_n319), .C1(KEYINPUT1), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n314), .A2(new_n316), .ZN(new_n322));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323));
  XOR2_X1   g122(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n271), .A2(new_n327), .A3(new_n284), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n271), .B2(new_n284), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT64), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT34), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n333), .B2(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n330), .B(new_n333), .C1(KEYINPUT75), .C2(new_n335), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n328), .B2(new_n329), .ZN(new_n340));
  NAND2_X1  g139(.A1(KEYINPUT73), .A2(KEYINPUT33), .ZN(new_n341));
  OR2_X1    g140(.A1(KEYINPUT73), .A2(KEYINPUT33), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(KEYINPUT32), .ZN(new_n344));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G71gat), .ZN(new_n346));
  INV_X1    g145(.A(G99gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n344), .B1(new_n343), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n339), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n343), .A2(new_n348), .ZN(new_n352));
  INV_X1    g151(.A(new_n344), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n338), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n351), .A2(new_n357), .A3(KEYINPUT93), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT93), .B1(new_n351), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n312), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT31), .B(G50gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G141gat), .ZN(new_n366));
  INV_X1    g165(.A(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G148gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G155gat), .ZN(new_n370));
  INV_X1    g169(.A(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n369), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n369), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n286), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n227), .A2(new_n381), .A3(new_n233), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n383));
  INV_X1    g182(.A(new_n202), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n229), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n202), .B(new_n206), .C1(new_n210), .C2(new_n215), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT89), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT90), .B1(new_n224), .B2(new_n202), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n224), .A2(new_n389), .A3(new_n202), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n385), .A2(new_n387), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n391), .B2(new_n286), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n382), .B1(new_n392), .B2(new_n378), .ZN(new_n393));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT88), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n394), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n218), .A2(new_n226), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n398), .B2(new_n286), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n376), .B2(new_n377), .ZN(new_n401));
  XNOR2_X1  g200(.A(G141gat), .B(G148gat), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n373), .B(new_n372), .C1(new_n402), .C2(KEYINPUT2), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n369), .A2(new_n374), .A3(new_n375), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(KEYINPUT84), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n382), .B(new_n397), .C1(new_n399), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n364), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT91), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n396), .A2(KEYINPUT91), .A3(new_n414), .A4(new_n408), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(new_n410), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n413), .A2(new_n415), .B1(new_n417), .B2(new_n363), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT35), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n403), .A2(KEYINPUT84), .A3(new_n404), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT84), .B1(new_n403), .B2(new_n404), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n326), .A3(new_n380), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n321), .A2(new_n325), .A3(new_n403), .A4(new_n404), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT4), .ZN(new_n426));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT85), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT86), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n406), .B2(new_n326), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT5), .B1(new_n433), .B2(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n430), .A3(KEYINPUT86), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G85gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT0), .B(G57gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT6), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n434), .A2(new_n430), .A3(KEYINPUT86), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n434), .B1(KEYINPUT86), .B2(new_n430), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n419), .A2(new_n420), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n360), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(KEYINPUT87), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n448), .A2(new_n443), .A3(new_n455), .A4(new_n449), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n445), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(new_n308), .A3(new_n306), .A4(new_n310), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n351), .A2(new_n357), .A3(KEYINPUT74), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT74), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n419), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT35), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT94), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(KEYINPUT35), .C1(new_n458), .C2(new_n461), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n453), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT39), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT39), .B1(new_n424), .B2(new_n426), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n428), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n433), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT39), .A3(new_n429), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n441), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n472), .A2(KEYINPUT92), .A3(new_n473), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT92), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n475), .A2(new_n476), .A3(new_n444), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n311), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n307), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n300), .A2(new_n301), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n235), .B1(new_n481), .B2(new_n287), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n287), .A2(new_n235), .A3(new_n289), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT37), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n295), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n445), .A3(new_n450), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n292), .A2(KEYINPUT37), .A3(new_n302), .A4(new_n303), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n296), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n304), .B1(new_n490), .B2(new_n486), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n478), .B(new_n419), .C1(new_n488), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n419), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n458), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n459), .A2(KEYINPUT36), .A3(new_n460), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n351), .A2(new_n357), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n492), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n466), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G183gat), .B(G211gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(new_n315), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(new_n370), .ZN(new_n503));
  NAND2_X1  g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n503), .B(new_n504), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT101), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n509), .A2(new_n510), .B1(G57gat), .B2(G64gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n510), .B2(new_n509), .ZN(new_n512));
  NAND2_X1  g311(.A1(G57gat), .A2(G64gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515));
  INV_X1    g314(.A(KEYINPUT102), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n512), .A2(new_n516), .A3(new_n515), .A4(new_n513), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT21), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT99), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(G1gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G8gat), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n528), .B(new_n531), .C1(G1gat), .C2(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT104), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n523), .A2(new_n533), .A3(KEYINPUT104), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n508), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n534), .A3(new_n507), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n522), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT103), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n537), .B2(new_n539), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n506), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n537), .A2(new_n539), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(new_n543), .A3(new_n505), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G85gat), .ZN(new_n551));
  INV_X1    g350(.A(G92gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT105), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT105), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n551), .B2(new_n552), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT105), .B(new_n559), .C1(new_n551), .C2(new_n552), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  OR2_X1    g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(G29gat), .A2(G36gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT14), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(KEYINPUT15), .B(new_n566), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n566), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n572), .B(KEYINPUT97), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(new_n569), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT17), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  AOI211_X1 g383(.A(KEYINPUT98), .B(new_n584), .C1(new_n574), .C2(new_n580), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n565), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n565), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n591), .A3(new_n588), .A4(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(new_n592), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n595), .A2(new_n598), .B1(KEYINPUT106), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(KEYINPUT106), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n593), .A2(new_n594), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n550), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n533), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n583), .B2(new_n585), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n533), .A2(new_n581), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n533), .A2(new_n581), .A3(KEYINPUT100), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT100), .B1(new_n533), .B2(new_n581), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n608), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n607), .A2(KEYINPUT18), .A3(new_n608), .A4(new_n609), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621));
  INV_X1    g420(.A(G197gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT11), .B(G169gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n612), .A2(new_n618), .A3(new_n626), .A4(new_n619), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G230gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n237), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n519), .A2(new_n520), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n563), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n565), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n587), .A2(new_n633), .A3(new_n635), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n587), .A2(new_n633), .A3(KEYINPUT10), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n632), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n632), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n637), .B2(new_n638), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n645), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n630), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n500), .A2(new_n605), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n457), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT108), .B(G1gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G8gat), .ZN(new_n658));
  OR4_X1    g457(.A1(new_n657), .A2(new_n653), .A3(new_n312), .A4(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n653), .A2(KEYINPUT109), .A3(new_n312), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT109), .B1(new_n653), .B2(new_n312), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n657), .B1(new_n662), .B2(G8gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n658), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n495), .A2(new_n667), .A3(new_n497), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n495), .B2(new_n497), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n653), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n653), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n358), .A2(new_n359), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n666), .B2(new_n676), .ZN(G1326gat));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n414), .A3(new_n493), .ZN(new_n678));
  OAI21_X1  g477(.A(G22gat), .B1(new_n653), .B2(new_n419), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(G1327gat));
  INV_X1    g481(.A(new_n603), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n550), .A2(new_n630), .A3(new_n651), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n500), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(G29gat), .A3(new_n457), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT45), .Z(new_n687));
  OAI21_X1  g486(.A(new_n683), .B1(new_n466), .B2(new_n499), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n492), .B(new_n494), .C1(new_n668), .C2(new_n669), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n690), .B(new_n683), .C1(new_n692), .C2(new_n466), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n684), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n457), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n687), .A2(new_n696), .ZN(G1328gat));
  NOR2_X1   g496(.A1(new_n685), .A2(G36gat), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT46), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n311), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n699), .A2(KEYINPUT46), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n695), .A2(KEYINPUT113), .A3(new_n312), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT113), .B1(new_n695), .B2(new_n312), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(G36gat), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(G1329gat));
  NAND2_X1  g506(.A1(new_n670), .A2(G43gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n685), .A2(new_n674), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n695), .A2(new_n708), .B1(new_n709), .B2(G43gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g510(.A1(new_n493), .A2(G50gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n685), .A2(new_n419), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n695), .A2(new_n712), .B1(new_n713), .B2(G50gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g514(.A1(new_n628), .A2(new_n629), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n463), .A2(new_n465), .ZN(new_n717));
  INV_X1    g516(.A(new_n453), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(new_n691), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n604), .A2(new_n650), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n457), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n722), .A2(KEYINPUT114), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n720), .A2(new_n728), .A3(new_n721), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n731));
  INV_X1    g530(.A(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n311), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT115), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n732), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n738), .A3(new_n675), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n671), .B1(new_n727), .B2(new_n729), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n738), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n742), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n744), .B(new_n739), .C1(new_n740), .C2(new_n738), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n493), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n550), .A2(new_n716), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n694), .A2(new_n651), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n457), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n724), .A2(new_n651), .A3(new_n551), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT117), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n603), .B1(new_n719), .B2(new_n691), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n754), .B2(new_n749), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n683), .B(new_n749), .C1(new_n692), .C2(new_n466), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n751), .A2(new_n759), .ZN(G1336gat));
  OAI21_X1  g559(.A(G92gat), .B1(new_n750), .B2(new_n312), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n312), .A2(G92gat), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n651), .B(new_n762), .C1(new_n755), .C2(new_n758), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n766), .A3(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1337gat));
  NOR3_X1   g567(.A1(new_n750), .A2(new_n347), .A3(new_n671), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n675), .B(new_n651), .C1(new_n755), .C2(new_n758), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n347), .B2(new_n770), .ZN(G1338gat));
  NOR2_X1   g570(.A1(new_n419), .A2(G106gat), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n651), .B(new_n772), .C1(new_n755), .C2(new_n758), .ZN(new_n773));
  INV_X1    g572(.A(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n749), .A2(new_n651), .ZN(new_n775));
  AOI211_X1 g574(.A(new_n419), .B(new_n775), .C1(new_n689), .C2(new_n693), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n774), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  OAI221_X1 g580(.A(new_n773), .B1(new_n779), .B2(KEYINPUT53), .C1(new_n774), .C2(new_n776), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(G1339gat));
  NAND2_X1  g582(.A1(new_n630), .A2(new_n650), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n604), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n640), .A2(KEYINPUT119), .A3(new_n632), .A4(new_n641), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n642), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n640), .A2(new_n641), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n643), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT54), .B(new_n786), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n649), .B1(new_n642), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n645), .A2(new_n648), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n615), .A2(new_n617), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n625), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n629), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n791), .A2(new_n793), .A3(KEYINPUT55), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n796), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n550), .B1(new_n803), .B2(new_n683), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n796), .A2(new_n716), .A3(new_n797), .A4(new_n802), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n651), .A2(new_n801), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n603), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n785), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n457), .A3(new_n493), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n459), .A2(new_n460), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n312), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT120), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(KEYINPUT120), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n630), .A2(G113gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n809), .A2(new_n312), .A3(new_n675), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n630), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1340gat));
  NOR2_X1   g618(.A1(new_n650), .A2(G120gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n813), .A2(new_n814), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n817), .B2(new_n650), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  INV_X1    g622(.A(new_n550), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n817), .A2(new_n315), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n812), .A2(new_n550), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n315), .ZN(G1342gat));
  NOR2_X1   g626(.A1(new_n603), .A2(new_n311), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT121), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n811), .A2(new_n313), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n817), .B2(new_n603), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n831), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(G1343gat));
  NAND3_X1  g634(.A1(new_n671), .A2(new_n724), .A3(new_n312), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n808), .A2(new_n419), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n716), .A2(new_n367), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(KEYINPUT124), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(KEYINPUT124), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n804), .A2(new_n807), .ZN(new_n845));
  INV_X1    g644(.A(new_n785), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n493), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n808), .A2(KEYINPUT57), .A3(new_n419), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n670), .A2(new_n457), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(KEYINPUT122), .A3(new_n312), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n850), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n716), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n843), .B1(new_n859), .B2(G141gat), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n850), .A2(new_n855), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n630), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n367), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n843), .A2(KEYINPUT58), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n860), .A2(new_n861), .B1(new_n864), .B2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(new_n839), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n365), .A3(new_n651), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT59), .B(G148gat), .C1(new_n862), .C2(new_n650), .ZN(new_n869));
  INV_X1    g668(.A(new_n858), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n365), .B1(new_n872), .B2(new_n651), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n868), .B(new_n869), .C1(new_n873), .C2(KEYINPUT59), .ZN(G1345gat));
  NAND3_X1  g673(.A1(new_n867), .A2(new_n370), .A3(new_n550), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n824), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n370), .ZN(G1346gat));
  NAND4_X1  g676(.A1(new_n838), .A2(new_n371), .A3(new_n853), .A4(new_n829), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n603), .B1(new_n870), .B2(new_n871), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n371), .ZN(G1347gat));
  NOR4_X1   g679(.A1(new_n808), .A2(new_n724), .A3(new_n312), .A4(new_n493), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n675), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n630), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n881), .A2(new_n810), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT125), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n881), .A2(new_n889), .A3(new_n810), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n716), .B1(new_n243), .B2(new_n242), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n885), .A2(new_n886), .B1(new_n891), .B2(new_n892), .ZN(G1348gat));
  INV_X1    g692(.A(G176gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n882), .A2(new_n894), .A3(new_n650), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n888), .A2(new_n651), .A3(new_n890), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n894), .ZN(G1349gat));
  OAI21_X1  g696(.A(new_n262), .B1(new_n882), .B2(new_n824), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n550), .B1(new_n277), .B2(new_n276), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g700(.A1(new_n888), .A2(new_n275), .A3(new_n683), .A4(new_n890), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n881), .A2(new_n683), .A3(new_n675), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(G190gat), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(new_n903), .A3(G190gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n670), .A2(new_n724), .A3(new_n312), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n850), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n630), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n838), .A2(new_n910), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n622), .A3(new_n716), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1352gat));
  INV_X1    g714(.A(G204gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n916), .A3(new_n651), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT62), .Z(new_n918));
  OAI21_X1  g717(.A(G204gat), .B1(new_n911), .B2(new_n650), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1353gat));
  OAI211_X1 g719(.A(new_n913), .B(new_n550), .C1(new_n208), .C2(new_n207), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n850), .A2(new_n550), .A3(new_n910), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n911), .B2(new_n603), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n913), .A2(new_n209), .A3(new_n683), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1355gat));
endmodule


