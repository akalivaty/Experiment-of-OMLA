

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XOR2_X1 U325 ( .A(G155GAT), .B(KEYINPUT3), .Z(n293) );
  XOR2_X1 U326 ( .A(n419), .B(n418), .Z(n294) );
  XNOR2_X1 U327 ( .A(KEYINPUT113), .B(KEYINPUT45), .ZN(n390) );
  XNOR2_X1 U328 ( .A(n391), .B(n390), .ZN(n392) );
  INV_X1 U329 ( .A(G106GAT), .ZN(n301) );
  XNOR2_X1 U330 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U331 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U332 ( .A(n426), .B(n425), .ZN(n429) );
  INV_X1 U333 ( .A(n521), .ZN(n467) );
  XNOR2_X1 U334 ( .A(n359), .B(n303), .ZN(n304) );
  XNOR2_X1 U335 ( .A(n432), .B(KEYINPUT55), .ZN(n451) );
  XOR2_X1 U336 ( .A(n312), .B(n311), .Z(n559) );
  XOR2_X1 U337 ( .A(KEYINPUT38), .B(n496), .Z(n504) );
  XNOR2_X1 U338 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U339 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n296) );
  XNOR2_X1 U341 ( .A(KEYINPUT66), .B(KEYINPUT78), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n312) );
  XOR2_X1 U343 ( .A(G99GAT), .B(G85GAT), .Z(n369) );
  XOR2_X1 U344 ( .A(KEYINPUT64), .B(n369), .Z(n298) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(n397), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n305) );
  XOR2_X1 U348 ( .A(G29GAT), .B(G43GAT), .Z(n300) );
  XNOR2_X1 U349 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n359) );
  NAND2_X1 U351 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U352 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U353 ( .A(G50GAT), .B(G162GAT), .Z(n418) );
  XOR2_X1 U354 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n307) );
  XNOR2_X1 U355 ( .A(G134GAT), .B(G92GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n418), .B(n308), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(G57GAT), .B(KEYINPUT1), .Z(n314) );
  XNOR2_X1 U360 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n334) );
  XOR2_X1 U362 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n316) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U365 ( .A(KEYINPUT87), .B(KEYINPUT91), .Z(n318) );
  XNOR2_X1 U366 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n332) );
  XNOR2_X1 U369 ( .A(KEYINPUT86), .B(KEYINPUT2), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n293), .B(n321), .ZN(n419) );
  XOR2_X1 U371 ( .A(G134GAT), .B(KEYINPUT0), .Z(n433) );
  XOR2_X1 U372 ( .A(n419), .B(n433), .Z(n323) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n330) );
  XOR2_X1 U375 ( .A(G85GAT), .B(G162GAT), .Z(n325) );
  XNOR2_X1 U376 ( .A(G127GAT), .B(G148GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(n326), .B(G120GAT), .Z(n328) );
  XOR2_X1 U379 ( .A(G113GAT), .B(G1GAT), .Z(n353) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n353), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(n334), .B(n333), .Z(n521) );
  XOR2_X1 U385 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n336) );
  XNOR2_X1 U386 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT13), .Z(n368) );
  XOR2_X1 U389 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XOR2_X1 U390 ( .A(n368), .B(n434), .Z(n338) );
  XNOR2_X1 U391 ( .A(G183GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U393 ( .A(n340), .B(n339), .Z(n342) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n350) );
  XOR2_X1 U396 ( .A(G155GAT), .B(G78GAT), .Z(n344) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G211GAT), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT80), .B(G64GAT), .Z(n346) );
  XNOR2_X1 U400 ( .A(G1GAT), .B(G8GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(n348), .B(n347), .Z(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n581) );
  XOR2_X1 U404 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n352) );
  XNOR2_X1 U405 ( .A(G15GAT), .B(G197GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n367) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G50GAT), .Z(n355) );
  XOR2_X1 U408 ( .A(G169GAT), .B(G8GAT), .Z(n402) );
  XNOR2_X1 U409 ( .A(n353), .B(n402), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XOR2_X1 U412 ( .A(n356), .B(n427), .Z(n365) );
  XOR2_X1 U413 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n358) );
  XNOR2_X1 U414 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U416 ( .A(n359), .B(KEYINPUT70), .Z(n361) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n561) );
  XOR2_X1 U422 ( .A(KEYINPUT75), .B(n368), .Z(n371) );
  XNOR2_X1 U423 ( .A(G204GAT), .B(n369), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U425 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n373) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U428 ( .A(n375), .B(n374), .Z(n377) );
  XOR2_X1 U429 ( .A(G120GAT), .B(G71GAT), .Z(n447) );
  XNOR2_X1 U430 ( .A(n447), .B(KEYINPUT73), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U432 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT76), .B(KEYINPUT74), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(n381), .B(n380), .Z(n385) );
  XNOR2_X1 U436 ( .A(G106GAT), .B(G78GAT), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n382), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U438 ( .A(G176GAT), .B(G92GAT), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n383), .B(G64GAT), .ZN(n398) );
  XNOR2_X1 U440 ( .A(n422), .B(n398), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n578) );
  XNOR2_X1 U442 ( .A(n578), .B(KEYINPUT41), .ZN(n565) );
  NOR2_X1 U443 ( .A1(n561), .A2(n565), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n386), .B(KEYINPUT46), .ZN(n387) );
  NOR2_X1 U445 ( .A1(n581), .A2(n387), .ZN(n388) );
  NAND2_X1 U446 ( .A1(n559), .A2(n388), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(KEYINPUT47), .ZN(n395) );
  INV_X1 U448 ( .A(n559), .ZN(n542) );
  XNOR2_X1 U449 ( .A(KEYINPUT36), .B(n542), .ZN(n586) );
  NAND2_X1 U450 ( .A1(n581), .A2(n586), .ZN(n391) );
  NAND2_X1 U451 ( .A1(n392), .A2(n561), .ZN(n393) );
  NOR2_X1 U452 ( .A1(n393), .A2(n578), .ZN(n394) );
  NOR2_X1 U453 ( .A1(n395), .A2(n394), .ZN(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT48), .B(n396), .Z(n529) );
  XOR2_X1 U455 ( .A(n398), .B(n397), .Z(n404) );
  XOR2_X1 U456 ( .A(KEYINPUT17), .B(KEYINPUT82), .Z(n400) );
  XNOR2_X1 U457 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U459 ( .A(KEYINPUT19), .B(n401), .Z(n437) );
  XNOR2_X1 U460 ( .A(n402), .B(n437), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n406) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U465 ( .A(n408), .B(n407), .Z(n415) );
  XOR2_X1 U466 ( .A(KEYINPUT21), .B(G204GAT), .Z(n410) );
  XNOR2_X1 U467 ( .A(G197GAT), .B(G211GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U469 ( .A(G218GAT), .B(KEYINPUT85), .Z(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n430) );
  INV_X1 U471 ( .A(n430), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n413), .B(KEYINPUT95), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n485) );
  INV_X1 U474 ( .A(n485), .ZN(n523) );
  AND2_X1 U475 ( .A1(n529), .A2(n523), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n416), .B(KEYINPUT54), .ZN(n417) );
  AND2_X1 U477 ( .A1(n467), .A2(n417), .ZN(n572) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n294), .B(n420), .ZN(n421) );
  XOR2_X1 U480 ( .A(n421), .B(KEYINPUT84), .Z(n426) );
  XNOR2_X1 U481 ( .A(n422), .B(KEYINPUT23), .ZN(n424) );
  INV_X1 U482 ( .A(KEYINPUT22), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n427), .B(KEYINPUT24), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n460) );
  NAND2_X1 U486 ( .A1(n572), .A2(n460), .ZN(n432) );
  XOR2_X1 U487 ( .A(G190GAT), .B(G99GAT), .Z(n436) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U491 ( .A(G43GAT), .B(G113GAT), .Z(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U493 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n442) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n450) );
  XOR2_X1 U497 ( .A(KEYINPUT65), .B(KEYINPUT81), .Z(n446) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(G176GAT), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n488) );
  INV_X1 U502 ( .A(n488), .ZN(n532) );
  NAND2_X1 U503 ( .A1(n451), .A2(n532), .ZN(n568) );
  NOR2_X1 U504 ( .A1(n559), .A2(n568), .ZN(n455) );
  XNOR2_X1 U505 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n453) );
  INV_X1 U506 ( .A(G190GAT), .ZN(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n477) );
  XNOR2_X1 U508 ( .A(n460), .B(KEYINPUT28), .ZN(n531) );
  INV_X1 U509 ( .A(n531), .ZN(n515) );
  INV_X1 U510 ( .A(n561), .ZN(n574) );
  NOR2_X1 U511 ( .A1(n574), .A2(n565), .ZN(n508) );
  NOR2_X1 U512 ( .A1(n485), .A2(n488), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT97), .B(n456), .ZN(n457) );
  NAND2_X1 U514 ( .A1(n457), .A2(n460), .ZN(n458) );
  XNOR2_X1 U515 ( .A(KEYINPUT25), .B(n458), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT98), .ZN(n465) );
  XNOR2_X1 U517 ( .A(n485), .B(KEYINPUT27), .ZN(n469) );
  INV_X1 U518 ( .A(KEYINPUT26), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n532), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT96), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n463), .B(n462), .ZN(n547) );
  NOR2_X1 U522 ( .A1(n469), .A2(n547), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT99), .ZN(n468) );
  AND2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n467), .A2(n469), .ZN(n528) );
  NAND2_X1 U527 ( .A1(n528), .A2(n531), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n532), .A2(n470), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n481) );
  NOR2_X1 U530 ( .A1(n481), .A2(n581), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n473), .A2(n586), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT37), .ZN(n494) );
  NAND2_X1 U533 ( .A1(n508), .A2(n494), .ZN(n475) );
  XOR2_X1 U534 ( .A(KEYINPUT110), .B(n475), .Z(n525) );
  NAND2_X1 U535 ( .A1(n515), .A2(n525), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n301), .B(n478), .ZN(G1339GAT) );
  NOR2_X1 U538 ( .A1(n578), .A2(n561), .ZN(n495) );
  INV_X1 U539 ( .A(n581), .ZN(n569) );
  NOR2_X1 U540 ( .A1(n569), .A2(n542), .ZN(n479) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U542 ( .A1(n481), .A2(n480), .ZN(n507) );
  NAND2_X1 U543 ( .A1(n495), .A2(n507), .ZN(n491) );
  NOR2_X1 U544 ( .A1(n467), .A2(n491), .ZN(n483) );
  XNOR2_X1 U545 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n484), .Z(G1324GAT) );
  NOR2_X1 U548 ( .A1(n485), .A2(n491), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U551 ( .A1(n488), .A2(n491), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n531), .A2(n491), .ZN(n492) );
  XOR2_X1 U555 ( .A(KEYINPUT102), .B(n492), .Z(n493) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U558 ( .A1(n495), .A2(n494), .ZN(n496) );
  NAND2_X1 U559 ( .A1(n521), .A2(n504), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XOR2_X1 U561 ( .A(G36GAT), .B(KEYINPUT103), .Z(n500) );
  NAND2_X1 U562 ( .A1(n504), .A2(n523), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n502) );
  NAND2_X1 U565 ( .A1(n532), .A2(n504), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U567 ( .A(G43GAT), .B(n503), .Z(G1330GAT) );
  XOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U569 ( .A1(n515), .A2(n504), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n511) );
  NAND2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT107), .B(n509), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n516), .A2(n521), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  NAND2_X1 U577 ( .A1(n523), .A2(n516), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n532), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT108), .Z(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n521), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT111), .Z(n527) );
  NAND2_X1 U591 ( .A1(n532), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(KEYINPUT114), .B(n530), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U596 ( .A1(n548), .A2(n533), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n543), .A2(n574), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n537) );
  INV_X1 U600 ( .A(n565), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n543), .A2(n535), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U605 ( .A1(n543), .A2(n581), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(n549), .Z(n558) );
  NOR2_X1 U614 ( .A1(n558), .A2(n561), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U617 ( .A1(n558), .A2(n565), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n569), .A2(n558), .ZN(n557) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n568), .ZN(n562) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n562), .Z(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n565), .A2(n568), .ZN(n566) );
  XOR2_X1 U633 ( .A(n567), .B(n566), .Z(G1349GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  INV_X1 U637 ( .A(n572), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n573), .A2(n547), .ZN(n587) );
  AND2_X1 U639 ( .A1(n574), .A2(n587), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n584) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT125), .B(n585), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(G1355GAT) );
endmodule

