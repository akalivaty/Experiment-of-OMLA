//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(G237), .A2(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G143), .A3(G214), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G131), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n195), .B2(G131), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT17), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT83), .ZN(new_n202));
  INV_X1    g016(.A(new_n195), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(new_n205), .A3(new_n206), .A4(new_n197), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  INV_X1    g025(.A(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G125), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT73), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n212), .A2(KEYINPUT73), .A3(G125), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n208), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n212), .A2(KEYINPUT73), .A3(G125), .ZN(new_n220));
  XNOR2_X1  g034(.A(G125), .B(G140), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(KEYINPUT73), .ZN(new_n222));
  OAI211_X1 g036(.A(G146), .B(new_n219), .C1(new_n222), .C2(new_n209), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n218), .A2(new_n223), .A3(KEYINPUT84), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT84), .B1(new_n218), .B2(new_n223), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n200), .B(new_n207), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n208), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n221), .A2(KEYINPUT75), .A3(new_n208), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n222), .A2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT18), .A2(G131), .ZN(new_n237));
  XOR2_X1   g051(.A(new_n237), .B(KEYINPUT82), .Z(new_n238));
  NAND2_X1  g052(.A1(new_n203), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n195), .B(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n236), .B(new_n239), .C1(new_n241), .C2(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(new_n229), .A3(new_n242), .ZN(new_n243));
  MUX2_X1   g057(.A(new_n221), .B(new_n222), .S(KEYINPUT19), .Z(new_n244));
  OAI21_X1  g058(.A(new_n223), .B1(new_n244), .B2(G146), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n202), .A2(new_n205), .A3(new_n197), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n229), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G475), .A2(G902), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n187), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n251), .ZN(new_n253));
  AOI211_X1 g067(.A(KEYINPUT20), .B(new_n253), .C1(new_n243), .C2(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n226), .A2(new_n242), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n248), .ZN(new_n256));
  AOI21_X1  g070(.A(G902), .B1(new_n256), .B2(new_n243), .ZN(new_n257));
  INV_X1    g071(.A(G475), .ZN(new_n258));
  OAI22_X1  g072(.A1(new_n252), .A2(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI221_X1 g075(.A(KEYINPUT85), .B1(new_n257), .B2(new_n258), .C1(new_n252), .C2(new_n254), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT9), .B(G234), .ZN(new_n264));
  OAI21_X1  g078(.A(G221), .B1(new_n264), .B2(G902), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G469), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  INV_X1    g086(.A(KEYINPUT10), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n208), .A2(G143), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G128), .ZN(new_n277));
  INV_X1    g091(.A(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n208), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n191), .A2(G146), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n276), .A2(new_n284), .A3(new_n279), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n277), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G101), .ZN(new_n287));
  INV_X1    g101(.A(G107), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G104), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n228), .A2(G107), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT77), .B1(new_n288), .B2(G104), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n228), .A3(G107), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n288), .A3(G104), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n292), .B1(new_n299), .B2(G101), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n273), .B1(new_n286), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT78), .B(new_n273), .C1(new_n286), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n299), .A2(new_n306), .A3(G101), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT4), .B1(new_n299), .B2(G101), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n299), .A2(G101), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n280), .A2(new_n281), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT0), .A2(G128), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT0), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(new_n278), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n280), .B(new_n281), .C1(new_n314), .C2(new_n278), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT70), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n315), .A2(new_n313), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n317), .B(KEYINPUT70), .C1(new_n320), .C2(new_n276), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n283), .A2(new_n285), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n312), .A2(new_n278), .B1(KEYINPUT1), .B2(new_n274), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n300), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n311), .A2(new_n322), .B1(new_n325), .B2(KEYINPUT10), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n305), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  INV_X1    g143(.A(G134), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G137), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(KEYINPUT11), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(G134), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT11), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT65), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(KEYINPUT65), .B(new_n334), .C1(new_n330), .C2(G137), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n332), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT66), .A2(G131), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n330), .A2(G137), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n333), .B2(new_n334), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT65), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n331), .B2(KEYINPUT11), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n345), .B2(new_n336), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n339), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n327), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n305), .A2(new_n326), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n272), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AND4_X1   g166(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n298), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n291), .B1(new_n353), .B2(new_n287), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n284), .B1(new_n276), .B2(new_n279), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n284), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n324), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n348), .B1(new_n358), .B2(new_n325), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT12), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT12), .B(new_n348), .C1(new_n358), .C2(new_n325), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n363), .A2(new_n351), .A3(new_n272), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n267), .B(new_n268), .C1(new_n352), .C2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n267), .A2(new_n268), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n351), .ZN(new_n369));
  INV_X1    g183(.A(new_n272), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n349), .A2(new_n351), .A3(new_n272), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT79), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(G469), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n266), .B1(new_n368), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n191), .A2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n278), .A2(G143), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(new_n330), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G122), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(G122), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(KEYINPUT14), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(KEYINPUT14), .B2(new_n384), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  XNOR2_X1  g202(.A(G116), .B(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n288), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n379), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(KEYINPUT13), .B2(new_n380), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(G134), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n381), .A2(new_n330), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n389), .B(new_n288), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n264), .A2(new_n400), .A3(G953), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n391), .A2(new_n398), .A3(new_n401), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  AOI211_X1 g225(.A(G953), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT21), .B(G898), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT87), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n268), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G214), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n420));
  INV_X1    g234(.A(G119), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(G116), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n383), .A2(KEYINPUT69), .A3(G119), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(KEYINPUT68), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G119), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n427), .A3(G116), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT2), .B(G113), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n430), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n424), .A3(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n299), .A2(new_n306), .A3(G101), .ZN(new_n435));
  INV_X1    g249(.A(new_n310), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n435), .C1(new_n436), .C2(new_n308), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT68), .B(G119), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(G116), .ZN(new_n440));
  OAI211_X1 g254(.A(G113), .B(new_n440), .C1(new_n429), .C2(new_n439), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n354), .A3(new_n433), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G122), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n443), .B(KEYINPUT8), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n433), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n300), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n447), .B2(new_n442), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n286), .A2(new_n210), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n316), .A2(G125), .A3(new_n317), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT80), .A2(KEYINPUT7), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G224), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G953), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n453), .B(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n449), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n435), .B1(new_n436), .B2(new_n308), .ZN(new_n461));
  INV_X1    g275(.A(new_n434), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n442), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n443), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n468), .A3(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n450), .A2(new_n451), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n455), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n459), .A2(new_n460), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n460), .B1(new_n459), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n419), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND4_X1   g290(.A1(new_n263), .A2(new_n378), .A3(new_n418), .A4(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n340), .B(new_n343), .C1(new_n345), .C2(new_n336), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n345), .A2(new_n336), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n339), .B1(new_n479), .B2(new_n332), .ZN(new_n480));
  INV_X1    g294(.A(new_n321), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n478), .A2(new_n480), .B1(new_n481), .B2(new_n318), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n346), .A2(new_n204), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n204), .B1(new_n333), .B2(new_n342), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n357), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n462), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n316), .A2(new_n317), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n348), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n462), .B1(new_n490), .B2(new_n486), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT28), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n487), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n193), .A2(G210), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT27), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT71), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT26), .B(G101), .Z(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n482), .A2(new_n486), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n434), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n493), .B1(new_n507), .B2(new_n487), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n499), .B(new_n504), .C1(new_n509), .C2(new_n496), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n482), .A2(KEYINPUT30), .A3(new_n486), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n484), .B1(new_n323), .B2(new_n324), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n348), .A2(new_n489), .B1(new_n512), .B2(new_n483), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n511), .B(new_n434), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n487), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(new_n504), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n517), .B2(new_n496), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G472), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT32), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n487), .A3(new_n504), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n515), .A2(KEYINPUT31), .A3(new_n487), .A4(new_n504), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n527));
  INV_X1    g341(.A(new_n504), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G902), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G472), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n521), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n533));
  NOR4_X1   g347(.A1(new_n533), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n520), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n218), .A2(new_n223), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n421), .A2(new_n278), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n438), .B2(new_n278), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT24), .B(G110), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n425), .A2(new_n427), .A3(new_n543), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n278), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G110), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n537), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G110), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n544), .A2(new_n550), .A3(new_n545), .A4(new_n546), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n538), .B(new_n540), .C1(new_n438), .C2(new_n278), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT74), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n223), .A3(new_n234), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n549), .B2(new_n557), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n536), .B(new_n268), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n400), .B1(G234), .B2(new_n268), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n549), .A2(new_n557), .ZN(new_n569));
  INV_X1    g383(.A(new_n562), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n563), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n536), .B1(new_n572), .B2(new_n268), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n567), .A2(G902), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n535), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n477), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT88), .B(G101), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G3));
  NAND2_X1  g394(.A1(new_n526), .A2(new_n529), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n531), .A3(new_n268), .ZN(new_n582));
  OAI21_X1  g396(.A(G472), .B1(new_n533), .B2(G902), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n378), .A2(new_n584), .A3(new_n576), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n261), .A2(new_n262), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n405), .A2(new_n408), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n403), .B2(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n403), .A2(new_n404), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n587), .B1(new_n593), .B2(new_n408), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n586), .A2(KEYINPUT91), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT89), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n602), .B(new_n419), .C1(new_n473), .C2(new_n474), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n417), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT92), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT91), .B1(new_n586), .B2(new_n595), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n597), .B(new_n594), .C1(new_n261), .C2(new_n262), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n604), .B(KEYINPUT92), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n585), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(new_n252), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n250), .A2(new_n187), .A3(new_n251), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT93), .B1(new_n252), .B2(new_n254), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT94), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n257), .B2(new_n258), .ZN(new_n620));
  INV_X1    g434(.A(new_n243), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n229), .B1(new_n226), .B2(new_n242), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n268), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(KEYINPUT94), .A3(G475), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n620), .A2(new_n624), .A3(new_n410), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n604), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n585), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT95), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT35), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT96), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n569), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n575), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n568), .B2(new_n573), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(KEYINPUT97), .B(new_n635), .C1(new_n568), .C2(new_n573), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n584), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n477), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n601), .B2(new_n603), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n412), .B(KEYINPUT98), .Z(new_n646));
  INV_X1    g460(.A(new_n416), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(G900), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n618), .A2(new_n625), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n535), .A2(new_n645), .A3(new_n378), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  AND3_X1   g466(.A1(new_n375), .A2(G469), .A3(new_n376), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n365), .A2(new_n367), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n265), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n656));
  XOR2_X1   g470(.A(new_n648), .B(new_n656), .Z(new_n657));
  OR2_X1    g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n530), .A2(new_n521), .A3(new_n531), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n522), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n504), .B1(new_n487), .B2(new_n507), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n268), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT100), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g481(.A(KEYINPUT100), .B(new_n666), .C1(new_n532), .C2(new_n534), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n473), .A2(new_n474), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n410), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n261), .B2(new_n262), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n419), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n675), .A2(new_n678), .A3(new_n679), .A4(new_n636), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n659), .A2(new_n671), .A3(new_n672), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  AOI211_X1 g496(.A(new_n594), .B(new_n649), .C1(new_n261), .C2(new_n262), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n535), .A3(new_n645), .A4(new_n378), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  NAND2_X1  g499(.A1(new_n535), .A2(new_n576), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n268), .B1(new_n352), .B2(new_n364), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(KEYINPUT102), .A3(new_n365), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n690), .A3(G469), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n265), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n605), .B2(new_n609), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  AOI21_X1  g511(.A(new_n266), .B1(new_n689), .B2(new_n691), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n577), .A2(new_n627), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AND3_X1   g514(.A1(new_n698), .A2(new_n263), .A3(new_n418), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n535), .A2(new_n645), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT103), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n698), .A2(new_n263), .A3(new_n418), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n535), .A2(new_n645), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NOR2_X1   g523(.A1(new_n693), .A2(new_n417), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n601), .A2(new_n603), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n678), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n526), .B1(new_n509), .B2(new_n504), .ZN(new_n713));
  NOR2_X1   g527(.A1(G472), .A2(G902), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n715), .A2(new_n576), .A3(new_n583), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  NAND2_X1  g532(.A1(new_n601), .A2(new_n603), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n715), .A2(new_n583), .A3(new_n636), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n683), .A2(new_n719), .A3(new_n698), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n673), .A2(new_n679), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n371), .A2(new_n372), .A3(G469), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n365), .A2(new_n367), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(new_n729), .A3(new_n265), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n729), .B1(new_n728), .B2(new_n265), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n726), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(KEYINPUT105), .B(new_n726), .C1(new_n730), .C2(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n725), .A2(new_n736), .A3(new_n577), .A4(new_n683), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n686), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n725), .B1(new_n738), .B2(new_n683), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n723), .B(new_n724), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n728), .A2(new_n265), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n728), .A2(new_n729), .A3(new_n265), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT105), .B1(new_n744), .B2(new_n726), .ZN(new_n745));
  INV_X1    g559(.A(new_n735), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n577), .B(new_n683), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n738), .A2(new_n725), .A3(new_n683), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT42), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n586), .A2(new_n595), .A3(new_n648), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n686), .B(new_n751), .C1(new_n734), .C2(new_n735), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT107), .B1(new_n752), .B2(KEYINPUT42), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n740), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  XNOR2_X1  g569(.A(new_n650), .B(KEYINPUT108), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n756), .B(new_n577), .C1(new_n745), .C2(new_n746), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  OAI21_X1  g573(.A(G469), .B1(new_n373), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n375), .A2(new_n376), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n759), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n366), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n365), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n265), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(new_n657), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n263), .A2(new_n595), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT110), .B1(new_n770), .B2(KEYINPUT109), .ZN(new_n773));
  MUX2_X1   g587(.A(new_n772), .B(KEYINPUT43), .S(new_n773), .Z(new_n774));
  INV_X1    g588(.A(new_n636), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n584), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(KEYINPUT44), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n769), .A2(new_n726), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT44), .B1(new_n774), .B2(new_n776), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n767), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n766), .A2(KEYINPUT47), .A3(new_n265), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n726), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n535), .A2(new_n751), .A3(new_n786), .A4(new_n576), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT111), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND3_X1  g604(.A1(new_n576), .A2(new_n265), .A3(new_n419), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT112), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n770), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT113), .Z(new_n794));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n692), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT114), .Z(new_n797));
  OAI21_X1  g611(.A(new_n675), .B1(new_n692), .B2(new_n795), .ZN(new_n798));
  OR4_X1    g612(.A1(new_n671), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n596), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n475), .A2(new_n417), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n586), .A2(new_n676), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n803), .A2(new_n804), .A3(new_n801), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n804), .B1(new_n803), .B2(new_n801), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n807), .A2(new_n585), .B1(new_n703), .B2(new_n707), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n477), .B1(new_n577), .B2(new_n640), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n699), .A3(new_n717), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n810), .A3(new_n695), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n683), .B(new_n720), .C1(new_n745), .C2(new_n746), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n786), .A2(new_n644), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n676), .A2(new_n620), .A3(new_n624), .A4(new_n648), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n618), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n813), .A2(new_n535), .A3(new_n378), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n757), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n684), .A2(new_n721), .A3(new_n651), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n728), .A2(new_n265), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n648), .B(KEYINPUT116), .Z(new_n822));
  NAND2_X1  g636(.A1(new_n775), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n719), .A2(new_n677), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n666), .B1(new_n532), .B2(new_n534), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n828), .B2(new_n668), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n819), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n751), .A2(new_n655), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n650), .A2(new_n378), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n702), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n719), .A2(new_n677), .A3(new_n821), .A4(new_n824), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n667), .B2(new_n669), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT52), .A4(new_n721), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n754), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT119), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n757), .A2(new_n812), .A3(new_n816), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n695), .A3(new_n810), .A4(new_n808), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n724), .B1(new_n737), .B2(new_n739), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n723), .B1(new_n747), .B2(new_n724), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n844), .B2(new_n740), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT53), .A4(new_n837), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n837), .A2(KEYINPUT117), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n830), .A2(new_n836), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n748), .A2(new_n749), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n753), .B1(new_n855), .B2(new_n724), .ZN(new_n856));
  AOI211_X1 g670(.A(KEYINPUT107), .B(KEYINPUT42), .C1(new_n748), .C2(new_n749), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n854), .B(new_n818), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n850), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n850), .A3(new_n859), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n848), .B(new_n849), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n845), .B2(new_n837), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n858), .A2(new_n859), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n864), .B1(new_n863), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n693), .A2(new_n786), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n670), .A2(new_n576), .A3(new_n412), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n598), .B2(new_n599), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n411), .A3(G953), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n698), .A2(new_n719), .ZN(new_n874));
  INV_X1    g688(.A(new_n646), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n774), .A2(new_n875), .A3(new_n716), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n774), .A2(new_n875), .A3(new_n870), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT48), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n877), .A2(new_n878), .A3(new_n577), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n877), .B2(new_n577), .ZN(new_n880));
  OAI221_X1 g694(.A(new_n873), .B1(new_n874), .B2(new_n876), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n263), .A2(new_n594), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT122), .B1(new_n871), .B2(new_n882), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n871), .A2(KEYINPUT122), .A3(new_n882), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n877), .A2(new_n720), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n675), .A2(new_n679), .A3(new_n698), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT50), .B1(new_n876), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(KEYINPUT50), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n692), .A2(new_n266), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n783), .A2(new_n784), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n892), .B2(new_n726), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n885), .B(new_n889), .C1(new_n876), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n881), .B1(new_n895), .B2(KEYINPUT51), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(KEYINPUT123), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT123), .B1(new_n894), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n868), .A2(new_n869), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n799), .B1(new_n902), .B2(new_n903), .ZN(G75));
  NAND2_X1  g718(.A1(new_n858), .A2(new_n859), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT118), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n861), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n848), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(G210), .A3(G902), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n467), .A2(new_n469), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n471), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n909), .B2(new_n910), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n189), .A2(G952), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G51));
  XOR2_X1   g731(.A(new_n366), .B(KEYINPUT124), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT57), .ZN(new_n919));
  INV_X1    g733(.A(new_n863), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n849), .B1(new_n907), .B2(new_n848), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n352), .A2(new_n364), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n906), .A2(new_n861), .B1(new_n839), .B2(new_n847), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n268), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n762), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n916), .B1(new_n924), .B2(new_n927), .ZN(G54));
  NAND2_X1  g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n926), .A2(new_n250), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n250), .B1(new_n926), .B2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n916), .ZN(G60));
  AND2_X1   g747(.A1(new_n591), .A2(new_n592), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n920), .B2(new_n921), .ZN(new_n938));
  INV_X1    g752(.A(new_n916), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n936), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n868), .B2(new_n869), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n942), .B2(new_n934), .ZN(G63));
  XNOR2_X1  g757(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n400), .A2(new_n268), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n908), .A2(new_n634), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n572), .ZN(new_n948));
  INV_X1    g762(.A(new_n946), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n925), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n950), .A3(new_n939), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G66));
  OAI21_X1  g767(.A(G953), .B1(new_n415), .B2(new_n454), .ZN(new_n954));
  INV_X1    g768(.A(new_n811), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n911), .B1(G898), .B2(new_n189), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT126), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  OAI21_X1  g773(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n244), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n658), .A2(new_n786), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n577), .C1(new_n800), .C2(new_n803), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n681), .A2(new_n721), .A3(new_n833), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  NAND4_X1  g779(.A1(new_n789), .A2(new_n780), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n966), .B2(new_n189), .ZN(new_n967));
  INV_X1    g781(.A(new_n757), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n686), .A2(new_n711), .A3(new_n678), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n968), .B(new_n820), .C1(new_n769), .C2(new_n969), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n754), .A2(new_n789), .A3(new_n780), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n189), .ZN(new_n972));
  INV_X1    g786(.A(new_n961), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(G900), .B2(G953), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n967), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n966), .B2(new_n811), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n528), .B1(new_n487), .B2(new_n515), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n916), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n517), .ZN(new_n983));
  INV_X1    g797(.A(new_n979), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n971), .B2(new_n955), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n865), .A2(new_n866), .ZN(new_n987));
  NOR4_X1   g801(.A1(new_n987), .A2(new_n517), .A3(new_n981), .A4(new_n984), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n986), .B1(new_n990), .B2(new_n991), .ZN(G57));
endmodule


