//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT66), .A3(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n198), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(new_n190), .A3(new_n192), .A4(new_n193), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  OAI211_X1 g022(.A(G128), .B(new_n205), .C1(new_n206), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n211), .A2(G137), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G134), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n204), .A2(G146), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n221), .B(new_n222), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n209), .A2(new_n217), .A3(new_n220), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n222), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  XNOR2_X1  g045(.A(G143), .B(G146), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n227), .ZN(new_n233));
  AND4_X1   g047(.A1(new_n231), .A2(new_n221), .A3(new_n222), .A4(new_n227), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n212), .A2(new_n214), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n219), .A2(G131), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n236), .A2(new_n237), .B1(new_n238), .B2(G131), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n203), .B(new_n225), .C1(new_n235), .C2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G237), .A2(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G210), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT64), .B1(new_n226), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n232), .A2(new_n231), .A3(new_n227), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n248), .A2(new_n249), .B1(new_n226), .B2(new_n229), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(G131), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n217), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n209), .A2(new_n224), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n217), .A2(new_n220), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n250), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n203), .B1(new_n255), .B2(KEYINPUT30), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  OAI22_X1  g072(.A1(new_n235), .A2(new_n239), .B1(new_n225), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n225), .A2(new_n258), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n246), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n240), .A2(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n250), .A2(new_n252), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n203), .A4(new_n225), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n269), .A3(new_n260), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n200), .A2(new_n202), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n265), .A2(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI22_X1  g086(.A1(new_n263), .A2(new_n264), .B1(new_n272), .B2(new_n245), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n263), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n256), .A2(new_n262), .ZN(new_n276));
  INV_X1    g090(.A(new_n246), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n264), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n273), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n265), .A2(new_n268), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n270), .A2(new_n271), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n245), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n263), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT31), .ZN(new_n290));
  AND4_X1   g104(.A1(new_n274), .A2(new_n276), .A3(new_n264), .A4(new_n277), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n274), .B1(new_n263), .B2(new_n264), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n288), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT68), .A3(new_n281), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n283), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n284), .A2(KEYINPUT69), .A3(new_n245), .A4(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  INV_X1    g112(.A(new_n240), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n256), .B2(new_n262), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n298), .C1(new_n245), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT69), .B1(new_n272), .B2(new_n245), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT70), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n276), .A2(new_n240), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n304), .B2(new_n287), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n286), .B2(new_n287), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n305), .A2(new_n307), .A3(new_n308), .A4(new_n297), .ZN(new_n309));
  INV_X1    g123(.A(new_n255), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n271), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n284), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n287), .A2(new_n298), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n303), .A2(new_n309), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G472), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n280), .A2(new_n295), .A3(new_n282), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n296), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(G234), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n326), .A3(G125), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(G146), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n335), .A3(G146), .A4(new_n332), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n327), .A2(new_n329), .A3(new_n207), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT73), .A4(new_n207), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n334), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n191), .B2(G128), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n191), .A2(G128), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G110), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n346), .A2(KEYINPUT71), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(G110), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n223), .A2(G119), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT24), .B(G110), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n330), .A2(new_n332), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n207), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n333), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n354), .A2(new_n355), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G110), .B2(new_n351), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n342), .A2(new_n357), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G137), .ZN(new_n364));
  INV_X1    g178(.A(G953), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n365), .A2(G221), .A3(G234), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n366), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT74), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT74), .B1(new_n367), .B2(new_n368), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n325), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n367), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n362), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n349), .A2(new_n352), .A3(new_n356), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n334), .A2(new_n336), .A3(new_n341), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n369), .A2(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(KEYINPUT75), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n372), .A2(new_n322), .A3(new_n374), .A4(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n357), .A2(new_n334), .A3(new_n336), .A4(new_n341), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n371), .B1(new_n384), .B2(new_n375), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n385), .A2(KEYINPUT75), .B1(new_n363), .B2(new_n373), .ZN(new_n386));
  INV_X1    g200(.A(new_n382), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n322), .A3(new_n372), .A4(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n324), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n323), .A2(G902), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT77), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n386), .A2(new_n391), .A3(new_n372), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT9), .B(G234), .ZN(new_n394));
  OAI21_X1  g208(.A(G221), .B1(new_n394), .B2(G902), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(G107), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G101), .ZN(new_n404));
  INV_X1    g218(.A(G101), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n398), .A2(new_n401), .A3(new_n405), .A4(new_n402), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(KEYINPUT4), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(new_n408), .A3(G101), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n250), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n397), .B2(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n400), .A2(KEYINPUT78), .A3(G104), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n402), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G101), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n224), .A3(new_n209), .A4(new_n406), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT10), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n415), .A2(new_n406), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n420), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n253), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n416), .B2(new_n417), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n252), .B(KEYINPUT80), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n419), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n365), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT83), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  INV_X1    g248(.A(new_n416), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n415), .A2(new_n406), .B1(new_n209), .B2(new_n224), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n252), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(KEYINPUT82), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n415), .A2(new_n406), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n209), .A2(new_n224), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n239), .B1(new_n443), .B2(new_n416), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n444), .B2(KEYINPUT12), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT12), .B(new_n252), .C1(new_n435), .C2(new_n436), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n449), .A3(KEYINPUT12), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n432), .A2(new_n434), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n419), .A2(new_n424), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n252), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n430), .B1(new_n455), .B2(new_n426), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G469), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n322), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n322), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n239), .B1(new_n419), .B2(new_n424), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n431), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n452), .A2(new_n426), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n429), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n465), .B2(G469), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n396), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n223), .A2(G143), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n211), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n204), .A2(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n223), .A2(G143), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n473), .B2(new_n468), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n472), .A3(new_n211), .ZN(new_n475));
  INV_X1    g289(.A(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G116), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n189), .A2(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n400), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n478), .A3(G107), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n474), .A2(new_n475), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n394), .A2(new_n321), .A3(G953), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n471), .A2(new_n472), .A3(new_n211), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n211), .B1(new_n471), .B2(new_n472), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n204), .A2(G128), .ZN(new_n488));
  OAI21_X1  g302(.A(G134), .B1(new_n469), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT94), .A3(new_n475), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n477), .A2(KEYINPUT14), .A3(G107), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n481), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT14), .A4(G107), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n491), .A2(KEYINPUT95), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n493), .A2(new_n494), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n487), .A2(new_n490), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n482), .B(new_n483), .C1(new_n496), .C2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT95), .B1(new_n491), .B2(new_n495), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n497), .A3(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n483), .B1(new_n506), .B2(new_n482), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n482), .B1(new_n496), .B2(new_n500), .ZN(new_n509));
  INV_X1    g323(.A(new_n483), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(KEYINPUT96), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n513), .A2(KEYINPUT97), .A3(new_n322), .A4(new_n516), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT91), .B(G475), .Z(new_n518));
  INV_X1    g332(.A(G237), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n365), .A3(G214), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n204), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n522));
  INV_X1    g336(.A(G214), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n523), .A2(G237), .A3(G953), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n524), .B2(G143), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(KEYINPUT88), .A3(new_n204), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n215), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(G143), .ZN(new_n531));
  AOI211_X1 g345(.A(G143), .B(new_n522), .C1(new_n241), .C2(G214), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT88), .B1(new_n520), .B2(new_n204), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n529), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n327), .A2(new_n329), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G146), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n530), .A2(new_n536), .B1(new_n341), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G131), .B1(new_n524), .B2(G143), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n532), .B2(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n534), .A2(G131), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n545), .B(new_n540), .C1(new_n532), .C2(new_n533), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n525), .A2(new_n526), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n215), .B1(new_n548), .B2(new_n531), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n360), .B1(new_n549), .B2(KEYINPUT17), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n539), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n397), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n547), .A2(new_n550), .ZN(new_n557));
  INV_X1    g371(.A(new_n539), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n554), .B2(new_n553), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n518), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n553), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n546), .B1(new_n527), .B2(new_n215), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n545), .B1(new_n548), .B2(new_n540), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n334), .A2(new_n336), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT90), .A4(new_n546), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n537), .B(KEYINPUT19), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n207), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n539), .A2(new_n553), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(G475), .A2(G902), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n562), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT20), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n553), .A2(new_n559), .B1(new_n572), .B2(new_n573), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n575), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n561), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n509), .A2(new_n510), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n502), .A3(new_n501), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(KEYINPUT97), .A3(new_n322), .A4(new_n511), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n515), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n517), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G210), .B1(G237), .B2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n407), .A2(new_n271), .A3(new_n409), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT5), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n191), .A3(G116), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n195), .B1(new_n591), .B2(KEYINPUT85), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT85), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(new_n590), .A3(new_n191), .A4(G116), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n592), .B(new_n594), .C1(new_n194), .C2(new_n590), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(new_n202), .A3(new_n406), .A4(new_n415), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(G110), .B(G122), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n589), .A2(new_n596), .A3(new_n598), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(KEYINPUT6), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n442), .A2(new_n328), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n250), .B2(new_n328), .ZN(new_n604));
  INV_X1    g418(.A(G224), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(G953), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT86), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n604), .B(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT6), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n597), .A2(new_n609), .A3(new_n599), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n602), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT87), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT7), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n603), .B(new_n613), .C1(new_n250), .C2(new_n328), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT7), .B1(new_n605), .B2(G953), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n598), .B(KEYINPUT8), .ZN(new_n617));
  INV_X1    g431(.A(new_n596), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n595), .A2(new_n202), .B1(new_n406), .B2(new_n415), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n601), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n322), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n588), .B1(new_n611), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n620), .A2(new_n601), .ZN(new_n624));
  INV_X1    g438(.A(new_n615), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n614), .B(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n602), .A2(new_n608), .A3(new_n610), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n587), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G214), .B1(G237), .B2(G902), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT84), .ZN(new_n632));
  NAND2_X1  g446(.A1(G234), .A2(G237), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(G952), .A3(new_n365), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(G902), .A3(G953), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT21), .B(G898), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n630), .A2(new_n632), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n586), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n320), .A2(new_n393), .A3(new_n467), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT98), .B(G101), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G3));
  XNOR2_X1  g459(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n583), .A2(new_n511), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n582), .A2(KEYINPUT33), .A3(new_n501), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n514), .A2(G902), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n583), .A2(new_n322), .A3(new_n511), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n514), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n577), .A2(new_n580), .ZN(new_n654));
  INV_X1    g468(.A(new_n561), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n631), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n623), .B2(new_n629), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n640), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n280), .B2(G902), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n283), .A2(new_n393), .A3(new_n662), .A4(new_n294), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(new_n663), .A3(new_n467), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NAND3_X1  g480(.A1(new_n659), .A2(new_n655), .A3(new_n640), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n584), .B(new_n516), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n579), .B1(new_n578), .B2(new_n575), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT100), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n654), .B2(KEYINPUT100), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n467), .A3(new_n663), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NAND3_X1  g489(.A1(new_n283), .A2(new_n662), .A3(new_n294), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n383), .A2(new_n388), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n323), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n379), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n378), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(new_n391), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n677), .A2(new_n642), .A3(new_n467), .A4(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT101), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  AOI211_X1 g502(.A(G469), .B(G902), .C1(new_n453), .C2(new_n457), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n455), .A2(new_n426), .A3(new_n430), .ZN(new_n690));
  INV_X1    g504(.A(new_n426), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n446), .B2(new_n451), .ZN(new_n692));
  OAI211_X1 g506(.A(G469), .B(new_n690), .C1(new_n692), .C2(new_n430), .ZN(new_n693));
  INV_X1    g507(.A(new_n461), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n395), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n684), .A2(new_n659), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n634), .B(KEYINPUT102), .Z(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(new_n637), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n561), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n668), .A2(new_n671), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n320), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XOR2_X1   g521(.A(new_n702), .B(KEYINPUT39), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n467), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n245), .B1(new_n311), .B2(new_n240), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n289), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n715), .B2(G902), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n296), .A2(new_n319), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT38), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n630), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n682), .B1(new_n678), .B2(new_n323), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n631), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n719), .A2(new_n581), .A3(new_n721), .A4(new_n668), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n710), .A2(new_n711), .A3(new_n717), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  INV_X1    g539(.A(new_n702), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n653), .A2(new_n725), .A3(new_n656), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n653), .A2(new_n656), .A3(new_n726), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n698), .A2(new_n320), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  AOI22_X1  g545(.A1(new_n431), .A2(KEYINPUT83), .B1(new_n446), .B2(new_n451), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n456), .B1(new_n732), .B2(new_n434), .ZN(new_n733));
  OAI21_X1  g547(.A(G469), .B1(new_n733), .B2(G902), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n393), .A2(new_n734), .A3(new_n460), .A4(new_n395), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n320), .A2(new_n661), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n672), .A2(new_n320), .A3(new_n735), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND3_X1  g554(.A1(new_n734), .A2(new_n460), .A3(new_n395), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n697), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n586), .A2(new_n639), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n320), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  INV_X1    g559(.A(new_n585), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n584), .A2(new_n515), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n656), .B(new_n659), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n639), .ZN(new_n749));
  INV_X1    g563(.A(new_n741), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n293), .A2(new_n322), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n312), .A2(new_n287), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n290), .B(new_n753), .C1(new_n291), .C2(new_n292), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n752), .A2(G472), .B1(new_n281), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n751), .B1(new_n755), .B2(new_n393), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n281), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n751), .A2(new_n393), .A3(new_n662), .A4(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n749), .B(new_n750), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NAND4_X1  g574(.A1(new_n742), .A2(new_n727), .A3(new_n729), .A4(new_n755), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  INV_X1    g577(.A(new_n393), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT32), .B1(new_n293), .B2(new_n281), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n318), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n763), .B(new_n764), .C1(new_n766), .C2(new_n317), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n623), .A2(new_n629), .A3(new_n395), .A4(new_n631), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT106), .B1(new_n431), .B2(new_n462), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n455), .A2(new_n770), .A3(new_n426), .A4(new_n430), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n429), .A2(new_n464), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n461), .B1(new_n772), .B2(G469), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n768), .B1(new_n773), .B2(new_n460), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n767), .A2(new_n727), .A3(new_n729), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n729), .A2(new_n727), .A3(new_n774), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n320), .A2(new_n393), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n763), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  NAND4_X1  g594(.A1(new_n320), .A2(new_n705), .A3(new_n393), .A4(new_n774), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  NOR2_X1   g596(.A1(new_n465), .A2(KEYINPUT45), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n459), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n772), .A2(KEYINPUT45), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n461), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n460), .B1(new_n786), .B2(KEYINPUT46), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n395), .B(new_n708), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n653), .A2(new_n581), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n676), .A3(new_n684), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n623), .A2(new_n629), .A3(new_n631), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n795), .B2(new_n796), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n791), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  NAND2_X1  g615(.A1(new_n729), .A2(new_n727), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n802), .A2(new_n320), .A3(new_n393), .A4(new_n798), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n395), .B1(new_n788), .B2(new_n789), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT47), .B(new_n395), .C1(new_n788), .C2(new_n789), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n326), .ZN(G42));
  NAND2_X1  g624(.A1(new_n734), .A2(new_n460), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT49), .Z(new_n812));
  INV_X1    g626(.A(new_n719), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n393), .A2(new_n395), .A3(new_n632), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n792), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n717), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n798), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n635), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n735), .ZN(new_n820));
  OR4_X1    g634(.A1(new_n656), .A2(new_n819), .A3(new_n653), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n794), .A2(new_n700), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT111), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n741), .A2(new_n798), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n684), .A2(new_n662), .A3(new_n757), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n821), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n756), .A2(new_n758), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n823), .B2(new_n824), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n813), .A2(new_n631), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n750), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT113), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(KEYINPUT113), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n750), .A3(new_n837), .A4(new_n833), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n830), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n832), .A2(new_n818), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n734), .A2(new_n460), .A3(new_n396), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n807), .A2(new_n808), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n365), .B2(G952), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n819), .A2(new_n657), .A3(new_n820), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n846), .B(new_n847), .C1(KEYINPUT114), .C2(new_n365), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n766), .A2(new_n317), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n393), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n827), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n832), .A2(new_n659), .A3(new_n750), .ZN(new_n854));
  INV_X1    g668(.A(new_n850), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT115), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n825), .A2(new_n855), .A3(new_n826), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n768), .B(new_n720), .C1(new_n460), .C2(new_n466), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n517), .A2(new_n703), .A3(new_n585), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT107), .B1(new_n864), .B2(new_n671), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n576), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n579), .A2(new_n562), .A3(new_n574), .A4(new_n575), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n669), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT100), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT107), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n668), .A2(new_n870), .A3(new_n871), .A4(new_n703), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n863), .A2(new_n320), .A3(new_n865), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n729), .A2(new_n774), .A3(new_n828), .A4(new_n727), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n781), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT108), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT108), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n873), .A2(new_n781), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n656), .A2(new_n652), .A3(new_n650), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n586), .ZN(new_n881));
  INV_X1    g695(.A(new_n641), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n467), .A3(new_n882), .A4(new_n663), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n759), .A2(new_n685), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n643), .A2(new_n739), .A3(new_n744), .A4(new_n736), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n879), .A2(new_n779), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n748), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n773), .A2(new_n460), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n684), .A2(new_n396), .A3(new_n702), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n717), .A2(new_n888), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n730), .A2(new_n761), .A3(new_n706), .A4(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT52), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n862), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n892), .B(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n759), .A2(new_n685), .A3(new_n883), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n643), .A2(new_n739), .A3(new_n744), .A4(new_n736), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n779), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n761), .A2(new_n706), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n862), .B1(new_n902), .B2(KEYINPUT52), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n897), .A2(new_n900), .A3(new_n879), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n894), .A2(new_n895), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT109), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n862), .B1(new_n901), .B2(new_n896), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n897), .A2(new_n900), .A3(new_n879), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n894), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT109), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n894), .A2(new_n904), .A3(new_n911), .A4(new_n895), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n914));
  INV_X1    g728(.A(new_n808), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n784), .A2(new_n785), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n694), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT46), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n460), .A3(new_n787), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT47), .B1(new_n920), .B2(new_n395), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT112), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n842), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n915), .A2(new_n921), .A3(KEYINPUT112), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n841), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n914), .B1(new_n839), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n861), .A2(new_n913), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n817), .B1(new_n927), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n365), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n322), .B1(new_n894), .B2(new_n904), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n932), .B2(G210), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n602), .A2(new_n610), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n608), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n931), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n936), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT116), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT116), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G51));
  AOI21_X1  g755(.A(new_n895), .B1(new_n894), .B2(new_n904), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n905), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n461), .B(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n458), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n932), .A2(new_n785), .A3(new_n784), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n930), .B1(new_n947), .B2(new_n948), .ZN(G54));
  AND2_X1   g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n932), .A2(new_n578), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n578), .B1(new_n932), .B2(new_n950), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n930), .ZN(G60));
  INV_X1    g767(.A(KEYINPUT118), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n647), .A2(new_n648), .ZN(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n514), .A2(new_n322), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n930), .B1(new_n944), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n895), .B1(new_n894), .B2(new_n908), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n894), .A2(new_n895), .A3(new_n904), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n911), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n958), .B1(new_n964), .B2(new_n906), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n954), .B(new_n961), .C1(new_n965), .C2(new_n955), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n955), .B1(new_n913), .B2(new_n959), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n963), .B2(new_n942), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n931), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT118), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n966), .A2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT119), .Z(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n894), .B2(new_n904), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n386), .A2(new_n372), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n930), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT120), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n976), .A2(new_n980), .A3(new_n681), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n976), .B2(new_n681), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT121), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n981), .B2(new_n982), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI221_X1 g801(.A(new_n979), .B1(new_n984), .B2(KEYINPUT61), .C1(new_n981), .C2(new_n982), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(G66));
  OAI21_X1  g803(.A(G953), .B1(new_n638), .B2(new_n605), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n886), .B2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n934), .B1(G898), .B2(new_n365), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  NAND3_X1  g807(.A1(new_n723), .A2(new_n901), .A3(new_n730), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT62), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n803), .B1(new_n915), .B2(new_n921), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n881), .A2(new_n818), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n998), .A2(new_n777), .A3(new_n709), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n997), .A2(new_n800), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT122), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n996), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n997), .A2(new_n800), .A3(new_n999), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT122), .B1(new_n995), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n365), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n262), .B1(new_n257), .B2(new_n310), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(new_n570), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n365), .B1(G227), .B2(G900), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n850), .A2(new_n748), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n791), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n901), .A2(new_n730), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n1014), .A3(new_n779), .A4(new_n781), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n791), .A2(new_n797), .A3(new_n799), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1017), .A2(new_n809), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1016), .A2(new_n1018), .A3(KEYINPUT123), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT123), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n997), .A2(new_n800), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(new_n1015), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1019), .A2(new_n365), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1008), .B1(G900), .B2(G953), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1011), .A2(new_n1010), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1011), .A2(new_n1010), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1008), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1029), .B1(new_n1005), .B2(new_n365), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1027), .B(new_n1028), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1026), .A2(new_n1032), .ZN(G72));
  NAND3_X1  g847(.A1(new_n1002), .A2(new_n886), .A3(new_n1004), .ZN(new_n1034));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  NAND2_X1  g850(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n245), .A3(new_n304), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1036), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n304), .A2(new_n287), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1039), .B1(new_n1040), .B2(new_n289), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n930), .B1(new_n909), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT125), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1019), .A2(new_n886), .A3(new_n1022), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1043), .B1(new_n1044), .B2(new_n1036), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1044), .A2(new_n1043), .A3(new_n1036), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n300), .A2(new_n287), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT126), .Z(new_n1048));
  NAND2_X1  g862(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1038), .B(new_n1042), .C1(new_n1045), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(G57));
endmodule


