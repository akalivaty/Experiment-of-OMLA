//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT72), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT27), .B(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  OR3_X1    g014(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  AND3_X1   g016(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(G183gat), .B(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(new_n223), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR3_X1   g029(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n231));
  OAI22_X1  g030(.A1(new_n230), .A2(new_n231), .B1(new_n218), .B2(new_n219), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT64), .B(new_n224), .C1(new_n225), .C2(new_n223), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n232), .B1(new_n233), .B2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n222), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n207), .B1(new_n242), .B2(KEYINPUT29), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244));
  INV_X1    g043(.A(G211gat), .ZN(new_n245));
  INV_X1    g044(.A(G218gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G197gat), .ZN(new_n248));
  INV_X1    g047(.A(G204gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(G197gat), .A2(G204gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n253));
  XOR2_X1   g052(.A(G211gat), .B(G218gat), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n253), .B(new_n255), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n236), .A2(new_n237), .B1(new_n240), .B2(new_n239), .ZN(new_n257));
  OAI211_X1 g056(.A(G226gat), .B(G233gat), .C1(new_n257), .C2(new_n222), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n207), .B1(new_n242), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n256), .B1(new_n263), .B2(new_n258), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n206), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n263), .A2(new_n258), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n259), .B(new_n205), .C1(new_n266), .C2(new_n256), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT30), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n260), .A2(new_n264), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n205), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT0), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  INV_X1    g078(.A(G155gat), .ZN(new_n280));
  INV_X1    g079(.A(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n279), .B1(new_n282), .B2(KEYINPUT2), .ZN(new_n283));
  INV_X1    g082(.A(G141gat), .ZN(new_n284));
  INV_X1    g083(.A(G148gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n290));
  OR2_X1    g089(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n292));
  AND4_X1   g091(.A1(new_n286), .A2(new_n291), .A3(new_n287), .A4(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT73), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G155gat), .B2(G162gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(new_n279), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n290), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n279), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n291), .A2(new_n286), .A3(new_n287), .A4(new_n292), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT75), .A4(new_n294), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n289), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G120gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G113gat), .A2(G120gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT4), .B1(new_n302), .B2(new_n310), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT77), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n317), .B(new_n318), .C1(new_n311), .C2(new_n312), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n301), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n288), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n310), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n312), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n302), .A2(KEYINPUT4), .A3(new_n310), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n327), .A2(new_n329), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n311), .ZN(new_n336));
  INV_X1    g135(.A(new_n329), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n328), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n320), .A2(new_n331), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n278), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(new_n338), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n330), .B1(new_n315), .B2(new_n319), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT80), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n327), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n315), .B2(new_n319), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT39), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n337), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n329), .A3(new_n311), .ZN(new_n352));
  OAI211_X1 g151(.A(KEYINPUT39), .B(new_n352), .C1(new_n348), .C2(new_n329), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT40), .A4(new_n277), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n277), .A3(new_n353), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT40), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n273), .A2(new_n346), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n256), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n302), .B1(new_n360), .B2(new_n324), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n256), .B1(new_n325), .B2(new_n261), .ZN(new_n362));
  OAI211_X1 g161(.A(G228gat), .B(G233gat), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n366));
  OAI221_X1 g165(.A(new_n247), .B1(new_n251), .B2(new_n250), .C1(new_n254), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n255), .A2(KEYINPUT78), .A3(new_n252), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n367), .A2(new_n368), .B1(new_n366), .B2(new_n254), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n324), .B1(new_n369), .B2(new_n262), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n370), .A2(new_n322), .B1(G228gat), .B2(G233gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(new_n364), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n363), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT31), .B(G50gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G22gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n375), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n363), .B(new_n379), .C1(new_n372), .C2(new_n373), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n376), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n206), .B1(new_n269), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n386), .A2(KEYINPUT83), .B1(new_n385), .B2(new_n269), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n206), .C1(new_n269), .C2(new_n385), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n384), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT6), .B1(new_n339), .B2(new_n277), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n341), .B2(new_n345), .ZN(new_n392));
  INV_X1    g191(.A(new_n339), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n278), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n206), .A2(new_n384), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n269), .B2(new_n385), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n256), .B1(new_n243), .B2(new_n258), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n263), .A2(new_n256), .A3(new_n258), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n397), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT37), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n392), .A2(new_n394), .A3(new_n403), .A4(new_n267), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n358), .B(new_n383), .C1(new_n390), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT36), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n238), .A2(new_n241), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT69), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n221), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT69), .B1(new_n257), .B2(new_n222), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n310), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n242), .A2(new_n408), .A3(new_n326), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G15gat), .B(G43gat), .Z(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n411), .B2(new_n415), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT34), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI211_X1 g224(.A(KEYINPUT34), .B(new_n414), .C1(new_n411), .C2(new_n415), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n416), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT32), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n421), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n416), .B2(new_n417), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n423), .A2(new_n424), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n426), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n428), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n428), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n406), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n428), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n428), .A2(new_n431), .A3(new_n435), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(KEYINPUT36), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n383), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n278), .B1(new_n343), .B2(new_n344), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n320), .A2(new_n331), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n277), .A3(new_n342), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n394), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n445), .B1(new_n452), .B2(new_n273), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n405), .A2(new_n444), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n436), .A2(new_n437), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n392), .A2(new_n394), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n457));
  NOR2_X1   g256(.A1(new_n273), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(new_n456), .A3(new_n383), .A4(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n450), .A2(new_n394), .B1(new_n268), .B2(new_n271), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n441), .A2(new_n460), .A3(new_n383), .A4(new_n442), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n454), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G57gat), .B(G64gat), .Z(new_n465));
  NAND2_X1  g264(.A1(G71gat), .A2(G78gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT94), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n466), .B(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(G71gat), .A2(G78gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G71gat), .B(G78gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n465), .A2(new_n469), .A3(new_n479), .A4(new_n471), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT21), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G231gat), .A2(G233gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(G127gat), .ZN(new_n486));
  INV_X1    g285(.A(G8gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(G1gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT16), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n488), .A2(G1gat), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT90), .B(new_n487), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n493), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(KEYINPUT90), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n487), .A2(KEYINPUT90), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(new_n491), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n481), .B2(new_n482), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n486), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(new_n280), .ZN(new_n503));
  XOR2_X1   g302(.A(G183gat), .B(G211gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n501), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(KEYINPUT12), .Z(new_n512));
  INV_X1    g311(.A(G50gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(G43gat), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(G50gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT86), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(G50gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(G43gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(KEYINPUT15), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT88), .B(G43gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n524), .B2(G50gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT87), .B(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n529), .B(new_n532), .C1(new_n534), .C2(new_n531), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n522), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G43gat), .ZN(new_n539));
  AOI21_X1  g338(.A(G50gat), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n523), .B(new_n526), .C1(new_n540), .C2(new_n514), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n522), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n529), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(G36gat), .B2(new_n533), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n499), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n494), .A2(new_n498), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n538), .A2(G43gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n513), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT15), .B1(new_n551), .B2(new_n518), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n552), .B2(new_n523), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n553), .A2(new_n522), .B1(new_n542), .B2(new_n544), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n536), .B2(new_n545), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n547), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT91), .Z(new_n561));
  AOI21_X1  g360(.A(KEYINPUT18), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(new_n548), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n499), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n561), .B(KEYINPUT13), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n561), .A2(KEYINPUT18), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n536), .A2(new_n545), .A3(new_n555), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n499), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n563), .B(new_n569), .C1(new_n571), .C2(new_n557), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n512), .B1(new_n562), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n566), .B1(new_n563), .B2(new_n564), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n559), .B2(new_n569), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n561), .B(new_n563), .C1(new_n571), .C2(new_n557), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n512), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(G92gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT95), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(G99gat), .A3(G106gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n598), .A3(KEYINPUT8), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n604));
  OR2_X1    g403(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(G92gat), .A3(new_n591), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT8), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n595), .B2(KEYINPUT95), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n606), .A2(new_n590), .B1(new_n608), .B2(new_n598), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n604), .B1(new_n609), .B2(new_n600), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n599), .ZN(new_n611));
  INV_X1    g410(.A(new_n600), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT97), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n603), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n558), .A2(new_n616), .A3(new_n570), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n615), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT98), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n617), .B2(new_n618), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n588), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n587), .A3(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n481), .B1(new_n603), .B2(new_n614), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n601), .B(KEYINPUT96), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n478), .A2(new_n480), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n612), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n635), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n629), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n603), .A2(new_n481), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n636), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n636), .B2(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR4_X1   g450(.A1(new_n506), .A2(new_n583), .A3(new_n628), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n464), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n451), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n489), .ZN(G1324gat));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n272), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(KEYINPUT42), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n656), .B2(new_n487), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n660), .B2(new_n663), .ZN(G1325gat));
  INV_X1    g463(.A(new_n455), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n653), .A2(G15gat), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n653), .B2(new_n444), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n383), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT101), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n454), .A2(KEYINPUT102), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n405), .A2(new_n444), .A3(new_n674), .A4(new_n453), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n459), .A2(new_n462), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n459), .B2(new_n462), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n628), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n506), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(new_n583), .A3(new_n651), .ZN(new_n685));
  INV_X1    g484(.A(new_n628), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n454), .B2(new_n463), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n533), .B1(new_n689), .B2(new_n451), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n685), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n452), .A3(new_n534), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(G1328gat));
  OAI21_X1  g494(.A(G36gat), .B1(new_n689), .B2(new_n272), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697));
  AOI21_X1  g496(.A(G36gat), .B1(new_n697), .B2(KEYINPUT46), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n692), .A2(new_n273), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(KEYINPUT46), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(new_n701), .ZN(G1329gat));
  OAI21_X1  g501(.A(new_n524), .B1(new_n691), .B2(new_n665), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n444), .A2(new_n524), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n689), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g505(.A(new_n513), .B1(new_n691), .B2(new_n383), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n445), .A2(G50gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n689), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT48), .ZN(G1331gat));
  OAI211_X1 g509(.A(new_n673), .B(new_n675), .C1(new_n678), .C2(new_n679), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n506), .A2(new_n628), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n583), .A2(new_n711), .A3(new_n712), .A4(new_n651), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n452), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n273), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT49), .B(G64gat), .Z(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(G1333gat));
  INV_X1    g518(.A(new_n444), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n665), .A2(G71gat), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n721), .A2(G71gat), .B1(new_n713), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n713), .A2(new_n445), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n684), .A2(new_n582), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n628), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n628), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(G85gat), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n452), .A4(new_n651), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n727), .A2(new_n651), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n683), .A2(new_n688), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n451), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(G1336gat));
  OAI21_X1  g538(.A(G92gat), .B1(new_n737), .B2(new_n272), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n273), .A2(new_n589), .A3(new_n651), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT105), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n737), .B2(new_n444), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n665), .A2(G99gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n651), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1338gat));
  INV_X1    g548(.A(new_n651), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n383), .A2(G106gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n750), .B(new_n752), .C1(new_n730), .C2(new_n731), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT107), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n732), .A2(new_n651), .A3(new_n751), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n683), .A2(new_n445), .A3(new_n688), .A4(new_n736), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT53), .B1(new_n758), .B2(G106gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n758), .A2(KEYINPUT106), .A3(G106gat), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT106), .B1(new_n758), .B2(G106gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n753), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(G1339gat));
  AOI21_X1  g564(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n639), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT54), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT55), .B1(new_n768), .B2(new_n643), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n639), .A2(new_n642), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n635), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n647), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT108), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n643), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n771), .B1(new_n639), .B2(new_n766), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n646), .B1(new_n643), .B2(new_n771), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n648), .B1(new_n574), .B2(new_n581), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT55), .B1(new_n777), .B2(new_n778), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT109), .B(KEYINPUT55), .C1(new_n777), .C2(new_n778), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n781), .B(new_n782), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n559), .A2(new_n561), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n565), .A2(new_n567), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n511), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n581), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n651), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n628), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n648), .B1(new_n625), .B2(new_n627), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n781), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n785), .A2(new_n786), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n506), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n712), .A2(new_n583), .A3(new_n750), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n451), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n800), .A2(new_n455), .A3(new_n383), .A4(new_n272), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT110), .Z(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n304), .A3(new_n582), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n445), .B1(new_n798), .B2(new_n799), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n273), .A2(new_n451), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n455), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n583), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(new_n808), .ZN(G1340gat));
  NAND2_X1  g608(.A1(new_n651), .A2(new_n305), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT111), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G120gat), .B1(new_n807), .B2(new_n750), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1341gat));
  NOR3_X1   g613(.A1(new_n801), .A2(G127gat), .A3(new_n506), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n804), .A2(new_n684), .A3(new_n806), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(G127gat), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT112), .Z(G1342gat));
  OAI21_X1  g617(.A(G134gat), .B1(new_n807), .B2(new_n686), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n801), .A2(G134gat), .A3(new_n686), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT113), .B1(new_n820), .B2(KEYINPUT56), .ZN(new_n822));
  OAI221_X1 g621(.A(new_n819), .B1(KEYINPUT56), .B2(new_n820), .C1(new_n821), .C2(new_n822), .ZN(G1343gat));
  AND2_X1   g622(.A1(new_n444), .A2(new_n805), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n445), .A2(KEYINPUT57), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n772), .B(new_n647), .C1(new_n768), .C2(new_n643), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n783), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n781), .A2(new_n829), .A3(new_n782), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n628), .B1(new_n832), .B2(new_n792), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n795), .A2(new_n796), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n833), .B2(KEYINPUT116), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n506), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n825), .B1(new_n837), .B2(new_n799), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n798), .A2(new_n799), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n445), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n824), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n583), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n720), .A2(new_n383), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n800), .A2(new_n272), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n582), .A2(new_n284), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT58), .ZN(G1344gat));
  OAI211_X1 g648(.A(new_n651), .B(new_n824), .C1(new_n838), .C2(new_n842), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n851), .A3(G148gat), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n506), .A2(new_n628), .A3(new_n582), .A4(new_n651), .ZN(new_n855));
  INV_X1    g654(.A(new_n792), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n562), .A2(new_n573), .A3(new_n512), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n580), .B1(new_n576), .B2(new_n579), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n649), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n774), .B2(new_n780), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n783), .B(KEYINPUT115), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n835), .B1(new_n862), .B2(new_n628), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n855), .B1(new_n863), .B2(new_n506), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT117), .B(new_n854), .C1(new_n864), .C2(new_n383), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n506), .B1(new_n833), .B2(new_n797), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n383), .B1(new_n867), .B2(new_n799), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n445), .A3(new_n840), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n824), .A2(new_n651), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G148gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n853), .B1(new_n875), .B2(KEYINPUT59), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n285), .B1(new_n871), .B2(new_n873), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n851), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n852), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n651), .A2(new_n285), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n846), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n882), .A3(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  INV_X1    g683(.A(new_n852), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n383), .B(new_n839), .C1(new_n798), .C2(new_n799), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n854), .B1(new_n864), .B2(new_n383), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n866), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n872), .B1(new_n888), .B2(new_n865), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n853), .B(KEYINPUT59), .C1(new_n889), .C2(new_n285), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT118), .B1(new_n877), .B2(new_n851), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(new_n881), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n883), .A2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n843), .B2(new_n506), .ZN(new_n895));
  INV_X1    g694(.A(new_n846), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n280), .A3(new_n684), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n843), .B2(new_n686), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n281), .A3(new_n628), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n452), .A2(new_n272), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n804), .A2(new_n455), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n583), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n452), .B1(new_n798), .B2(new_n799), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n665), .A2(new_n445), .A3(new_n272), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n582), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n905), .B1(new_n913), .B2(new_n904), .ZN(G1348gat));
  INV_X1    g713(.A(G176gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n915), .A3(new_n651), .ZN(new_n916));
  OAI21_X1  g715(.A(G176gat), .B1(new_n903), .B2(new_n750), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1349gat));
  NOR2_X1   g717(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n912), .A2(new_n208), .A3(new_n684), .ZN(new_n920));
  OAI21_X1  g719(.A(G183gat), .B1(new_n903), .B2(new_n506), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT122), .Z(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n924), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n919), .B(new_n926), .C1(new_n920), .C2(new_n921), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n925), .A2(new_n927), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n903), .B2(new_n686), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT61), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n910), .A2(new_n209), .A3(new_n628), .A4(new_n911), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n930), .B(new_n937), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n720), .A2(new_n383), .A3(new_n272), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n910), .A2(KEYINPUT125), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n908), .B2(new_n909), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n941), .A2(new_n248), .A3(new_n582), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n871), .A2(new_n444), .A3(new_n902), .ZN(new_n946));
  OAI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n583), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT126), .ZN(G1352gat));
  OAI21_X1  g748(.A(G204gat), .B1(new_n946), .B2(new_n750), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n651), .A2(new_n249), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT62), .B1(new_n942), .B2(new_n951), .ZN(new_n952));
  OR3_X1    g751(.A1(new_n942), .A2(KEYINPUT62), .A3(new_n951), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(G1353gat));
  NAND4_X1  g753(.A1(new_n941), .A2(new_n245), .A3(new_n684), .A4(new_n944), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n946), .A2(new_n506), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n245), .B1(new_n956), .B2(KEYINPUT127), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n946), .B2(new_n506), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n957), .A2(KEYINPUT63), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  NAND4_X1  g761(.A1(new_n941), .A2(new_n246), .A3(new_n628), .A4(new_n944), .ZN(new_n963));
  OAI21_X1  g762(.A(G218gat), .B1(new_n946), .B2(new_n686), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


