

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710;

  INV_X1 U363 ( .A(G953), .ZN(n701) );
  XNOR2_X2 U364 ( .A(n581), .B(KEYINPUT2), .ZN(n635) );
  XNOR2_X2 U365 ( .A(n694), .B(n349), .ZN(n385) );
  XNOR2_X2 U366 ( .A(n348), .B(n444), .ZN(n694) );
  OR2_X1 U367 ( .A1(n666), .A2(n561), .ZN(n546) );
  NOR2_X1 U368 ( .A1(n555), .A2(n471), .ZN(n543) );
  XNOR2_X1 U369 ( .A(n394), .B(G134), .ZN(n444) );
  INV_X1 U370 ( .A(KEYINPUT70), .ZN(n343) );
  NAND2_X2 U371 ( .A1(n484), .A2(n639), .ZN(n572) );
  NOR2_X2 U372 ( .A1(n518), .A2(n637), .ZN(n692) );
  XNOR2_X2 U373 ( .A(n492), .B(n359), .ZN(n542) );
  XOR2_X2 U374 ( .A(KEYINPUT106), .B(n503), .Z(n710) );
  NOR2_X2 U375 ( .A1(n526), .A2(n502), .ZN(n503) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(G131), .Z(n430) );
  INV_X1 U377 ( .A(KEYINPUT65), .ZN(n346) );
  XNOR2_X1 U378 ( .A(n695), .B(n425), .ZN(n432) );
  XNOR2_X1 U379 ( .A(n543), .B(KEYINPUT33), .ZN(n666) );
  XNOR2_X1 U380 ( .A(n580), .B(n579), .ZN(n606) );
  NOR2_X1 U381 ( .A1(n494), .A2(n486), .ZN(n487) );
  OR2_X1 U382 ( .A1(n498), .A2(n499), .ZN(n529) );
  NOR2_X1 U383 ( .A1(n636), .A2(n492), .ZN(n559) );
  BUF_X1 U384 ( .A(n544), .Z(n561) );
  XNOR2_X1 U385 ( .A(n385), .B(n384), .ZN(n584) );
  INV_X1 U386 ( .A(KEYINPUT67), .ZN(n482) );
  AND2_X1 U387 ( .A1(n539), .A2(n707), .ZN(n340) );
  XOR2_X1 U388 ( .A(n534), .B(KEYINPUT48), .Z(n341) );
  AND2_X1 U389 ( .A1(G214), .A2(n423), .ZN(n342) );
  INV_X1 U390 ( .A(KEYINPUT83), .ZN(n505) );
  XNOR2_X1 U391 ( .A(n506), .B(n505), .ZN(n509) );
  NOR2_X2 U392 ( .A1(n509), .A2(n508), .ZN(n510) );
  INV_X1 U393 ( .A(G137), .ZN(n344) );
  INV_X1 U394 ( .A(G110), .ZN(n362) );
  XNOR2_X1 U395 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U396 ( .A(n424), .B(n342), .ZN(n425) );
  XNOR2_X1 U397 ( .A(n365), .B(n364), .ZN(n368) );
  XNOR2_X1 U398 ( .A(n514), .B(KEYINPUT36), .ZN(n515) );
  XNOR2_X1 U399 ( .A(n420), .B(KEYINPUT0), .ZN(n544) );
  BUF_X1 U400 ( .A(n624), .Z(n628) );
  NOR2_X1 U401 ( .A1(n521), .A2(n491), .ZN(n683) );
  XNOR2_X2 U402 ( .A(n343), .B(KEYINPUT4), .ZN(n391) );
  XNOR2_X1 U403 ( .A(n391), .B(n344), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n345), .B(n430), .ZN(n348) );
  XNOR2_X2 U405 ( .A(G143), .B(G128), .ZN(n347) );
  XNOR2_X2 U406 ( .A(n347), .B(n346), .ZN(n394) );
  INV_X1 U407 ( .A(G146), .ZN(n349) );
  XNOR2_X1 U408 ( .A(G107), .B(G104), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n350), .B(G110), .ZN(n352) );
  XNOR2_X1 U410 ( .A(G101), .B(KEYINPUT77), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n401) );
  XOR2_X1 U412 ( .A(G140), .B(KEYINPUT78), .Z(n354) );
  AND2_X1 U413 ( .A1(G227), .A2(n701), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n401), .B(n355), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n385), .B(n356), .ZN(n630) );
  INV_X1 U417 ( .A(G902), .ZN(n447) );
  NAND2_X1 U418 ( .A1(n630), .A2(n447), .ZN(n358) );
  INV_X1 U419 ( .A(G469), .ZN(n357) );
  XNOR2_X2 U420 ( .A(n358), .B(n357), .ZN(n492) );
  INV_X1 U421 ( .A(KEYINPUT1), .ZN(n359) );
  INV_X1 U422 ( .A(n542), .ZN(n637) );
  XOR2_X1 U423 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n361) );
  XNOR2_X1 U424 ( .A(G119), .B(KEYINPUT94), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n365) );
  XNOR2_X1 U426 ( .A(G128), .B(G137), .ZN(n363) );
  NAND2_X1 U427 ( .A1(G234), .A2(n701), .ZN(n366) );
  XOR2_X1 U428 ( .A(KEYINPUT8), .B(n366), .Z(n437) );
  NAND2_X1 U429 ( .A1(n437), .A2(G221), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n371) );
  INV_X1 U431 ( .A(G146), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n369), .B(G125), .ZN(n393) );
  XNOR2_X1 U433 ( .A(n393), .B(KEYINPUT10), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n370), .B(G140), .ZN(n695) );
  XNOR2_X1 U435 ( .A(n371), .B(n695), .ZN(n619) );
  NAND2_X1 U436 ( .A1(n619), .A2(n447), .ZN(n375) );
  XNOR2_X1 U437 ( .A(KEYINPUT15), .B(G902), .ZN(n582) );
  NAND2_X1 U438 ( .A1(G234), .A2(n582), .ZN(n372) );
  XNOR2_X1 U439 ( .A(KEYINPUT20), .B(n372), .ZN(n450) );
  NAND2_X1 U440 ( .A1(G217), .A2(n450), .ZN(n373) );
  XNOR2_X1 U441 ( .A(KEYINPUT25), .B(n373), .ZN(n374) );
  XNOR2_X2 U442 ( .A(n375), .B(n374), .ZN(n639) );
  INV_X1 U443 ( .A(n639), .ZN(n465) );
  NOR2_X1 U444 ( .A1(n637), .A2(n465), .ZN(n387) );
  XOR2_X1 U445 ( .A(G101), .B(KEYINPUT5), .Z(n377) );
  XNOR2_X1 U446 ( .A(KEYINPUT96), .B(KEYINPUT76), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n377), .B(n376), .ZN(n379) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n423) );
  NAND2_X1 U449 ( .A1(n423), .A2(G210), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U451 ( .A(G116), .B(G113), .ZN(n381) );
  XNOR2_X1 U452 ( .A(KEYINPUT3), .B(G119), .ZN(n380) );
  XNOR2_X1 U453 ( .A(n381), .B(n380), .ZN(n400) );
  INV_X1 U454 ( .A(n400), .ZN(n382) );
  XNOR2_X1 U455 ( .A(n383), .B(n382), .ZN(n384) );
  NAND2_X1 U456 ( .A1(n584), .A2(n447), .ZN(n386) );
  XNOR2_X2 U457 ( .A(n386), .B(G472), .ZN(n480) );
  XNOR2_X1 U458 ( .A(n480), .B(KEYINPUT6), .ZN(n471) );
  NAND2_X1 U459 ( .A1(n387), .A2(n471), .ZN(n458) );
  XNOR2_X1 U460 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n389) );
  NAND2_X1 U461 ( .A1(n701), .A2(G224), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U463 ( .A(n391), .B(n390), .ZN(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT79), .B(KEYINPUT88), .ZN(n392) );
  XNOR2_X1 U465 ( .A(n393), .B(n392), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n403) );
  XNOR2_X1 U468 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n398), .B(G122), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n612) );
  XNOR2_X1 U472 ( .A(n403), .B(n612), .ZN(n591) );
  NAND2_X1 U473 ( .A1(n591), .A2(n582), .ZN(n408) );
  OR2_X1 U474 ( .A1(G237), .A2(G902), .ZN(n409) );
  NAND2_X1 U475 ( .A1(n409), .A2(G210), .ZN(n406) );
  INV_X1 U476 ( .A(KEYINPUT82), .ZN(n404) );
  XNOR2_X1 U477 ( .A(n404), .B(KEYINPUT89), .ZN(n405) );
  XNOR2_X1 U478 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X2 U479 ( .A(n408), .B(n407), .ZN(n478) );
  NAND2_X1 U480 ( .A1(n409), .A2(G214), .ZN(n411) );
  INV_X1 U481 ( .A(KEYINPUT90), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n411), .B(n410), .ZN(n650) );
  OR2_X2 U483 ( .A1(n478), .A2(n650), .ZN(n511) );
  XNOR2_X2 U484 ( .A(n511), .B(KEYINPUT19), .ZN(n490) );
  XOR2_X1 U485 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n413) );
  NAND2_X1 U486 ( .A1(G234), .A2(G237), .ZN(n412) );
  XNOR2_X1 U487 ( .A(n413), .B(n412), .ZN(n415) );
  AND2_X1 U488 ( .A1(G902), .A2(n415), .ZN(n466) );
  NOR2_X1 U489 ( .A1(G898), .A2(n701), .ZN(n613) );
  NAND2_X1 U490 ( .A1(n466), .A2(n613), .ZN(n414) );
  XOR2_X1 U491 ( .A(KEYINPUT92), .B(n414), .Z(n417) );
  NAND2_X1 U492 ( .A1(n415), .A2(G952), .ZN(n416) );
  XNOR2_X1 U493 ( .A(n416), .B(KEYINPUT91), .ZN(n663) );
  AND2_X1 U494 ( .A1(n663), .A2(n701), .ZN(n469) );
  NOR2_X1 U495 ( .A1(n417), .A2(n469), .ZN(n418) );
  XNOR2_X1 U496 ( .A(n418), .B(KEYINPUT93), .ZN(n419) );
  NAND2_X1 U497 ( .A1(n490), .A2(n419), .ZN(n420) );
  INV_X1 U498 ( .A(n544), .ZN(n455) );
  XNOR2_X1 U499 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n434) );
  XOR2_X1 U500 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n422) );
  XNOR2_X1 U501 ( .A(G122), .B(KEYINPUT100), .ZN(n421) );
  XNOR2_X1 U502 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U503 ( .A(KEYINPUT12), .B(G104), .Z(n427) );
  XNOR2_X1 U504 ( .A(G143), .B(G113), .ZN(n426) );
  XNOR2_X1 U505 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U506 ( .A(n428), .B(KEYINPUT99), .ZN(n429) );
  XOR2_X1 U507 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U508 ( .A(n432), .B(n431), .ZN(n598) );
  NOR2_X1 U509 ( .A1(G902), .A2(n598), .ZN(n433) );
  XNOR2_X1 U510 ( .A(n434), .B(n433), .ZN(n436) );
  INV_X1 U511 ( .A(G475), .ZN(n435) );
  XNOR2_X1 U512 ( .A(n436), .B(n435), .ZN(n498) );
  XOR2_X1 U513 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n439) );
  NAND2_X1 U514 ( .A1(G217), .A2(n437), .ZN(n438) );
  XNOR2_X1 U515 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U516 ( .A(KEYINPUT7), .B(G122), .Z(n441) );
  XNOR2_X1 U517 ( .A(G116), .B(G107), .ZN(n440) );
  XOR2_X1 U518 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U519 ( .A(n443), .B(n442), .ZN(n446) );
  INV_X1 U520 ( .A(n444), .ZN(n445) );
  XNOR2_X1 U521 ( .A(n446), .B(n445), .ZN(n626) );
  NAND2_X1 U522 ( .A1(n626), .A2(n447), .ZN(n449) );
  INV_X1 U523 ( .A(G478), .ZN(n448) );
  XNOR2_X1 U524 ( .A(n449), .B(n448), .ZN(n473) );
  AND2_X1 U525 ( .A1(n498), .A2(n473), .ZN(n653) );
  AND2_X1 U526 ( .A1(n450), .A2(G221), .ZN(n452) );
  XNOR2_X1 U527 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U528 ( .A(n452), .B(n451), .ZN(n640) );
  INV_X1 U529 ( .A(n640), .ZN(n453) );
  AND2_X1 U530 ( .A1(n653), .A2(n453), .ZN(n454) );
  NAND2_X1 U531 ( .A1(n455), .A2(n454), .ZN(n457) );
  XNOR2_X1 U532 ( .A(KEYINPUT68), .B(KEYINPUT22), .ZN(n456) );
  XNOR2_X1 U533 ( .A(n457), .B(n456), .ZN(n461) );
  NOR2_X1 U534 ( .A1(n458), .A2(n461), .ZN(n460) );
  XNOR2_X1 U535 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n459) );
  XNOR2_X1 U536 ( .A(n460), .B(n459), .ZN(n574) );
  XOR2_X1 U537 ( .A(G119), .B(n574), .Z(G21) );
  OR2_X2 U538 ( .A1(n461), .A2(n542), .ZN(n481) );
  INV_X1 U539 ( .A(n471), .ZN(n462) );
  NOR2_X1 U540 ( .A1(n481), .A2(n462), .ZN(n463) );
  XNOR2_X1 U541 ( .A(n463), .B(KEYINPUT86), .ZN(n464) );
  NAND2_X1 U542 ( .A1(n464), .A2(n465), .ZN(n564) );
  XNOR2_X1 U543 ( .A(n564), .B(G101), .ZN(G3) );
  NOR2_X1 U544 ( .A1(n640), .A2(n465), .ZN(n470) );
  NAND2_X1 U545 ( .A1(G953), .A2(n466), .ZN(n467) );
  NOR2_X1 U546 ( .A1(G900), .A2(n467), .ZN(n468) );
  OR2_X1 U547 ( .A1(n469), .A2(n468), .ZN(n493) );
  NAND2_X1 U548 ( .A1(n470), .A2(n493), .ZN(n486) );
  NOR2_X1 U549 ( .A1(n486), .A2(n471), .ZN(n472) );
  XNOR2_X1 U550 ( .A(n472), .B(KEYINPUT104), .ZN(n474) );
  INV_X1 U551 ( .A(n473), .ZN(n499) );
  INV_X1 U552 ( .A(n529), .ZN(n686) );
  NAND2_X1 U553 ( .A1(n474), .A2(n686), .ZN(n475) );
  XNOR2_X1 U554 ( .A(n475), .B(KEYINPUT105), .ZN(n513) );
  NOR2_X1 U555 ( .A1(n650), .A2(n542), .ZN(n476) );
  NAND2_X1 U556 ( .A1(n513), .A2(n476), .ZN(n477) );
  XNOR2_X1 U557 ( .A(KEYINPUT43), .B(n477), .ZN(n479) );
  NAND2_X1 U558 ( .A1(n479), .A2(n478), .ZN(n539) );
  XNOR2_X1 U559 ( .A(n539), .B(G140), .ZN(G42) );
  INV_X1 U560 ( .A(n480), .ZN(n494) );
  INV_X1 U561 ( .A(n494), .ZN(n643) );
  NOR2_X2 U562 ( .A1(n481), .A2(n643), .ZN(n483) );
  XNOR2_X1 U563 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U564 ( .A(G110), .B(KEYINPUT112), .ZN(n485) );
  XNOR2_X1 U565 ( .A(n572), .B(n485), .ZN(G12) );
  XNOR2_X1 U566 ( .A(n487), .B(KEYINPUT28), .ZN(n489) );
  XNOR2_X1 U567 ( .A(n492), .B(KEYINPUT107), .ZN(n488) );
  NAND2_X1 U568 ( .A1(n489), .A2(n488), .ZN(n521) );
  INV_X1 U569 ( .A(n490), .ZN(n491) );
  NAND2_X1 U570 ( .A1(n498), .A2(n499), .ZN(n675) );
  NAND2_X1 U571 ( .A1(n529), .A2(n675), .ZN(n655) );
  NAND2_X1 U572 ( .A1(n683), .A2(n655), .ZN(n507) );
  NAND2_X1 U573 ( .A1(n507), .A2(KEYINPUT47), .ZN(n504) );
  OR2_X1 U574 ( .A1(n640), .A2(n639), .ZN(n636) );
  AND2_X1 U575 ( .A1(n493), .A2(n559), .ZN(n497) );
  NOR2_X1 U576 ( .A1(n494), .A2(n650), .ZN(n495) );
  XNOR2_X1 U577 ( .A(n495), .B(KEYINPUT30), .ZN(n496) );
  NAND2_X1 U578 ( .A1(n497), .A2(n496), .ZN(n526) );
  INV_X1 U579 ( .A(n498), .ZN(n500) );
  AND2_X1 U580 ( .A1(n500), .A2(n499), .ZN(n547) );
  INV_X1 U581 ( .A(n478), .ZN(n501) );
  NAND2_X1 U582 ( .A1(n547), .A2(n501), .ZN(n502) );
  NAND2_X1 U583 ( .A1(n504), .A2(n710), .ZN(n506) );
  NOR2_X1 U584 ( .A1(KEYINPUT47), .A2(n507), .ZN(n508) );
  XNOR2_X1 U585 ( .A(n510), .B(KEYINPUT74), .ZN(n520) );
  INV_X1 U586 ( .A(n511), .ZN(n512) );
  NAND2_X1 U587 ( .A1(n513), .A2(n512), .ZN(n516) );
  XOR2_X1 U588 ( .A(KEYINPUT87), .B(KEYINPUT109), .Z(n514) );
  XNOR2_X1 U589 ( .A(n516), .B(n515), .ZN(n517) );
  INV_X1 U590 ( .A(n517), .ZN(n518) );
  XNOR2_X1 U591 ( .A(n692), .B(KEYINPUT85), .ZN(n519) );
  NAND2_X1 U592 ( .A1(n520), .A2(n519), .ZN(n533) );
  XOR2_X1 U593 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n524) );
  INV_X1 U594 ( .A(KEYINPUT38), .ZN(n522) );
  XNOR2_X1 U595 ( .A(n478), .B(n522), .ZN(n651) );
  NOR2_X1 U596 ( .A1(n651), .A2(n650), .ZN(n656) );
  NAND2_X1 U597 ( .A1(n653), .A2(n656), .ZN(n523) );
  XNOR2_X1 U598 ( .A(n524), .B(n523), .ZN(n667) );
  NOR2_X1 U599 ( .A1(n521), .A2(n667), .ZN(n525) );
  XNOR2_X1 U600 ( .A(n525), .B(KEYINPUT42), .ZN(n709) );
  NOR2_X1 U601 ( .A1(n526), .A2(n651), .ZN(n528) );
  XNOR2_X1 U602 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n527) );
  XNOR2_X1 U603 ( .A(n528), .B(n527), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U605 ( .A(KEYINPUT40), .B(n530), .ZN(n706) );
  NOR2_X1 U606 ( .A1(n709), .A2(n706), .ZN(n531) );
  XOR2_X1 U607 ( .A(KEYINPUT46), .B(n531), .Z(n532) );
  NOR2_X2 U608 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U609 ( .A(KEYINPUT84), .ZN(n534) );
  XNOR2_X1 U610 ( .A(n535), .B(n341), .ZN(n540) );
  NOR2_X1 U611 ( .A1(n536), .A2(n675), .ZN(n538) );
  INV_X1 U612 ( .A(KEYINPUT110), .ZN(n537) );
  XNOR2_X1 U613 ( .A(n538), .B(n537), .ZN(n707) );
  NAND2_X1 U614 ( .A1(n540), .A2(n340), .ZN(n699) );
  INV_X1 U615 ( .A(n636), .ZN(n541) );
  NAND2_X1 U616 ( .A1(n542), .A2(n541), .ZN(n555) );
  XNOR2_X1 U617 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n545) );
  XNOR2_X1 U618 ( .A(n546), .B(n545), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n547), .B(KEYINPUT80), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X2 U621 ( .A(n550), .B(KEYINPUT35), .ZN(n605) );
  NOR2_X1 U622 ( .A1(n574), .A2(KEYINPUT69), .ZN(n551) );
  NAND2_X1 U623 ( .A1(n551), .A2(n572), .ZN(n552) );
  NOR2_X1 U624 ( .A1(n605), .A2(n552), .ZN(n554) );
  INV_X1 U625 ( .A(KEYINPUT44), .ZN(n553) );
  NOR2_X1 U626 ( .A1(n554), .A2(n553), .ZN(n567) );
  OR2_X1 U627 ( .A1(n555), .A2(n494), .ZN(n646) );
  OR2_X1 U628 ( .A1(n646), .A2(n561), .ZN(n558) );
  XNOR2_X1 U629 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n556) );
  XOR2_X1 U630 ( .A(n556), .B(KEYINPUT97), .Z(n557) );
  XNOR2_X1 U631 ( .A(n558), .B(n557), .ZN(n690) );
  INV_X1 U632 ( .A(n559), .ZN(n560) );
  OR2_X1 U633 ( .A1(n643), .A2(n560), .ZN(n562) );
  NOR2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n676) );
  OR2_X1 U635 ( .A1(n690), .A2(n676), .ZN(n563) );
  NAND2_X1 U636 ( .A1(n563), .A2(n655), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n578) );
  INV_X1 U639 ( .A(n605), .ZN(n569) );
  NOR2_X1 U640 ( .A1(KEYINPUT69), .A2(KEYINPUT44), .ZN(n568) );
  NAND2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n605), .A2(KEYINPUT69), .ZN(n570) );
  NAND2_X1 U643 ( .A1(n571), .A2(n570), .ZN(n576) );
  INV_X1 U644 ( .A(n572), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n579) );
  NOR2_X2 U649 ( .A1(n699), .A2(n606), .ZN(n581) );
  NOR2_X2 U650 ( .A1(n635), .A2(n582), .ZN(n624) );
  NAND2_X1 U651 ( .A1(n624), .A2(G472), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n583) );
  XNOR2_X1 U653 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n586), .B(n585), .ZN(n588) );
  INV_X1 U655 ( .A(G952), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n587), .A2(G953), .ZN(n622) );
  NAND2_X1 U657 ( .A1(n588), .A2(n622), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n589), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U659 ( .A1(n624), .A2(G210), .ZN(n593) );
  XOR2_X1 U660 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n590) );
  XNOR2_X1 U661 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n593), .B(n592), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n594), .A2(n622), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n595) );
  XNOR2_X1 U665 ( .A(n596), .B(n595), .ZN(G51) );
  INV_X1 U666 ( .A(KEYINPUT60), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n624), .A2(G475), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n597) );
  XNOR2_X1 U669 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n601), .A2(n622), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n603), .B(n602), .ZN(G60) );
  XNOR2_X1 U673 ( .A(G122), .B(KEYINPUT125), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(G24) );
  BUF_X1 U675 ( .A(n606), .Z(n607) );
  NOR2_X1 U676 ( .A1(n607), .A2(G953), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G953), .A2(G224), .ZN(n608) );
  XNOR2_X1 U678 ( .A(KEYINPUT61), .B(n608), .ZN(n609) );
  AND2_X1 U679 ( .A1(n609), .A2(G898), .ZN(n610) );
  NOR2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n617) );
  INV_X1 U681 ( .A(n612), .ZN(n615) );
  INV_X1 U682 ( .A(n613), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U684 ( .A(n617), .B(n616), .ZN(G69) );
  NAND2_X1 U685 ( .A1(n628), .A2(G217), .ZN(n621) );
  XNOR2_X1 U686 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U689 ( .A(n622), .ZN(n633) );
  NOR2_X1 U690 ( .A1(n623), .A2(n633), .ZN(G66) );
  NAND2_X1 U691 ( .A1(n624), .A2(G478), .ZN(n625) );
  XOR2_X1 U692 ( .A(n626), .B(n625), .Z(n627) );
  NOR2_X1 U693 ( .A1(n627), .A2(n633), .ZN(G63) );
  NAND2_X1 U694 ( .A1(n628), .A2(G469), .ZN(n632) );
  XNOR2_X1 U695 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n629) );
  XNOR2_X1 U696 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U697 ( .A(n632), .B(n631), .ZN(n634) );
  NOR2_X1 U698 ( .A1(n634), .A2(n633), .ZN(G54) );
  NAND2_X1 U699 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U700 ( .A(n638), .B(KEYINPUT50), .ZN(n645) );
  NAND2_X1 U701 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U702 ( .A(KEYINPUT49), .B(n641), .ZN(n642) );
  NOR2_X1 U703 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U704 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U705 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U706 ( .A(KEYINPUT51), .B(n648), .ZN(n649) );
  NOR2_X1 U707 ( .A1(n667), .A2(n649), .ZN(n661) );
  NAND2_X1 U708 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U709 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U710 ( .A(n654), .B(KEYINPUT117), .ZN(n658) );
  AND2_X1 U711 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U712 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U713 ( .A1(n659), .A2(n666), .ZN(n660) );
  NOR2_X1 U714 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U715 ( .A(n662), .B(KEYINPUT52), .Z(n664) );
  NAND2_X1 U716 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U717 ( .A1(n665), .A2(n701), .ZN(n670) );
  NOR2_X1 U718 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U719 ( .A(n668), .B(KEYINPUT118), .ZN(n669) );
  NOR2_X1 U720 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U721 ( .A1(n635), .A2(n671), .ZN(n673) );
  XNOR2_X1 U722 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n672) );
  XNOR2_X1 U723 ( .A(n673), .B(n672), .ZN(G75) );
  NAND2_X1 U724 ( .A1(n676), .A2(n686), .ZN(n674) );
  XNOR2_X1 U725 ( .A(n674), .B(G104), .ZN(G6) );
  XOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n678) );
  INV_X1 U727 ( .A(n675), .ZN(n689) );
  NAND2_X1 U728 ( .A1(n676), .A2(n689), .ZN(n677) );
  XNOR2_X1 U729 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U730 ( .A(G107), .B(n679), .ZN(G9) );
  XOR2_X1 U731 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n681) );
  NAND2_X1 U732 ( .A1(n683), .A2(n689), .ZN(n680) );
  XNOR2_X1 U733 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U734 ( .A(G128), .B(n682), .Z(G30) );
  NAND2_X1 U735 ( .A1(n683), .A2(n686), .ZN(n684) );
  XNOR2_X1 U736 ( .A(n684), .B(KEYINPUT114), .ZN(n685) );
  XNOR2_X1 U737 ( .A(G146), .B(n685), .ZN(G48) );
  XOR2_X1 U738 ( .A(G113), .B(KEYINPUT115), .Z(n688) );
  NAND2_X1 U739 ( .A1(n686), .A2(n690), .ZN(n687) );
  XNOR2_X1 U740 ( .A(n688), .B(n687), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U742 ( .A(n691), .B(G116), .ZN(G18) );
  XNOR2_X1 U743 ( .A(G125), .B(n692), .ZN(n693) );
  XNOR2_X1 U744 ( .A(n693), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U745 ( .A(n694), .B(n695), .ZN(n700) );
  XNOR2_X1 U746 ( .A(G227), .B(n700), .ZN(n696) );
  NAND2_X1 U747 ( .A1(n696), .A2(G900), .ZN(n697) );
  NAND2_X1 U748 ( .A1(G953), .A2(n697), .ZN(n698) );
  XNOR2_X1 U749 ( .A(n698), .B(KEYINPUT124), .ZN(n704) );
  XNOR2_X1 U750 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U751 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U752 ( .A1(n704), .A2(n703), .ZN(G72) );
  XOR2_X1 U753 ( .A(G131), .B(KEYINPUT126), .Z(n705) );
  XNOR2_X1 U754 ( .A(n706), .B(n705), .ZN(G33) );
  XNOR2_X1 U755 ( .A(G134), .B(n707), .ZN(n708) );
  XNOR2_X1 U756 ( .A(n708), .B(KEYINPUT116), .ZN(G36) );
  XOR2_X1 U757 ( .A(G137), .B(n709), .Z(G39) );
  XNOR2_X1 U758 ( .A(G143), .B(n710), .ZN(G45) );
endmodule

