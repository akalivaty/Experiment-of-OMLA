//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G50gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n217), .A3(new_n203), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n207), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n214), .A2(new_n207), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT17), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT16), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n224), .A2(G1gat), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n227), .A2(new_n228), .A3(G8gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XOR2_X1   g029(.A(G15gat), .B(G22gat), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n225), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n226), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n207), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n211), .A2(new_n213), .B1(new_n218), .B2(new_n219), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n236), .B(new_n237), .C1(new_n238), .C2(new_n207), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT91), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n221), .A2(new_n222), .ZN(new_n244));
  OAI21_X1  g043(.A(G8gat), .B1(new_n227), .B2(new_n228), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n232), .A2(new_n230), .A3(new_n233), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n240), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(KEYINPUT92), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n244), .B(new_n247), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n242), .B(KEYINPUT13), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G197gat), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT11), .B(G169gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT12), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n251), .A2(new_n264), .A3(new_n253), .A4(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G148gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT80), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G148gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n273), .A3(G141gat), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n270), .A2(G141gat), .ZN(new_n275));
  AND2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278));
  INV_X1    g077(.A(G155gat), .ZN(new_n279));
  INV_X1    g078(.A(G162gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n274), .A2(new_n275), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT79), .B1(new_n283), .B2(new_n276), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT78), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT2), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n278), .A2(KEYINPUT78), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n277), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n270), .A2(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n279), .A2(new_n280), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n282), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(G113gat), .A2(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G113gat), .A2(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(KEYINPUT73), .A3(new_n302), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G127gat), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n309), .A2(KEYINPUT72), .A3(G134gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n298), .B2(KEYINPUT72), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n304), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n312), .A3(KEYINPUT82), .A4(new_n297), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n278), .A2(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n286), .A2(KEYINPUT2), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n276), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n291), .B1(new_n319), .B2(new_n285), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n283), .A2(KEYINPUT79), .A3(new_n276), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n295), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n282), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n311), .ZN(new_n325));
  INV_X1    g124(.A(new_n304), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT4), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n315), .A2(new_n316), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n312), .B1(new_n324), .B2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n333), .A3(new_n323), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n327), .B1(new_n296), .B2(new_n333), .ZN(new_n336));
  AOI211_X1 g135(.A(KEYINPUT3), .B(new_n282), .C1(new_n292), .C2(new_n295), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n336), .A2(KEYINPUT81), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n329), .B(new_n330), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n330), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n327), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n296), .A2(new_n312), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT81), .B1(new_n336), .B2(new_n337), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n352), .A2(KEYINPUT79), .B1(new_n275), .B2(new_n290), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n294), .B1(new_n353), .B2(new_n289), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(new_n354), .B2(new_n282), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(new_n331), .A3(new_n327), .A4(new_n334), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n351), .A2(new_n356), .B1(new_n313), .B2(new_n328), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n269), .B1(new_n346), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n339), .A2(new_n345), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n350), .B1(new_n361), .B2(KEYINPUT87), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n340), .B1(new_n351), .B2(new_n356), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n344), .B1(new_n363), .B2(new_n329), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n328), .A2(new_n313), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n365), .B(new_n358), .C1(new_n335), .C2(new_n338), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n360), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n346), .A2(new_n366), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n350), .A3(new_n269), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT67), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(G169gat), .A3(G176gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT68), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT68), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382));
  NOR2_X1   g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n379), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT69), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT69), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(G183gat), .A3(G190gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT24), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(G183gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT70), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT70), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G183gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n394), .B(new_n395), .C1(G190gat), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n389), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n395), .A2(KEYINPUT66), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n395), .A2(KEYINPUT66), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n378), .B(new_n402), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n409));
  AOI22_X1  g208(.A1(new_n388), .A2(new_n401), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT26), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n383), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n378), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n389), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G190gat), .ZN(new_n415));
  AND2_X1   g214(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT28), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT28), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n400), .B2(KEYINPUT27), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(G190gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n312), .B1(new_n410), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n426), .B(KEYINPUT64), .Z(new_n427));
  NAND4_X1  g226(.A1(new_n401), .A2(new_n381), .A3(new_n379), .A4(new_n387), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n409), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n389), .ZN(new_n431));
  INV_X1    g230(.A(new_n412), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n378), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT71), .ZN(new_n434));
  INV_X1    g233(.A(new_n417), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT70), .B(G183gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT28), .B1(new_n438), .B2(new_n415), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n433), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n430), .A2(new_n440), .A3(new_n327), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n427), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(KEYINPUT74), .A3(new_n443), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n442), .B2(KEYINPUT32), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n450), .A2(new_n443), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n442), .A2(KEYINPUT32), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT75), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n442), .A2(new_n456), .A3(KEYINPUT32), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n425), .A2(new_n441), .ZN(new_n460));
  INV_X1    g259(.A(new_n427), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n461), .B2(KEYINPUT76), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n460), .B(new_n461), .C1(KEYINPUT76), .C2(new_n463), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n410), .B2(new_n424), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(G197gat), .A2(G204gat), .ZN(new_n479));
  AND2_X1   g278(.A1(G197gat), .A2(G204gat), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n478), .B(KEYINPUT77), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G211gat), .B(G218gat), .Z(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n480), .A2(new_n479), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(new_n477), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n486), .A2(new_n481), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n483), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT29), .B1(new_n430), .B2(new_n440), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n476), .B(new_n488), .C1(new_n489), .C2(new_n475), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n420), .A2(new_n423), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n433), .B1(new_n428), .B2(new_n429), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n474), .B1(new_n493), .B2(KEYINPUT29), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n488), .B1(new_n494), .B2(new_n476), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n473), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n482), .B1(new_n486), .B2(new_n481), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n489), .A2(new_n475), .ZN(new_n500));
  INV_X1    g299(.A(new_n476), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n490), .A3(new_n472), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n503), .A3(KEYINPUT30), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n491), .A2(new_n495), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n472), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n467), .A2(new_n452), .A3(new_n458), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n469), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n497), .B2(new_n498), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n333), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n324), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n499), .B1(new_n337), .B2(KEYINPUT29), .ZN(new_n517));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n488), .B1(new_n334), .B2(new_n513), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n296), .B1(new_n514), .B2(new_n333), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G50gat), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n520), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n512), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n524), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n519), .B1(new_n516), .B2(new_n517), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n521), .A2(new_n522), .A3(new_n518), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n511), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT85), .B(G22gat), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n527), .B2(new_n533), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT88), .B(KEYINPUT35), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n373), .A2(new_n510), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT84), .ZN(new_n542));
  INV_X1    g341(.A(new_n350), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n366), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n542), .B(new_n268), .C1(new_n544), .C2(new_n364), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n350), .B1(new_n364), .B2(new_n367), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n346), .A2(new_n359), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n542), .B1(new_n548), .B2(new_n268), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n372), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n535), .A2(new_n536), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n467), .A2(new_n452), .A3(new_n458), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n467), .B1(new_n452), .B2(new_n458), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n550), .A2(new_n508), .A3(new_n551), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n373), .A2(new_n510), .A3(new_n538), .A4(KEYINPUT89), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(new_n508), .ZN(new_n559));
  INV_X1    g358(.A(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(KEYINPUT36), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n552), .B2(new_n553), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n351), .A2(new_n356), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n330), .B1(new_n565), .B2(new_n365), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n341), .A2(new_n342), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT39), .B1(new_n567), .B2(new_n340), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT39), .ZN(new_n570));
  AOI211_X1 g369(.A(KEYINPUT86), .B(new_n350), .C1(new_n566), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n365), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n570), .A3(new_n340), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n574), .B2(new_n543), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n569), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n543), .B1(new_n371), .B2(new_n368), .ZN(new_n579));
  INV_X1    g378(.A(new_n369), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n508), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(KEYINPUT40), .B(new_n569), .C1(new_n571), .C2(new_n575), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT37), .B1(new_n491), .B2(new_n495), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n502), .A2(new_n585), .A3(new_n490), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n586), .A3(new_n473), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n587), .A2(KEYINPUT38), .B1(new_n505), .B2(new_n472), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n587), .A2(KEYINPUT38), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n370), .A2(new_n588), .A3(new_n372), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n583), .A2(new_n590), .A3(new_n551), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n564), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n267), .B1(new_n558), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n550), .ZN(new_n594));
  XOR2_X1   g393(.A(G71gat), .B(G78gat), .Z(new_n595));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G57gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(G64gat), .ZN(new_n601));
  INV_X1    g400(.A(G64gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(G57gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G71gat), .B(G78gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT93), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n601), .A2(KEYINPUT94), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n605), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n235), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n610), .A2(new_n605), .A3(new_n611), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n619), .A2(new_n609), .B1(new_n599), .B2(new_n606), .ZN(new_n620));
  INV_X1    g419(.A(G231gat), .ZN(new_n621));
  INV_X1    g420(.A(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n620), .A2(KEYINPUT21), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n613), .B2(new_n614), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT96), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G183gat), .B(G211gat), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n629), .B1(new_n624), .B2(new_n626), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n633), .B1(new_n631), .B2(new_n634), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n618), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n617), .A3(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(KEYINPUT8), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT7), .ZN(new_n645));
  OAI211_X1 g444(.A(G85gat), .B(G92gat), .C1(new_n645), .C2(KEYINPUT97), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(KEYINPUT7), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(KEYINPUT97), .A3(KEYINPUT98), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n644), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(G99gat), .A2(G106gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n646), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n649), .A2(new_n650), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n651), .ZN(new_n662));
  INV_X1    g461(.A(new_n657), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n644), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n223), .A3(new_n239), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n244), .A2(new_n658), .A3(new_n664), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  NAND3_X1  g467(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  XOR2_X1   g474(.A(G190gat), .B(G218gat), .Z(new_n676));
  XNOR2_X1  g475(.A(G134gat), .B(G162gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n674), .B2(new_n675), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n641), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n613), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n620), .A2(new_n658), .A3(new_n664), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(G230gat), .A3(G233gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G120gat), .B(G148gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(G176gat), .B(G204gat), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n686), .B(new_n687), .Z(new_n688));
  AND2_X1   g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(G230gat), .A2(G233gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n683), .A2(KEYINPUT100), .A3(KEYINPUT10), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n682), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n693), .B(KEYINPUT101), .Z(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n692), .A2(new_n682), .A3(new_n694), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n685), .ZN(new_n701));
  INV_X1    g500(.A(new_n688), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI211_X1 g502(.A(KEYINPUT102), .B(new_n688), .C1(new_n700), .C2(new_n685), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n696), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n593), .A2(new_n594), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT103), .B(G1gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1324gat));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n593), .A2(new_n706), .ZN(new_n711));
  OAI21_X1  g510(.A(G8gat), .B1(new_n711), .B2(new_n508), .ZN(new_n712));
  INV_X1    g511(.A(new_n508), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT16), .B(G8gat), .Z(new_n714));
  NAND4_X1  g513(.A1(new_n593), .A2(new_n713), .A3(new_n706), .A4(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n710), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n710), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT104), .ZN(G1325gat));
  NAND2_X1  g517(.A1(new_n561), .A2(new_n563), .ZN(new_n719));
  OAI21_X1  g518(.A(G15gat), .B1(new_n711), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n554), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(G15gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n711), .B2(new_n722), .ZN(G1326gat));
  NOR2_X1   g522(.A1(new_n711), .A2(new_n551), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT43), .B(G22gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  NOR2_X1   g525(.A1(new_n679), .A2(new_n680), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n558), .B2(new_n592), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n705), .A2(new_n267), .A3(new_n641), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n212), .A3(new_n594), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n558), .A2(new_n592), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT44), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n737), .B(new_n728), .C1(new_n558), .C2(new_n592), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n730), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(new_n594), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n741), .B2(new_n212), .ZN(G1328gat));
  NAND3_X1  g541(.A1(new_n732), .A2(new_n208), .A3(new_n713), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n740), .A2(new_n713), .ZN(new_n748));
  OAI221_X1 g547(.A(new_n747), .B1(new_n745), .B2(new_n743), .C1(new_n748), .C2(new_n208), .ZN(G1329gat));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n727), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n737), .ZN(new_n752));
  INV_X1    g551(.A(new_n719), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n729), .A2(KEYINPUT44), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n730), .A4(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(G43gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n732), .A2(new_n203), .A3(new_n554), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n750), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(KEYINPUT47), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n203), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n739), .A2(KEYINPUT106), .A3(new_n753), .A4(new_n730), .ZN(new_n763));
  AOI211_X1 g562(.A(KEYINPUT107), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n755), .A2(new_n761), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n763), .A3(G43gat), .ZN(new_n767));
  INV_X1    g566(.A(new_n760), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n759), .B1(new_n764), .B2(new_n769), .ZN(G1330gat));
  AOI21_X1  g569(.A(new_n551), .B1(new_n215), .B2(new_n217), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n740), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n215), .B(new_n217), .C1(new_n731), .C2(new_n551), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g574(.A(new_n696), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n701), .A2(new_n702), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT102), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n701), .A2(new_n697), .A3(new_n702), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n681), .A2(new_n266), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n735), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n594), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g583(.A(new_n508), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT108), .Z(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1333gat));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n753), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n721), .A2(G71gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(G71gat), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g592(.A1(new_n782), .A2(new_n560), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g594(.A1(new_n641), .A2(new_n266), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n780), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n752), .A2(new_n594), .A3(new_n754), .A4(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n739), .A2(KEYINPUT109), .A3(new_n594), .A4(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(G85gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n751), .B2(new_n797), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n805), .A2(KEYINPUT110), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n729), .A2(KEYINPUT51), .A3(new_n796), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(KEYINPUT110), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n550), .A2(G85gat), .A3(new_n780), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n803), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1336gat));
  AND3_X1   g614(.A1(new_n752), .A2(new_n754), .A3(new_n798), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n713), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G92gat), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n780), .A2(G92gat), .A3(new_n508), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n806), .A2(new_n808), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n817), .A2(G92gat), .B1(new_n823), .B2(new_n821), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n820), .A2(new_n822), .B1(new_n824), .B2(new_n819), .ZN(G1337gat));
  NAND2_X1  g624(.A1(new_n816), .A2(new_n753), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G99gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n721), .A2(G99gat), .A3(new_n780), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n806), .A2(new_n808), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1338gat));
  NOR3_X1   g633(.A1(new_n551), .A2(G106gat), .A3(new_n780), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n823), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n752), .A2(new_n560), .A3(new_n754), .A4(new_n798), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(G106gat), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT53), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(G106gat), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n806), .A2(new_n808), .A3(new_n835), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n839), .B1(new_n842), .B2(new_n845), .ZN(G1339gat));
  NAND2_X1  g645(.A1(new_n694), .A2(new_n682), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT10), .B1(new_n683), .B2(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n698), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n695), .A3(KEYINPUT54), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n847), .A2(new_n848), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n699), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT55), .A4(new_n702), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n696), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n702), .A3(new_n853), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n727), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n254), .A2(new_n255), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n243), .B1(new_n240), .B2(new_n248), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n261), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n265), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n780), .B2(new_n863), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n855), .A2(new_n266), .A3(new_n858), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  INV_X1    g666(.A(new_n863), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n705), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n727), .B1(new_n870), .B2(KEYINPUT117), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n865), .A2(new_n866), .A3(new_n872), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n864), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n706), .B2(new_n267), .ZN(new_n876));
  NOR4_X1   g675(.A1(new_n681), .A2(new_n705), .A3(KEYINPUT115), .A4(new_n266), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n874), .A2(new_n641), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n551), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n594), .A3(new_n510), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n267), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n780), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(G120gat), .Z(G1341gat));
  INV_X1    g683(.A(new_n641), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(new_n309), .ZN(G1342gat));
  OAI21_X1  g686(.A(G134gat), .B1(new_n880), .B2(new_n728), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n727), .A2(new_n508), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n721), .A2(new_n889), .A3(G134gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n879), .A2(new_n594), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n719), .A2(new_n594), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n713), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n551), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n266), .A2(new_n854), .A3(new_n696), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT55), .B1(new_n856), .B2(KEYINPUT118), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n850), .A2(new_n853), .A3(new_n902), .A4(new_n702), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n780), .A2(new_n863), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n728), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n864), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT119), .B(new_n728), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n641), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n876), .A2(new_n877), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT120), .B(new_n899), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n266), .A2(new_n696), .A3(new_n854), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n849), .A2(new_n695), .A3(KEYINPUT54), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n702), .B1(new_n700), .B2(KEYINPUT54), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT118), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n857), .A3(new_n903), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n914), .A2(new_n918), .B1(new_n705), .B2(new_n868), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n907), .B1(new_n919), .B2(new_n727), .ZN(new_n920));
  INV_X1    g719(.A(new_n864), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n909), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n911), .B1(new_n922), .B2(new_n885), .ZN(new_n923));
  INV_X1    g722(.A(new_n899), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n912), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n878), .B2(new_n560), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n266), .B(new_n897), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G141gat), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n878), .A2(new_n560), .ZN(new_n930));
  INV_X1    g729(.A(new_n896), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n267), .A2(G141gat), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n930), .A2(new_n508), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT58), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1344gat));
  NAND2_X1  g737(.A1(new_n271), .A2(new_n273), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n780), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n930), .A2(new_n508), .A3(new_n931), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n897), .A2(new_n705), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n863), .B1(new_n859), .B2(KEYINPUT121), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(KEYINPUT121), .B2(new_n859), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n906), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n946), .A2(new_n885), .B1(new_n267), .B2(new_n706), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n898), .B1(new_n947), .B2(new_n551), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n878), .A2(new_n899), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n270), .B1(new_n950), .B2(KEYINPUT122), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n705), .B(new_n897), .C1(new_n926), .C2(new_n927), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(new_n942), .A3(new_n939), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n941), .B1(new_n953), .B2(new_n955), .ZN(G1345gat));
  OAI211_X1 g755(.A(new_n641), .B(new_n897), .C1(new_n926), .C2(new_n927), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G155gat), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n885), .A2(G155gat), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n930), .A2(new_n508), .A3(new_n931), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n958), .A2(KEYINPUT123), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1346gat));
  OAI211_X1 g764(.A(new_n727), .B(new_n897), .C1(new_n926), .C2(new_n927), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G162gat), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n889), .A2(G162gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n930), .A2(new_n931), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n967), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1347gat));
  NOR2_X1   g773(.A1(new_n594), .A2(new_n508), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n976), .A2(new_n721), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n879), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(G169gat), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(new_n267), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n878), .A2(new_n550), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n560), .A2(new_n721), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n713), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n981), .A2(new_n266), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n980), .B1(new_n979), .B2(new_n987), .ZN(G1348gat));
  OAI21_X1  g787(.A(G176gat), .B1(new_n978), .B2(new_n780), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n981), .A2(new_n986), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n780), .A2(G176gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(G1349gat));
  OAI21_X1  g791(.A(new_n400), .B1(new_n978), .B2(new_n885), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n416), .A2(new_n417), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n981), .A2(new_n994), .A3(new_n641), .A4(new_n986), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(KEYINPUT60), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT60), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n993), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n997), .A2(new_n999), .ZN(G1350gat));
  NOR3_X1   g799(.A1(new_n990), .A2(G190gat), .A3(new_n728), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n879), .A2(new_n727), .A3(new_n977), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1002), .B1(new_n1003), .B2(G190gat), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT61), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1003), .A2(G190gat), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT61), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(G1351gat));
  NOR3_X1   g810(.A1(new_n753), .A2(new_n508), .A3(new_n551), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n267), .A2(G197gat), .ZN(new_n1013));
  AND4_X1   g812(.A1(new_n550), .A2(new_n878), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n948), .A2(new_n949), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n976), .A2(new_n753), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1015), .A2(new_n266), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1014), .B1(new_n1017), .B2(G197gat), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT127), .ZN(G1352gat));
  NAND2_X1  g818(.A1(new_n981), .A2(new_n1012), .ZN(new_n1020));
  INV_X1    g819(.A(G204gat), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n705), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g821(.A(KEYINPUT62), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OR3_X1    g822(.A1(new_n1020), .A2(KEYINPUT62), .A3(new_n1022), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1025));
  AND2_X1   g824(.A1(new_n1025), .A2(new_n705), .ZN(new_n1026));
  OAI211_X1 g825(.A(new_n1023), .B(new_n1024), .C1(new_n1026), .C2(new_n1021), .ZN(G1353gat));
  OR3_X1    g826(.A1(new_n1020), .A2(G211gat), .A3(new_n885), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1015), .A2(new_n641), .A3(new_n1016), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G1354gat));
  AND2_X1   g831(.A1(new_n1025), .A2(new_n727), .ZN(new_n1033));
  INV_X1    g832(.A(G218gat), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n727), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g834(.A1(new_n1033), .A2(new_n1034), .B1(new_n1020), .B2(new_n1035), .ZN(G1355gat));
endmodule


