

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U555 ( .A1(n528), .A2(G2104), .ZN(n883) );
  NOR2_X2 U556 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X1 U557 ( .A(n657), .B(n656), .ZN(n660) );
  OR2_X1 U558 ( .A1(n692), .A2(n700), .ZN(n520) );
  AND2_X1 U559 ( .A1(n703), .A2(n702), .ZN(n521) );
  AND2_X1 U560 ( .A1(n690), .A2(n994), .ZN(n522) );
  NOR2_X1 U561 ( .A1(n676), .A2(n605), .ZN(n606) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n656) );
  NOR2_X1 U563 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U564 ( .A1(n584), .A2(G651), .ZN(n795) );
  XNOR2_X1 U565 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n523) );
  INV_X1 U566 ( .A(KEYINPUT87), .ZN(n538) );
  XNOR2_X1 U567 ( .A(n524), .B(n523), .ZN(n527) );
  INV_X1 U568 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U569 ( .A1(G101), .A2(n883), .ZN(n524) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U571 ( .A1(G113), .A2(n887), .ZN(n525) );
  XNOR2_X1 U572 ( .A(n525), .B(KEYINPUT66), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n533) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n528), .ZN(n888) );
  NAND2_X1 U575 ( .A1(G125), .A2(n888), .ZN(n531) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n529), .Z(n884) );
  NAND2_X1 U577 ( .A1(G137), .A2(n884), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U579 ( .A1(n533), .A2(n532), .ZN(G160) );
  NAND2_X1 U580 ( .A1(G114), .A2(n887), .ZN(n535) );
  NAND2_X1 U581 ( .A1(G126), .A2(n888), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n541) );
  NAND2_X1 U583 ( .A1(G138), .A2(n884), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G102), .A2(n883), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U586 ( .A(n539), .B(n538), .ZN(n540) );
  NOR2_X1 U587 ( .A1(n541), .A2(n540), .ZN(G164) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n584) );
  NAND2_X1 U589 ( .A1(n795), .A2(G51), .ZN(n542) );
  XNOR2_X1 U590 ( .A(KEYINPUT79), .B(n542), .ZN(n546) );
  XNOR2_X1 U591 ( .A(G651), .B(KEYINPUT67), .ZN(n550) );
  NOR2_X1 U592 ( .A1(G543), .A2(n550), .ZN(n543) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n543), .Z(n794) );
  NAND2_X1 U594 ( .A1(n794), .A2(G63), .ZN(n544) );
  XOR2_X1 U595 ( .A(KEYINPUT78), .B(n544), .Z(n545) );
  NOR2_X1 U596 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U597 ( .A(n547), .B(KEYINPUT6), .ZN(n555) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n548) );
  XNOR2_X1 U599 ( .A(n548), .B(KEYINPUT64), .ZN(n799) );
  NAND2_X1 U600 ( .A1(G89), .A2(n799), .ZN(n549) );
  XNOR2_X1 U601 ( .A(n549), .B(KEYINPUT4), .ZN(n552) );
  NOR2_X1 U602 ( .A1(n584), .A2(n550), .ZN(n798) );
  NAND2_X1 U603 ( .A1(G76), .A2(n798), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U605 ( .A(KEYINPUT5), .B(n553), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U607 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U608 ( .A1(n798), .A2(G77), .ZN(n557) );
  XNOR2_X1 U609 ( .A(n557), .B(KEYINPUT70), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G90), .A2(n799), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U612 ( .A(n560), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U613 ( .A1(G64), .A2(n794), .ZN(n561) );
  NAND2_X1 U614 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U615 ( .A1(G52), .A2(n795), .ZN(n563) );
  XNOR2_X1 U616 ( .A(KEYINPUT69), .B(n563), .ZN(n564) );
  NOR2_X1 U617 ( .A1(n565), .A2(n564), .ZN(G171) );
  NAND2_X1 U618 ( .A1(G78), .A2(n798), .ZN(n566) );
  XNOR2_X1 U619 ( .A(n566), .B(KEYINPUT72), .ZN(n573) );
  NAND2_X1 U620 ( .A1(G65), .A2(n794), .ZN(n568) );
  NAND2_X1 U621 ( .A1(G53), .A2(n795), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U623 ( .A1(G91), .A2(n799), .ZN(n569) );
  XNOR2_X1 U624 ( .A(KEYINPUT71), .B(n569), .ZN(n570) );
  NOR2_X1 U625 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n573), .A2(n572), .ZN(G299) );
  NAND2_X1 U627 ( .A1(n799), .A2(G88), .ZN(n574) );
  XNOR2_X1 U628 ( .A(n574), .B(KEYINPUT82), .ZN(n576) );
  NAND2_X1 U629 ( .A1(n794), .A2(G62), .ZN(n575) );
  NAND2_X1 U630 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U631 ( .A1(G50), .A2(n795), .ZN(n578) );
  NAND2_X1 U632 ( .A1(G75), .A2(n798), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U634 ( .A1(n580), .A2(n579), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G49), .A2(n795), .ZN(n582) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U640 ( .A1(n794), .A2(n583), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n584), .A2(G87), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G73), .A2(n798), .ZN(n587) );
  XNOR2_X1 U644 ( .A(n587), .B(KEYINPUT2), .ZN(n594) );
  NAND2_X1 U645 ( .A1(G61), .A2(n794), .ZN(n589) );
  NAND2_X1 U646 ( .A1(G48), .A2(n795), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U648 ( .A1(G86), .A2(n799), .ZN(n590) );
  XNOR2_X1 U649 ( .A(KEYINPUT81), .B(n590), .ZN(n591) );
  NOR2_X1 U650 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U651 ( .A1(n594), .A2(n593), .ZN(G305) );
  NAND2_X1 U652 ( .A1(n795), .A2(G47), .ZN(n596) );
  NAND2_X1 U653 ( .A1(G85), .A2(n799), .ZN(n595) );
  NAND2_X1 U654 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U655 ( .A1(n798), .A2(G72), .ZN(n597) );
  XOR2_X1 U656 ( .A(KEYINPUT68), .B(n597), .Z(n598) );
  NOR2_X1 U657 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U658 ( .A1(n794), .A2(G60), .ZN(n600) );
  NAND2_X1 U659 ( .A1(n601), .A2(n600), .ZN(G290) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n705) );
  NAND2_X1 U661 ( .A1(G40), .A2(G160), .ZN(n602) );
  XNOR2_X1 U662 ( .A(n602), .B(KEYINPUT88), .ZN(n706) );
  INV_X1 U663 ( .A(n706), .ZN(n603) );
  NAND2_X2 U664 ( .A1(n705), .A2(n603), .ZN(n661) );
  NAND2_X1 U665 ( .A1(G8), .A2(n661), .ZN(n700) );
  NOR2_X1 U666 ( .A1(G2084), .A2(n661), .ZN(n676) );
  NOR2_X1 U667 ( .A1(G1966), .A2(n700), .ZN(n604) );
  XOR2_X1 U668 ( .A(KEYINPUT92), .B(n604), .Z(n678) );
  NAND2_X1 U669 ( .A1(G8), .A2(n678), .ZN(n605) );
  XOR2_X1 U670 ( .A(KEYINPUT30), .B(n606), .Z(n607) );
  NOR2_X1 U671 ( .A1(G168), .A2(n607), .ZN(n613) );
  XOR2_X1 U672 ( .A(G2078), .B(KEYINPUT25), .Z(n941) );
  NOR2_X1 U673 ( .A1(n941), .A2(n661), .ZN(n608) );
  XOR2_X1 U674 ( .A(KEYINPUT94), .B(n608), .Z(n610) );
  XNOR2_X1 U675 ( .A(KEYINPUT93), .B(G1961), .ZN(n964) );
  NAND2_X1 U676 ( .A1(n661), .A2(n964), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n610), .A2(n609), .ZN(n658) );
  NOR2_X1 U678 ( .A1(G171), .A2(n658), .ZN(n611) );
  XNOR2_X1 U679 ( .A(n611), .B(KEYINPUT98), .ZN(n612) );
  XOR2_X1 U680 ( .A(KEYINPUT31), .B(n614), .Z(n674) );
  INV_X1 U681 ( .A(n661), .ZN(n642) );
  NAND2_X1 U682 ( .A1(n642), .A2(G2072), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n615), .B(KEYINPUT27), .ZN(n617) );
  INV_X1 U684 ( .A(G1956), .ZN(n965) );
  NOR2_X1 U685 ( .A1(n965), .A2(n642), .ZN(n616) );
  NOR2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n651) );
  INV_X1 U687 ( .A(G299), .ZN(n998) );
  NOR2_X1 U688 ( .A1(n651), .A2(n998), .ZN(n619) );
  XNOR2_X1 U689 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n655) );
  XNOR2_X1 U691 ( .A(G1996), .B(KEYINPUT96), .ZN(n940) );
  NAND2_X1 U692 ( .A1(n940), .A2(n642), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(KEYINPUT26), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n661), .A2(G1341), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n633) );
  NAND2_X1 U696 ( .A1(n794), .A2(G56), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n623), .B(KEYINPUT14), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G43), .A2(n795), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n631) );
  NAND2_X1 U700 ( .A1(G81), .A2(n799), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT12), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G68), .A2(n798), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U704 ( .A(KEYINPUT13), .B(n629), .Z(n630) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U706 ( .A(KEYINPUT76), .B(n632), .Z(n997) );
  NOR2_X1 U707 ( .A1(n633), .A2(n997), .ZN(n646) );
  NAND2_X1 U708 ( .A1(G79), .A2(n798), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n794), .A2(G66), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G92), .A2(n799), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G54), .A2(n795), .ZN(n636) );
  XNOR2_X1 U713 ( .A(KEYINPUT77), .B(n636), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(KEYINPUT15), .ZN(n1011) );
  INV_X1 U717 ( .A(n1011), .ZN(n771) );
  NOR2_X1 U718 ( .A1(G2067), .A2(n661), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n642), .A2(G1348), .ZN(n643) );
  NOR2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n771), .A2(n647), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n649) );
  OR2_X1 U723 ( .A1(n647), .A2(n771), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT97), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n651), .A2(n998), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n658), .A2(G171), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n675) );
  INV_X1 U731 ( .A(G8), .ZN(n666) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n700), .ZN(n663) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n661), .ZN(n662) );
  NOR2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(G303), .ZN(n665) );
  OR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n668) );
  AND2_X1 U737 ( .A1(n675), .A2(n668), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n674), .A2(n667), .ZN(n672) );
  INV_X1 U739 ( .A(n668), .ZN(n670) );
  AND2_X1 U740 ( .A1(G286), .A2(G8), .ZN(n669) );
  OR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT32), .ZN(n696) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n680) );
  NAND2_X1 U745 ( .A1(G8), .A2(n676), .ZN(n677) );
  AND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n697) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  AND2_X1 U749 ( .A1(n697), .A2(n1001), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n696), .A2(n681), .ZN(n685) );
  INV_X1 U751 ( .A(n1001), .ZN(n683) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n691) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U754 ( .A1(n691), .A2(n682), .ZN(n1002) );
  OR2_X1 U755 ( .A1(n683), .A2(n1002), .ZN(n684) );
  AND2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U757 ( .A1(n700), .A2(n686), .ZN(n687) );
  NOR2_X1 U758 ( .A1(KEYINPUT33), .A2(n687), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT99), .ZN(n690) );
  XOR2_X1 U760 ( .A(G1981), .B(KEYINPUT100), .Z(n689) );
  XNOR2_X1 U761 ( .A(G305), .B(n689), .ZN(n994) );
  NAND2_X1 U762 ( .A1(n691), .A2(KEYINPUT33), .ZN(n692) );
  NAND2_X1 U763 ( .A1(n522), .A2(n520), .ZN(n704) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U765 ( .A(n693), .B(KEYINPUT24), .Z(n694) );
  OR2_X1 U766 ( .A1(n700), .A2(n694), .ZN(n703) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U768 ( .A1(G8), .A2(n695), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n704), .A2(n521), .ZN(n739) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n751) );
  XNOR2_X1 U774 ( .A(G1986), .B(G290), .ZN(n1007) );
  NAND2_X1 U775 ( .A1(n751), .A2(n1007), .ZN(n726) );
  NAND2_X1 U776 ( .A1(G117), .A2(n887), .ZN(n708) );
  NAND2_X1 U777 ( .A1(G129), .A2(n888), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n883), .A2(G105), .ZN(n709) );
  XOR2_X1 U780 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U782 ( .A(n712), .B(KEYINPUT90), .ZN(n714) );
  NAND2_X1 U783 ( .A1(G141), .A2(n884), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n877) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n877), .ZN(n715) );
  XNOR2_X1 U786 ( .A(n715), .B(KEYINPUT91), .ZN(n723) );
  XNOR2_X1 U787 ( .A(KEYINPUT89), .B(G1991), .ZN(n952) );
  NAND2_X1 U788 ( .A1(G95), .A2(n883), .ZN(n717) );
  NAND2_X1 U789 ( .A1(G131), .A2(n884), .ZN(n716) );
  NAND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U791 ( .A1(G107), .A2(n887), .ZN(n719) );
  NAND2_X1 U792 ( .A1(G119), .A2(n888), .ZN(n718) );
  NAND2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U794 ( .A1(n721), .A2(n720), .ZN(n894) );
  NOR2_X1 U795 ( .A1(n952), .A2(n894), .ZN(n722) );
  NOR2_X1 U796 ( .A1(n723), .A2(n722), .ZN(n932) );
  INV_X1 U797 ( .A(n751), .ZN(n724) );
  NOR2_X1 U798 ( .A1(n932), .A2(n724), .ZN(n742) );
  INV_X1 U799 ( .A(n742), .ZN(n725) );
  NAND2_X1 U800 ( .A1(n726), .A2(n725), .ZN(n737) );
  NAND2_X1 U801 ( .A1(G104), .A2(n883), .ZN(n728) );
  NAND2_X1 U802 ( .A1(G140), .A2(n884), .ZN(n727) );
  NAND2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U804 ( .A(KEYINPUT34), .B(n729), .ZN(n734) );
  NAND2_X1 U805 ( .A1(G116), .A2(n887), .ZN(n731) );
  NAND2_X1 U806 ( .A1(G128), .A2(n888), .ZN(n730) );
  NAND2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U808 ( .A(KEYINPUT35), .B(n732), .Z(n733) );
  NOR2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U810 ( .A(KEYINPUT36), .B(n735), .ZN(n899) );
  XNOR2_X1 U811 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  NOR2_X1 U812 ( .A1(n899), .A2(n748), .ZN(n918) );
  NAND2_X1 U813 ( .A1(n751), .A2(n918), .ZN(n745) );
  INV_X1 U814 ( .A(n745), .ZN(n736) );
  NOR2_X1 U815 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U816 ( .A1(n739), .A2(n738), .ZN(n754) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n877), .ZN(n922) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n740) );
  AND2_X1 U819 ( .A1(n952), .A2(n894), .ZN(n914) );
  NOR2_X1 U820 ( .A1(n740), .A2(n914), .ZN(n741) );
  NOR2_X1 U821 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U822 ( .A1(n922), .A2(n743), .ZN(n744) );
  XNOR2_X1 U823 ( .A(n744), .B(KEYINPUT39), .ZN(n746) );
  NAND2_X1 U824 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U825 ( .A(KEYINPUT101), .B(n747), .Z(n749) );
  NAND2_X1 U826 ( .A1(n899), .A2(n748), .ZN(n919) );
  NAND2_X1 U827 ( .A1(n749), .A2(n919), .ZN(n750) );
  NAND2_X1 U828 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U829 ( .A(n752), .B(KEYINPUT102), .ZN(n753) );
  NAND2_X1 U830 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U831 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U832 ( .A(KEYINPUT105), .B(G2446), .Z(n757) );
  XNOR2_X1 U833 ( .A(KEYINPUT103), .B(G2451), .ZN(n756) );
  XNOR2_X1 U834 ( .A(n757), .B(n756), .ZN(n758) );
  XOR2_X1 U835 ( .A(n758), .B(G2430), .Z(n760) );
  XNOR2_X1 U836 ( .A(G1348), .B(G1341), .ZN(n759) );
  XNOR2_X1 U837 ( .A(n760), .B(n759), .ZN(n764) );
  XOR2_X1 U838 ( .A(G2438), .B(G2435), .Z(n762) );
  XNOR2_X1 U839 ( .A(KEYINPUT104), .B(G2454), .ZN(n761) );
  XNOR2_X1 U840 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U841 ( .A(n764), .B(n763), .Z(n766) );
  XNOR2_X1 U842 ( .A(G2443), .B(G2427), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n766), .B(n765), .ZN(n767) );
  AND2_X1 U844 ( .A1(n767), .A2(G14), .ZN(G401) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G860), .ZN(n793) );
  OR2_X1 U847 ( .A1(n793), .A2(n997), .ZN(G153) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  XOR2_X1 U849 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n769) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U851 ( .A(n769), .B(n768), .ZN(G223) );
  INV_X1 U852 ( .A(G223), .ZN(n831) );
  NAND2_X1 U853 ( .A1(n831), .A2(G567), .ZN(n770) );
  XOR2_X1 U854 ( .A(KEYINPUT11), .B(n770), .Z(G234) );
  INV_X1 U855 ( .A(G171), .ZN(G301) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n773) );
  INV_X1 U857 ( .A(G868), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n771), .A2(n775), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(G284) );
  NOR2_X1 U860 ( .A1(G868), .A2(G299), .ZN(n774) );
  XNOR2_X1 U861 ( .A(n774), .B(KEYINPUT80), .ZN(n777) );
  NOR2_X1 U862 ( .A1(n775), .A2(G286), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n793), .A2(G559), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n778), .A2(n1011), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(n997), .A2(G868), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G868), .A2(n1011), .ZN(n780) );
  NOR2_X1 U869 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G123), .A2(n888), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT18), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n883), .A2(G99), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G111), .A2(n887), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G135), .A2(n884), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n913) );
  XNOR2_X1 U879 ( .A(G2096), .B(n913), .ZN(n791) );
  INV_X1 U880 ( .A(G2100), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G559), .A2(n1011), .ZN(n792) );
  XOR2_X1 U883 ( .A(n997), .B(n792), .Z(n810) );
  NAND2_X1 U884 ( .A1(n793), .A2(n810), .ZN(n804) );
  NAND2_X1 U885 ( .A1(G67), .A2(n794), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G55), .A2(n795), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n798), .A2(G80), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G93), .A2(n799), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n812) );
  XOR2_X1 U892 ( .A(n804), .B(n812), .Z(G145) );
  XNOR2_X1 U893 ( .A(G288), .B(KEYINPUT19), .ZN(n806) );
  XNOR2_X1 U894 ( .A(G166), .B(n998), .ZN(n805) );
  XNOR2_X1 U895 ( .A(n806), .B(n805), .ZN(n807) );
  XOR2_X1 U896 ( .A(n812), .B(n807), .Z(n808) );
  XNOR2_X1 U897 ( .A(G305), .B(n808), .ZN(n809) );
  XNOR2_X1 U898 ( .A(n809), .B(G290), .ZN(n904) );
  XNOR2_X1 U899 ( .A(n810), .B(n904), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n811), .A2(G868), .ZN(n814) );
  OR2_X1 U901 ( .A1(G868), .A2(n812), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XOR2_X1 U908 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  XNOR2_X1 U909 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n819) );
  XNOR2_X1 U912 ( .A(KEYINPUT22), .B(n819), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n820), .A2(G96), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n821), .A2(G218), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT83), .ZN(n836) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n836), .ZN(n823) );
  XNOR2_X1 U917 ( .A(KEYINPUT84), .B(n823), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U919 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U920 ( .A1(G108), .A2(n825), .ZN(n837) );
  NAND2_X1 U921 ( .A1(G567), .A2(n837), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n838) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n828) );
  XOR2_X1 U924 ( .A(KEYINPUT85), .B(n828), .Z(n829) );
  NOR2_X1 U925 ( .A1(n838), .A2(n829), .ZN(n835) );
  NAND2_X1 U926 ( .A1(G36), .A2(n835), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n830), .B(KEYINPUT86), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n832) );
  XOR2_X1 U930 ( .A(KEYINPUT106), .B(n832), .Z(n833) );
  NAND2_X1 U931 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n838), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2084), .Z(n840) );
  XNOR2_X1 U942 ( .A(G2090), .B(G2067), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U944 ( .A(n841), .B(G2096), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2072), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2678), .Z(n845) );
  XNOR2_X1 U948 ( .A(KEYINPUT107), .B(G2100), .ZN(n844) );
  XNOR2_X1 U949 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U950 ( .A(n847), .B(n846), .Z(G227) );
  XOR2_X1 U951 ( .A(G1991), .B(G1981), .Z(n849) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1996), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U955 ( .A(G1986), .B(KEYINPUT110), .ZN(n850) );
  XNOR2_X1 U956 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U957 ( .A(G1976), .B(G1971), .Z(n853) );
  XNOR2_X1 U958 ( .A(G1961), .B(G1956), .ZN(n852) );
  XNOR2_X1 U959 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U960 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U961 ( .A(KEYINPUT109), .B(G2474), .ZN(n856) );
  XNOR2_X1 U962 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G124), .A2(n888), .ZN(n860) );
  XOR2_X1 U965 ( .A(KEYINPUT111), .B(n860), .Z(n861) );
  XNOR2_X1 U966 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U967 ( .A1(G136), .A2(n884), .ZN(n862) );
  NAND2_X1 U968 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G112), .A2(n887), .ZN(n865) );
  NAND2_X1 U970 ( .A1(G100), .A2(n883), .ZN(n864) );
  NAND2_X1 U971 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U973 ( .A(KEYINPUT112), .B(n868), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G118), .A2(n887), .ZN(n870) );
  NAND2_X1 U975 ( .A1(G130), .A2(n888), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G106), .A2(n883), .ZN(n872) );
  NAND2_X1 U978 ( .A1(G142), .A2(n884), .ZN(n871) );
  NAND2_X1 U979 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n873), .Z(n874) );
  NOR2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U982 ( .A(G164), .B(n876), .ZN(n898) );
  XNOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U984 ( .A(n877), .B(KEYINPUT113), .ZN(n878) );
  XNOR2_X1 U985 ( .A(n879), .B(n878), .ZN(n882) );
  XOR2_X1 U986 ( .A(G160), .B(n913), .Z(n880) );
  XNOR2_X1 U987 ( .A(G162), .B(n880), .ZN(n881) );
  XOR2_X1 U988 ( .A(n882), .B(n881), .Z(n896) );
  NAND2_X1 U989 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U990 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G115), .A2(n887), .ZN(n890) );
  NAND2_X1 U993 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n924) );
  XNOR2_X1 U997 ( .A(n894), .B(n924), .ZN(n895) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n901), .ZN(G395) );
  XOR2_X1 U1002 ( .A(KEYINPUT114), .B(G286), .Z(n903) );
  XNOR2_X1 U1003 ( .A(G171), .B(n1011), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n906) );
  XOR2_X1 U1005 ( .A(n997), .B(n904), .Z(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n909), .ZN(n910) );
  AND2_X1 U1011 ( .A1(G319), .A2(n910), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(KEYINPUT55), .ZN(n937) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n931) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n923), .Z(n929) );
  XOR2_X1 U1025 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT50), .B(n927), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n934), .B(KEYINPUT115), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n935), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n938), .A2(G29), .ZN(n993) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(G29), .ZN(n962) );
  XNOR2_X1 U1037 ( .A(G2084), .B(G34), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(n939), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n957) );
  XOR2_X1 U1040 ( .A(n940), .B(G32), .Z(n944) );
  XOR2_X1 U1041 ( .A(n941), .B(KEYINPUT116), .Z(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(G27), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT117), .B(n945), .ZN(n947) );
  XOR2_X1 U1045 ( .A(G2072), .B(G33), .Z(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G26), .B(G2067), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(KEYINPUT118), .B(n950), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n951), .A2(G28), .ZN(n954) );
  XOR2_X1 U1051 ( .A(G25), .B(n952), .Z(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n958), .B(KEYINPUT119), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n1022) );
  INV_X1 U1057 ( .A(n1022), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n963), .ZN(n991) );
  XNOR2_X1 U1060 ( .A(G5), .B(n964), .ZN(n979) );
  XOR2_X1 U1061 ( .A(G1966), .B(G21), .Z(n976) );
  XNOR2_X1 U1062 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G20), .B(n965), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(G1348), .Z(n970) );
  XNOR2_X1 U1069 ( .A(G4), .B(n970), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(n974), .B(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(KEYINPUT125), .B(n977), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(G24), .B(G1986), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1078 ( .A(G1976), .B(G23), .Z(n982) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1082 ( .A(KEYINPUT61), .B(n987), .Z(n988) );
  NOR2_X1 U1083 ( .A1(G16), .A2(n988), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(n989), .B(KEYINPUT126), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1026) );
  XNOR2_X1 U1087 ( .A(KEYINPUT56), .B(G16), .ZN(n1021) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G168), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(KEYINPUT57), .B(n996), .ZN(n1019) );
  XOR2_X1 U1091 ( .A(n997), .B(G1341), .Z(n1016) );
  XNOR2_X1 U1092 ( .A(G1956), .B(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(G1971), .A2(G303), .ZN(n999) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1097 ( .A(KEYINPUT120), .B(n1005), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT121), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1100 ( .A(G171), .B(G1961), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(G1348), .B(n1011), .Z(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT122), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(KEYINPUT123), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(KEYINPUT55), .A2(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n1027) );
  XNOR2_X1 U1113 ( .A(n1028), .B(n1027), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

