//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n462), .A2(G136), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n461), .A2(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G162));
  OAI211_X1 g052(.A(G138), .B(new_n463), .C1(new_n459), .C2(new_n460), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n459), .A2(new_n460), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(G126), .A3(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n480), .B1(new_n478), .B2(new_n479), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n479), .B2(new_n478), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G164));
  XNOR2_X1  g065(.A(KEYINPUT5), .B(G543), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n491), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n492));
  INV_X1    g067(.A(G651), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G50), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n499), .A2(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n494), .A2(new_n507), .ZN(G303));
  INV_X1    g083(.A(G303), .ZN(G166));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT7), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n512), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G89), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n505), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(G63), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n491), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g093(.A(G51), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n496), .B2(new_n497), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G51), .B1(new_n491), .B2(new_n517), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n498), .A2(new_n491), .A3(G89), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n527), .ZN(G168));
  NOR2_X1   g103(.A1(new_n502), .A2(new_n501), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  INV_X1    g105(.A(G77), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n522), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT72), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n534), .B1(new_n531), .B2(new_n522), .C1(new_n529), .C2(new_n530), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(G651), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n505), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT73), .B(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n537), .A2(G90), .B1(new_n523), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n491), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n493), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n499), .A2(new_n544), .B1(new_n505), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n523), .A2(G53), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n491), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G91), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n493), .B1(new_n558), .B2(new_n505), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n556), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  NAND2_X1  g136(.A1(new_n537), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n491), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n523), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n491), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n493), .ZN(new_n567));
  INV_X1    g142(.A(G48), .ZN(new_n568));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n499), .A2(new_n568), .B1(new_n505), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT75), .Z(G305));
  INV_X1    g147(.A(G47), .ZN(new_n573));
  INV_X1    g148(.A(G85), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n499), .A2(new_n573), .B1(new_n505), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n491), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n493), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(KEYINPUT77), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G301), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n498), .A2(new_n491), .A3(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n529), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n587), .A2(KEYINPUT78), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(KEYINPUT78), .B1(new_n587), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n585), .B1(new_n595), .B2(new_n584), .ZN(G284));
  AOI21_X1  g171(.A(new_n585), .B1(new_n595), .B2(new_n584), .ZN(G321));
  MUX2_X1   g172(.A(G286), .B(G299), .S(new_n584), .Z(G297));
  MUX2_X1   g173(.A(G286), .B(G299), .S(new_n584), .Z(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n595), .B1(new_n600), .B2(G860), .ZN(G148));
  INV_X1    g176(.A(new_n547), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n594), .A2(G559), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT79), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(G868), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n482), .A2(new_n464), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT80), .B(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n462), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n472), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n463), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G1341), .B(G1348), .Z(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G14), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n630), .A2(new_n633), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  INV_X1    g220(.A(new_n638), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2096), .B(G2100), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n655));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n652), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(new_n654), .ZN(new_n663));
  MUX2_X1   g238(.A(new_n663), .B(new_n662), .S(new_n657), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XOR2_X1   g242(.A(G1981), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n667), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G29), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G26), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT92), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n462), .A2(G140), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT91), .Z(new_n679));
  OAI21_X1  g254(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n680));
  INV_X1    g255(.A(G116), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(G2105), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n472), .B2(G128), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n677), .B1(new_n684), .B2(G29), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2067), .ZN(new_n686));
  NOR2_X1   g261(.A1(G29), .A2(G33), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT25), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n462), .A2(G139), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(new_n463), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n687), .B1(new_n696), .B2(G29), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(G2072), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G20), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT23), .Z(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G299), .B2(G16), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1956), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(G2072), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n686), .A2(new_n698), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G164), .A2(new_n674), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G27), .B2(new_n674), .ZN(new_n707));
  INV_X1    g282(.A(G2078), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n674), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n674), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT29), .B(G2090), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n707), .A2(new_n708), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n709), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n547), .A2(new_n699), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n699), .B2(G19), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT24), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n674), .B1(new_n719), .B2(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(G34), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G160), .B2(G29), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n718), .A2(G1341), .B1(G2084), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(G2084), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n674), .A2(G32), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n462), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n472), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n674), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G28), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n674), .B1(new_n737), .B2(G28), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(new_n738), .B2(new_n739), .C1(new_n618), .C2(new_n674), .ZN(new_n740));
  INV_X1    g315(.A(G1341), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n717), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n723), .A2(new_n724), .A3(new_n734), .A4(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n705), .A2(new_n715), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n699), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1961), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G21), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G168), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1966), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT89), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n595), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT90), .B(G1348), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n744), .A2(new_n748), .A3(new_n752), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n699), .A2(G22), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G166), .B2(new_n699), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1971), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n699), .A2(G23), .ZN(new_n762));
  INV_X1    g337(.A(G288), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n699), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT33), .B(G1976), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n764), .B(new_n765), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n699), .A2(G6), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n571), .B(KEYINPUT75), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n699), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT32), .B(G1981), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n767), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT34), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n674), .A2(G25), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n472), .A2(G119), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT86), .Z(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n779));
  INV_X1    g354(.A(G107), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G2105), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n462), .B2(G131), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n699), .A2(G24), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT87), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G290), .B2(G16), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1986), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(G1986), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT34), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n767), .A2(new_n794), .A3(new_n773), .A4(new_n772), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n793), .A2(KEYINPUT88), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(KEYINPUT88), .B1(new_n793), .B2(new_n795), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n775), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT36), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(new_n775), .C1(new_n796), .C2(new_n797), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n758), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(G311));
  INV_X1    g379(.A(new_n802), .ZN(G150));
  NOR2_X1   g380(.A1(new_n594), .A2(new_n600), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT38), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n537), .A2(G93), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n491), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT97), .B(G55), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(new_n493), .B2(new_n809), .C1(new_n499), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n547), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n807), .B(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n815), .A2(new_n816), .A3(G860), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n811), .A2(G860), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  XNOR2_X1  g395(.A(new_n783), .B(new_n609), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n462), .A2(G142), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n472), .A2(G130), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n463), .A2(G118), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n821), .B(new_n826), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n684), .A2(new_n489), .ZN(new_n828));
  NAND3_X1  g403(.A1(G164), .A2(new_n679), .A3(new_n683), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n696), .ZN(new_n831));
  INV_X1    g406(.A(new_n696), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n832), .A2(new_n828), .A3(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n833), .A3(new_n731), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n731), .B1(new_n831), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n827), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n836), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n821), .B(new_n826), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n840), .A2(new_n841), .A3(new_n834), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT99), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n840), .A2(new_n841), .A3(new_n844), .A4(new_n834), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n827), .B(KEYINPUT98), .C1(new_n835), .C2(new_n836), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n839), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(G160), .B(new_n618), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n476), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n837), .A2(new_n851), .A3(new_n842), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n812), .B(KEYINPUT100), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n605), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n605), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n587), .A2(new_n591), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n556), .A2(new_n559), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n863), .A2(new_n864), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(KEYINPUT41), .A3(new_n865), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n857), .B1(new_n861), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n865), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n861), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n861), .A2(new_n857), .A3(new_n873), .ZN(new_n878));
  XNOR2_X1  g453(.A(G303), .B(G288), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n581), .A2(new_n769), .A3(new_n582), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n769), .B1(new_n581), .B2(new_n582), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n879), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n877), .A2(new_n878), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n877), .B2(new_n878), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n811), .A2(new_n584), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(G331));
  NAND3_X1  g469(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT103), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(G301), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(G168), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n900));
  NAND3_X1  g475(.A1(G168), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n896), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(G168), .B2(new_n897), .ZN(new_n903));
  AOI211_X1 g478(.A(KEYINPUT103), .B(KEYINPUT104), .C1(new_n521), .C2(new_n527), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n895), .A2(G301), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n813), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n899), .A2(new_n896), .A3(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n812), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n887), .B1(new_n873), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n871), .A2(new_n865), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n908), .A2(new_n909), .A3(new_n915), .A4(new_n812), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .A4(new_n907), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n912), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n853), .ZN(new_n922));
  INV_X1    g497(.A(new_n887), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n907), .A2(new_n916), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n914), .A4(new_n913), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n918), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n873), .A2(new_n911), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n913), .A2(new_n916), .A3(new_n907), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n876), .B2(KEYINPUT41), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n914), .A2(new_n933), .A3(new_n862), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n866), .A2(KEYINPUT41), .A3(new_n871), .A4(new_n867), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n907), .A2(new_n914), .A3(new_n910), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT43), .B1(new_n939), .B2(new_n887), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n921), .A3(new_n853), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT108), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n927), .B2(new_n912), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n940), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n930), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(KEYINPUT44), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n939), .A2(new_n887), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n927), .A2(new_n928), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n948), .B(new_n943), .C1(new_n951), .C2(new_n923), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n952), .B2(KEYINPUT109), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n922), .A2(new_n929), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n955), .A3(new_n948), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n947), .B1(KEYINPUT44), .B2(new_n957), .ZN(G397));
  INV_X1    g533(.A(G8), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n489), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n465), .A2(G40), .A3(new_n469), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n486), .B2(new_n488), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(KEYINPUT115), .A2(G2084), .ZN(new_n968));
  AND2_X1   g543(.A1(KEYINPUT115), .A2(G2084), .ZN(new_n969));
  OR3_X1    g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT114), .B(new_n963), .C1(new_n964), .C2(KEYINPUT45), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n751), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n959), .B1(new_n970), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(G168), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT116), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n981), .A3(G168), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1971), .ZN(new_n984));
  INV_X1    g559(.A(new_n974), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n971), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT110), .B(G2090), .Z(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n967), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT111), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n986), .B(new_n991), .C1(new_n967), .C2(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G166), .B2(new_n959), .ZN(new_n994));
  NAND3_X1  g569(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n990), .A2(new_n992), .A3(G8), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n571), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(G1981), .B1(new_n567), .B2(new_n570), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n964), .A2(new_n963), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(KEYINPUT49), .A3(new_n1002), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1005), .A2(G8), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1006), .B(G8), .C1(new_n1009), .C2(G288), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n763), .B2(G1976), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1008), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n999), .A2(KEYINPUT63), .A3(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n990), .A2(G8), .A3(new_n992), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n983), .B(new_n1019), .C1(new_n1020), .C2(new_n996), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT63), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n989), .A2(G8), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n994), .A2(new_n995), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n999), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n980), .B2(new_n982), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1022), .B1(new_n1027), .B2(KEYINPUT117), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(new_n1026), .C1(new_n982), .C2(new_n980), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1021), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1961), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n967), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n708), .A2(KEYINPUT53), .ZN(new_n1034));
  INV_X1    g609(.A(new_n963), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n961), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n708), .A3(new_n974), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1042));
  OAI221_X1 g617(.A(new_n1033), .B1(new_n976), .B2(new_n1034), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(new_n1026), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G168), .A2(new_n959), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT120), .Z(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n978), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1046), .A2(KEYINPUT51), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n978), .B2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n751), .B2(new_n976), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT121), .B(new_n1050), .C1(new_n1054), .C2(new_n959), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1054), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1046), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1056), .A2(KEYINPUT62), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT62), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1045), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n985), .A2(new_n971), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n967), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n556), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n1067), .B2(KEYINPUT118), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(G299), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT61), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .A4(KEYINPUT119), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(new_n999), .A3(new_n1018), .A4(new_n1025), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1006), .A2(G2067), .ZN(new_n1077));
  INV_X1    g652(.A(G1348), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n967), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(KEYINPUT60), .B2(new_n595), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT58), .B(G1341), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n1006), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1037), .A2(new_n974), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(G1996), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n547), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT59), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1069), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT61), .A3(new_n1070), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n594), .B2(new_n1079), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1076), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1098));
  NAND3_X1  g673(.A1(new_n1062), .A2(KEYINPUT53), .A3(new_n708), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1033), .B(new_n1099), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT125), .B1(new_n1100), .B2(G171), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1044), .A2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1100), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1100), .A2(G171), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(KEYINPUT54), .C1(G171), .C2(new_n1043), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1097), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1006), .A2(G8), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1008), .A2(new_n1009), .A3(new_n763), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1001), .ZN(new_n1111));
  INV_X1    g686(.A(new_n999), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1018), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1031), .A2(new_n1061), .A3(new_n1108), .A4(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n684), .B(G2067), .Z(new_n1115));
  XOR2_X1   g690(.A(new_n730), .B(G1996), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n783), .B(new_n785), .Z(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G290), .A2(G1986), .ZN(new_n1120));
  OR2_X1    g695(.A1(G290), .A2(G1986), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n963), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1114), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(KEYINPUT48), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(KEYINPUT48), .B2(new_n1129), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1124), .B1(new_n1115), .B2(new_n731), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT46), .B1(new_n1124), .B2(G1996), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1124), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT47), .Z(new_n1136));
  NAND3_X1  g711(.A1(new_n778), .A2(new_n785), .A3(new_n782), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1117), .A2(new_n1137), .B1(G2067), .B2(new_n684), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1125), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1131), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1127), .A2(new_n1140), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n1143));
  OAI211_X1 g717(.A(new_n650), .B(G319), .C1(new_n635), .C2(new_n636), .ZN(new_n1144));
  NOR2_X1   g718(.A1(G229), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g719(.A(new_n1145), .B(KEYINPUT126), .ZN(new_n1146));
  AOI21_X1  g720(.A(new_n1146), .B1(new_n850), .B2(new_n854), .ZN(new_n1147));
  AND3_X1   g721(.A1(new_n946), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g722(.A(new_n1143), .B1(new_n946), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n1149), .ZN(G308));
  NAND2_X1  g724(.A1(new_n946), .A2(new_n1147), .ZN(G225));
endmodule


