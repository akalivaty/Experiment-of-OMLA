

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n601), .A2(n600), .ZN(n637) );
  INV_X1 U558 ( .A(KEYINPUT94), .ZN(n598) );
  XNOR2_X1 U559 ( .A(n660), .B(n598), .ZN(n644) );
  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n638) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n642) );
  XNOR2_X1 U562 ( .A(n643), .B(n642), .ZN(n649) );
  NOR2_X1 U563 ( .A1(n691), .A2(n690), .ZN(n703) );
  NOR2_X1 U564 ( .A1(n571), .A2(G651), .ZN(n795) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(n529), .Z(n892) );
  NOR2_X1 U566 ( .A1(n540), .A2(n539), .ZN(G164) );
  INV_X1 U567 ( .A(G2105), .ZN(n523) );
  AND2_X1 U568 ( .A1(n523), .A2(G2104), .ZN(n891) );
  NAND2_X1 U569 ( .A1(G101), .A2(n891), .ZN(n524) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n524), .Z(n528) );
  NOR2_X1 U571 ( .A1(n523), .A2(G2104), .ZN(n525) );
  XNOR2_X2 U572 ( .A(n525), .B(KEYINPUT64), .ZN(n897) );
  NAND2_X1 U573 ( .A1(n897), .A2(G125), .ZN(n526) );
  XOR2_X1 U574 ( .A(n526), .B(KEYINPUT65), .Z(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n533) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G137), .A2(n892), .ZN(n531) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U579 ( .A1(G113), .A2(n895), .ZN(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U581 ( .A1(n533), .A2(n532), .ZN(G160) );
  NAND2_X1 U582 ( .A1(n892), .A2(G138), .ZN(n536) );
  NAND2_X1 U583 ( .A1(n897), .A2(G126), .ZN(n534) );
  XOR2_X1 U584 ( .A(n534), .B(KEYINPUT85), .Z(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U586 ( .A1(G102), .A2(n891), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G114), .A2(n895), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n571) );
  NAND2_X1 U590 ( .A1(G52), .A2(n795), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n541), .B(KEYINPUT67), .ZN(n551) );
  NOR2_X1 U592 ( .A1(G543), .A2(G651), .ZN(n799) );
  NAND2_X1 U593 ( .A1(G90), .A2(n799), .ZN(n543) );
  INV_X1 U594 ( .A(G651), .ZN(n545) );
  NOR2_X1 U595 ( .A1(n571), .A2(n545), .ZN(n800) );
  NAND2_X1 U596 ( .A1(G77), .A2(n800), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n544), .B(KEYINPUT9), .ZN(n549) );
  NOR2_X1 U599 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n546), .Z(n547) );
  XNOR2_X1 U601 ( .A(KEYINPUT66), .B(n547), .ZN(n796) );
  NAND2_X1 U602 ( .A1(G64), .A2(n796), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U605 ( .A1(G89), .A2(n799), .ZN(n552) );
  XOR2_X1 U606 ( .A(KEYINPUT71), .B(n552), .Z(n553) );
  XNOR2_X1 U607 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G76), .A2(n800), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n556), .B(KEYINPUT5), .ZN(n562) );
  NAND2_X1 U611 ( .A1(n795), .A2(G51), .ZN(n557) );
  XNOR2_X1 U612 ( .A(n557), .B(KEYINPUT72), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G63), .A2(n796), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U617 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G88), .A2(n799), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G75), .A2(n800), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U622 ( .A(KEYINPUT80), .B(n566), .Z(n570) );
  NAND2_X1 U623 ( .A1(n796), .A2(G62), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n795), .A2(G50), .ZN(n567) );
  AND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(G303) );
  NAND2_X1 U627 ( .A1(G87), .A2(n571), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT78), .ZN(n577) );
  NAND2_X1 U629 ( .A1(G49), .A2(n795), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U632 ( .A1(n796), .A2(n575), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U634 ( .A1(n795), .A2(G48), .ZN(n584) );
  NAND2_X1 U635 ( .A1(G86), .A2(n799), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G61), .A2(n796), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n800), .A2(G73), .ZN(n580) );
  XOR2_X1 U639 ( .A(KEYINPUT2), .B(n580), .Z(n581) );
  NOR2_X1 U640 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U642 ( .A(KEYINPUT79), .B(n585), .Z(G305) );
  NAND2_X1 U643 ( .A1(G85), .A2(n799), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G60), .A2(n796), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U646 ( .A1(G72), .A2(n800), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G47), .A2(n795), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(n590) );
  OR2_X1 U649 ( .A1(n591), .A2(n590), .ZN(G290) );
  NAND2_X1 U650 ( .A1(n795), .A2(G53), .ZN(n593) );
  NAND2_X1 U651 ( .A1(G65), .A2(n796), .ZN(n592) );
  NAND2_X1 U652 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U653 ( .A1(G91), .A2(n799), .ZN(n595) );
  NAND2_X1 U654 ( .A1(G78), .A2(n800), .ZN(n594) );
  NAND2_X1 U655 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U656 ( .A1(n597), .A2(n596), .ZN(n946) );
  AND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n723) );
  NOR2_X1 U658 ( .A1(G164), .A2(G1384), .ZN(n724) );
  NAND2_X1 U659 ( .A1(n723), .A2(n724), .ZN(n660) );
  NAND2_X1 U660 ( .A1(n644), .A2(G2072), .ZN(n599) );
  XNOR2_X1 U661 ( .A(n599), .B(KEYINPUT27), .ZN(n601) );
  INV_X1 U662 ( .A(G1956), .ZN(n972) );
  NOR2_X1 U663 ( .A1(n644), .A2(n972), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n946), .A2(n637), .ZN(n636) );
  NAND2_X1 U665 ( .A1(n660), .A2(G1348), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G2067), .A2(n644), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n603), .A2(n602), .ZN(n628) );
  INV_X1 U668 ( .A(G1996), .ZN(n604) );
  NOR2_X1 U669 ( .A1(n660), .A2(n604), .ZN(n605) );
  XOR2_X1 U670 ( .A(n605), .B(KEYINPUT26), .Z(n607) );
  NAND2_X1 U671 ( .A1(n660), .A2(G1341), .ZN(n606) );
  AND2_X1 U672 ( .A1(n607), .A2(n606), .ZN(n630) );
  NAND2_X1 U673 ( .A1(n799), .A2(G81), .ZN(n608) );
  XNOR2_X1 U674 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U675 ( .A1(G68), .A2(n800), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n612) );
  XOR2_X1 U677 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n611) );
  XNOR2_X1 U678 ( .A(n612), .B(n611), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G56), .A2(n796), .ZN(n613) );
  XOR2_X1 U680 ( .A(KEYINPUT14), .B(n613), .Z(n614) );
  NOR2_X1 U681 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U682 ( .A1(n795), .A2(G43), .ZN(n616) );
  NAND2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n964) );
  INV_X1 U684 ( .A(n964), .ZN(n631) );
  NAND2_X1 U685 ( .A1(G54), .A2(n795), .ZN(n624) );
  NAND2_X1 U686 ( .A1(G79), .A2(n800), .ZN(n619) );
  NAND2_X1 U687 ( .A1(G66), .A2(n796), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G92), .A2(n799), .ZN(n620) );
  XNOR2_X1 U690 ( .A(KEYINPUT69), .B(n620), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(KEYINPUT15), .ZN(n913) );
  AND2_X1 U694 ( .A1(n631), .A2(n913), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n630), .A2(n626), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(KEYINPUT96), .ZN(n634) );
  AND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U699 ( .A1(n632), .A2(n913), .ZN(n633) );
  NAND2_X1 U700 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n641) );
  NOR2_X1 U702 ( .A1(n637), .A2(n946), .ZN(n639) );
  XNOR2_X1 U703 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U704 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U705 ( .A(G2078), .B(KEYINPUT25), .ZN(n930) );
  NAND2_X1 U706 ( .A1(n644), .A2(n930), .ZN(n646) );
  INV_X1 U707 ( .A(G1961), .ZN(n971) );
  NAND2_X1 U708 ( .A1(n971), .A2(n660), .ZN(n645) );
  NAND2_X1 U709 ( .A1(n646), .A2(n645), .ZN(n653) );
  AND2_X1 U710 ( .A1(n653), .A2(G171), .ZN(n647) );
  XNOR2_X1 U711 ( .A(n647), .B(KEYINPUT95), .ZN(n648) );
  NAND2_X1 U712 ( .A1(n649), .A2(n648), .ZN(n658) );
  NAND2_X1 U713 ( .A1(G8), .A2(n660), .ZN(n699) );
  NOR2_X1 U714 ( .A1(G1966), .A2(n699), .ZN(n673) );
  NOR2_X1 U715 ( .A1(G2084), .A2(n660), .ZN(n669) );
  NOR2_X1 U716 ( .A1(n673), .A2(n669), .ZN(n650) );
  NAND2_X1 U717 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U719 ( .A1(G168), .A2(n652), .ZN(n655) );
  NOR2_X1 U720 ( .A1(G171), .A2(n653), .ZN(n654) );
  NOR2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U722 ( .A(KEYINPUT31), .B(n656), .Z(n657) );
  NAND2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n671) );
  NAND2_X1 U724 ( .A1(n671), .A2(G286), .ZN(n659) );
  XOR2_X1 U725 ( .A(KEYINPUT97), .B(n659), .Z(n665) );
  NOR2_X1 U726 ( .A1(G1971), .A2(n699), .ZN(n662) );
  NOR2_X1 U727 ( .A1(G2090), .A2(n660), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n663), .A2(G303), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n666), .B(KEYINPUT98), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(G8), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n668), .B(KEYINPUT32), .ZN(n677) );
  NAND2_X1 U734 ( .A1(G8), .A2(n669), .ZN(n670) );
  XOR2_X1 U735 ( .A(KEYINPUT93), .B(n670), .Z(n675) );
  INV_X1 U736 ( .A(n671), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n694) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n679) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n962) );
  XOR2_X1 U743 ( .A(G1981), .B(G305), .Z(n943) );
  INV_X1 U744 ( .A(n943), .ZN(n682) );
  NAND2_X1 U745 ( .A1(n679), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n699), .A2(n680), .ZN(n681) );
  OR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n686) );
  INV_X1 U748 ( .A(n686), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n683), .A2(KEYINPUT33), .ZN(n689) );
  AND2_X1 U750 ( .A1(n962), .A2(n689), .ZN(n684) );
  AND2_X1 U751 ( .A1(n694), .A2(n684), .ZN(n691) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n947) );
  INV_X1 U753 ( .A(n699), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n947), .A2(n685), .ZN(n687) );
  OR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  AND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U757 ( .A1(G2090), .A2(G303), .ZN(n692) );
  XOR2_X1 U758 ( .A(KEYINPUT99), .B(n692), .Z(n693) );
  NAND2_X1 U759 ( .A1(G8), .A2(n693), .ZN(n695) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n696), .A2(n699), .ZN(n701) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U763 ( .A(n697), .B(KEYINPUT24), .Z(n698) );
  OR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n739) );
  NAND2_X1 U767 ( .A1(G105), .A2(n891), .ZN(n704) );
  XNOR2_X1 U768 ( .A(n704), .B(KEYINPUT88), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(KEYINPUT38), .ZN(n707) );
  NAND2_X1 U770 ( .A1(G117), .A2(n895), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U772 ( .A1(n892), .A2(G141), .ZN(n709) );
  NAND2_X1 U773 ( .A1(G129), .A2(n897), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U776 ( .A(KEYINPUT89), .B(n712), .ZN(n887) );
  NAND2_X1 U777 ( .A1(G1996), .A2(n887), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n713), .B(KEYINPUT90), .ZN(n721) );
  NAND2_X1 U779 ( .A1(G95), .A2(n891), .ZN(n715) );
  NAND2_X1 U780 ( .A1(G107), .A2(n895), .ZN(n714) );
  NAND2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U782 ( .A1(n892), .A2(G131), .ZN(n717) );
  NAND2_X1 U783 ( .A1(G119), .A2(n897), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n874) );
  NAND2_X1 U786 ( .A1(G1991), .A2(n874), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U788 ( .A(KEYINPUT91), .B(n722), .ZN(n1020) );
  INV_X1 U789 ( .A(n1020), .ZN(n726) );
  INV_X1 U790 ( .A(n723), .ZN(n725) );
  NOR2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n755) );
  NAND2_X1 U792 ( .A1(n726), .A2(n755), .ZN(n744) );
  XNOR2_X1 U793 ( .A(KEYINPUT37), .B(G2067), .ZN(n743) );
  NAND2_X1 U794 ( .A1(G104), .A2(n891), .ZN(n728) );
  NAND2_X1 U795 ( .A1(G140), .A2(n892), .ZN(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n730) );
  XOR2_X1 U797 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n729) );
  XNOR2_X1 U798 ( .A(n730), .B(n729), .ZN(n735) );
  NAND2_X1 U799 ( .A1(n895), .A2(G116), .ZN(n732) );
  NAND2_X1 U800 ( .A1(G128), .A2(n897), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U802 ( .A(KEYINPUT35), .B(n733), .Z(n734) );
  NOR2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U804 ( .A(KEYINPUT36), .B(n736), .ZN(n907) );
  NOR2_X1 U805 ( .A1(n743), .A2(n907), .ZN(n1011) );
  NAND2_X1 U806 ( .A1(n755), .A2(n1011), .ZN(n751) );
  NAND2_X1 U807 ( .A1(n744), .A2(n751), .ZN(n737) );
  XNOR2_X1 U808 ( .A(n737), .B(KEYINPUT92), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n742) );
  XNOR2_X1 U810 ( .A(G1986), .B(G290), .ZN(n950) );
  NAND2_X1 U811 ( .A1(n755), .A2(n950), .ZN(n740) );
  XNOR2_X1 U812 ( .A(KEYINPUT86), .B(n740), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n742), .A2(n741), .ZN(n758) );
  NAND2_X1 U814 ( .A1(n743), .A2(n907), .ZN(n1008) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n887), .ZN(n1022) );
  INV_X1 U816 ( .A(n744), .ZN(n747) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n874), .ZN(n1010) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U819 ( .A1(n1010), .A2(n745), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n1022), .A2(n748), .ZN(n749) );
  XNOR2_X1 U822 ( .A(KEYINPUT100), .B(n749), .ZN(n750) );
  XNOR2_X1 U823 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U825 ( .A(KEYINPUT101), .B(n753), .Z(n754) );
  NAND2_X1 U826 ( .A1(n1008), .A2(n754), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U829 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U830 ( .A(G2451), .B(G2435), .ZN(n769) );
  XOR2_X1 U831 ( .A(G2446), .B(KEYINPUT103), .Z(n761) );
  XNOR2_X1 U832 ( .A(G2454), .B(G2430), .ZN(n760) );
  XNOR2_X1 U833 ( .A(n761), .B(n760), .ZN(n765) );
  XOR2_X1 U834 ( .A(KEYINPUT102), .B(G2427), .Z(n763) );
  XNOR2_X1 U835 ( .A(G1341), .B(G1348), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n763), .B(n762), .ZN(n764) );
  XOR2_X1 U837 ( .A(n765), .B(n764), .Z(n767) );
  XNOR2_X1 U838 ( .A(G2443), .B(G2438), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n767), .B(n766), .ZN(n768) );
  XNOR2_X1 U840 ( .A(n769), .B(n768), .ZN(n770) );
  AND2_X1 U841 ( .A1(n770), .A2(G14), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(n946), .ZN(G299) );
  INV_X1 U844 ( .A(G120), .ZN(G236) );
  INV_X1 U845 ( .A(G69), .ZN(G235) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  INV_X1 U848 ( .A(G82), .ZN(G220) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U850 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U851 ( .A(G567), .ZN(n832) );
  NOR2_X1 U852 ( .A1(n832), .A2(G223), .ZN(n772) );
  XNOR2_X1 U853 ( .A(n772), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n778) );
  OR2_X1 U855 ( .A1(n964), .A2(n778), .ZN(G153) );
  INV_X1 U856 ( .A(G171), .ZN(G301) );
  INV_X1 U857 ( .A(n913), .ZN(n952) );
  INV_X1 U858 ( .A(G868), .ZN(n818) );
  NAND2_X1 U859 ( .A1(n952), .A2(n818), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT70), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(G284) );
  NOR2_X1 U863 ( .A1(G286), .A2(n818), .ZN(n777) );
  NOR2_X1 U864 ( .A1(G868), .A2(G299), .ZN(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U866 ( .A1(n778), .A2(G559), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n779), .A2(n913), .ZN(n780) );
  XNOR2_X1 U868 ( .A(n780), .B(KEYINPUT73), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT16), .B(n781), .Z(G148) );
  NOR2_X1 U870 ( .A1(G868), .A2(n964), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n913), .A2(G868), .ZN(n782) );
  NOR2_X1 U872 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G99), .A2(n891), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G111), .A2(n895), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n897), .A2(G123), .ZN(n787) );
  XNOR2_X1 U878 ( .A(n787), .B(KEYINPUT74), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(KEYINPUT18), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G135), .A2(n892), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n1014) );
  XOR2_X1 U883 ( .A(n1014), .B(G2096), .Z(n793) );
  NOR2_X1 U884 ( .A1(G2100), .A2(n793), .ZN(n794) );
  XNOR2_X1 U885 ( .A(KEYINPUT75), .B(n794), .ZN(G156) );
  NAND2_X1 U886 ( .A1(n795), .A2(G55), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G67), .A2(n796), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G93), .A2(n799), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G80), .A2(n800), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U892 ( .A(KEYINPUT77), .B(n803), .Z(n804) );
  OR2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n819) );
  NAND2_X1 U894 ( .A1(G559), .A2(n913), .ZN(n806) );
  XOR2_X1 U895 ( .A(n964), .B(n806), .Z(n815) );
  XOR2_X1 U896 ( .A(n815), .B(KEYINPUT76), .Z(n807) );
  NOR2_X1 U897 ( .A1(G860), .A2(n807), .ZN(n808) );
  XOR2_X1 U898 ( .A(n819), .B(n808), .Z(G145) );
  INV_X1 U899 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U900 ( .A(n819), .B(G166), .ZN(n809) );
  XNOR2_X1 U901 ( .A(n809), .B(G305), .ZN(n810) );
  XNOR2_X1 U902 ( .A(KEYINPUT19), .B(n810), .ZN(n812) );
  XNOR2_X1 U903 ( .A(G288), .B(KEYINPUT81), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U905 ( .A(n813), .B(G290), .ZN(n814) );
  XNOR2_X1 U906 ( .A(n814), .B(G299), .ZN(n910) );
  XNOR2_X1 U907 ( .A(n815), .B(n910), .ZN(n816) );
  XNOR2_X1 U908 ( .A(KEYINPUT82), .B(n816), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n821) );
  NOR2_X1 U910 ( .A1(G868), .A2(n819), .ZN(n820) );
  NOR2_X1 U911 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U913 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U914 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U918 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U919 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U920 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G96), .A2(n828), .ZN(n842) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n842), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n829), .B(KEYINPUT83), .ZN(n834) );
  NOR2_X1 U924 ( .A1(G235), .A2(G236), .ZN(n830) );
  NAND2_X1 U925 ( .A1(G108), .A2(n830), .ZN(n831) );
  NOR2_X1 U926 ( .A1(G237), .A2(n831), .ZN(n844) );
  NOR2_X1 U927 ( .A1(n832), .A2(n844), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(G319) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n836) );
  INV_X1 U930 ( .A(G319), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n837), .B(KEYINPUT84), .ZN(n841) );
  NAND2_X1 U933 ( .A1(G36), .A2(n841), .ZN(G176) );
  INV_X1 U934 ( .A(G223), .ZN(n838) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U937 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U939 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U940 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(n842), .ZN(n843) );
  NAND2_X1 U944 ( .A1(n844), .A2(n843), .ZN(G261) );
  INV_X1 U945 ( .A(G261), .ZN(G325) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1981), .Z(n846) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1956), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n847), .B(KEYINPUT106), .Z(n849) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1961), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U956 ( .A(KEYINPUT105), .B(G2474), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2096), .B(KEYINPUT43), .Z(n857) );
  XNOR2_X1 U959 ( .A(G2090), .B(G2678), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(n858), .B(KEYINPUT104), .Z(n860) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U964 ( .A(KEYINPUT42), .B(G2100), .Z(n862) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U968 ( .A1(G100), .A2(n891), .ZN(n866) );
  NAND2_X1 U969 ( .A1(G112), .A2(n895), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n892), .A2(G136), .ZN(n867) );
  XNOR2_X1 U972 ( .A(KEYINPUT107), .B(n867), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G124), .A2(n897), .ZN(n868) );
  XOR2_X1 U974 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  NOR2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U976 ( .A(KEYINPUT108), .B(n871), .Z(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n874), .B(KEYINPUT112), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n877), .ZN(n889) );
  NAND2_X1 U982 ( .A1(n895), .A2(G118), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G130), .A2(n897), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G106), .A2(n891), .ZN(n881) );
  NAND2_X1 U986 ( .A1(G142), .A2(n892), .ZN(n880) );
  NAND2_X1 U987 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U988 ( .A(KEYINPUT45), .B(n882), .ZN(n883) );
  XNOR2_X1 U989 ( .A(KEYINPUT109), .B(n883), .ZN(n884) );
  NOR2_X1 U990 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U992 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U993 ( .A(G160), .B(n890), .ZN(n906) );
  NAND2_X1 U994 ( .A1(G103), .A2(n891), .ZN(n894) );
  NAND2_X1 U995 ( .A1(G139), .A2(n892), .ZN(n893) );
  NAND2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U997 ( .A1(n895), .A2(G115), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n896), .B(KEYINPUT110), .ZN(n899) );
  NAND2_X1 U999 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1001 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n1004) );
  XOR2_X1 U1003 ( .A(n1004), .B(G162), .Z(n904) );
  XNOR2_X1 U1004 ( .A(G164), .B(n1014), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1009 ( .A(KEYINPUT113), .B(n910), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G171), .B(G286), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n964), .B(n913), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n916), .ZN(G397) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n917) );
  XOR2_X1 U1016 ( .A(KEYINPUT49), .B(n917), .Z(n918) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT114), .B(n920), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1023 ( .A(G2090), .B(G35), .Z(n936) );
  XOR2_X1 U1024 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n934) );
  XNOR2_X1 U1025 ( .A(G1996), .B(G32), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n923) );
  NOR2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n929) );
  XOR2_X1 U1028 ( .A(G1991), .B(G25), .Z(n925) );
  NAND2_X1 U1029 ( .A1(n925), .A2(G28), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(G26), .B(G2067), .ZN(n926) );
  NOR2_X1 U1031 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1033 ( .A(G27), .B(n930), .Z(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(n934), .B(n933), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G34), .B(G2084), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT54), .B(n937), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1040 ( .A(KEYINPUT55), .B(n940), .Z(n942) );
  XOR2_X1 U1041 ( .A(G29), .B(KEYINPUT119), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n1001) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .ZN(n970) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G168), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(n945), .B(KEYINPUT57), .ZN(n968) );
  XNOR2_X1 U1047 ( .A(n946), .B(G1956), .ZN(n948) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n960) );
  AND2_X1 U1049 ( .A1(G303), .A2(G1971), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G171), .B(G1961), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT121), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(G1348), .B(KEYINPUT120), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(n953), .B(n952), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(n956), .B(KEYINPUT122), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1060 ( .A(KEYINPUT123), .B(n963), .Z(n966) );
  XNOR2_X1 U1061 ( .A(G1341), .B(n964), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n999) );
  INV_X1 U1065 ( .A(G16), .ZN(n997) );
  XNOR2_X1 U1066 ( .A(n971), .B(G5), .ZN(n993) );
  XOR2_X1 U1067 ( .A(G1966), .B(G21), .Z(n984) );
  XNOR2_X1 U1068 ( .A(n972), .B(G20), .ZN(n980) );
  XOR2_X1 U1069 ( .A(G1341), .B(G19), .Z(n975) );
  XOR2_X1 U1070 ( .A(G6), .B(KEYINPUT124), .Z(n973) );
  XNOR2_X1 U1071 ( .A(G1981), .B(n973), .ZN(n974) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1073 ( .A(KEYINPUT59), .B(G1348), .Z(n976) );
  XNOR2_X1 U1074 ( .A(G4), .B(n976), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(n981), .B(KEYINPUT125), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n982), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n985) );
  NOR2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n988) );
  XOR2_X1 U1083 ( .A(G1976), .B(G23), .Z(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n989), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1088 ( .A(n994), .B(KEYINPUT126), .ZN(n995) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(n995), .Z(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(G11), .A2(n1002), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(n1003), .B(KEYINPUT127), .ZN(n1031) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT50), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G160), .B(G2084), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT116), .B(n1016), .Z(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1025) );
  XOR2_X1 U1107 ( .A(G2090), .B(G162), .Z(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT51), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1026), .Z(n1027) );
  NOR2_X1 U1112 ( .A1(KEYINPUT55), .A2(n1027), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT117), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(G29), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

