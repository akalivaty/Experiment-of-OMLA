//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n210), .A2(G50), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n209), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  AOI21_X1  g0043(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G97), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n228), .A2(G1698), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G226), .B2(G1698), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n245), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n215), .B1(KEYINPUT68), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G33), .A3(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n244), .A2(new_n253), .B1(new_n261), .B2(G238), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n263));
  INV_X1    g0063(.A(new_n215), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT67), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT67), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n255), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n265), .A2(new_n268), .A3(new_n269), .A4(G274), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n258), .B2(new_n260), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT67), .A2(G41), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT67), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n277), .B2(new_n255), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT69), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n262), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n270), .A2(new_n271), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT69), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(new_n262), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G200), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n281), .A2(new_n290), .A3(new_n286), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT64), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT64), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n296), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n214), .A2(new_n299), .A3(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n300), .A3(G77), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n215), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT11), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(KEYINPUT11), .A3(new_n307), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n269), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OR3_X1    g0116(.A1(new_n316), .A2(KEYINPUT12), .A3(G68), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT12), .B1(new_n316), .B2(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n314), .B2(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n303), .B1(new_n269), .B2(G20), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n310), .A2(new_n311), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT75), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n310), .A2(new_n324), .A3(new_n311), .A4(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n292), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n284), .A2(new_n285), .A3(new_n262), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n285), .B1(new_n284), .B2(new_n262), .ZN(new_n329));
  OAI21_X1  g0129(.A(G169), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT14), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n287), .A2(new_n332), .A3(G169), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n281), .A2(G179), .A3(new_n286), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n331), .B(new_n333), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n326), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n327), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n298), .A2(new_n300), .A3(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n302), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n307), .ZN(new_n346));
  INV_X1    g0146(.A(new_n316), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n202), .B1(new_n269), .B2(G20), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n347), .A2(new_n202), .B1(new_n319), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n261), .A2(G226), .ZN(new_n353));
  MUX2_X1   g0153(.A(G222), .B(G223), .S(G1698), .Z(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n252), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT3), .B(G33), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n244), .B1(new_n356), .B2(G77), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n284), .B(new_n353), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n351), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT72), .B(G179), .Z(new_n360));
  OR2_X1    g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT9), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n350), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n358), .A2(new_n290), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n358), .A2(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n350), .A2(new_n364), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT10), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n365), .B(KEYINPUT74), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n368), .A2(new_n370), .A3(new_n369), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT10), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n363), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n261), .A2(G232), .ZN(new_n378));
  OR2_X1    g0178(.A1(G223), .A2(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G1698), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(G226), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G87), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n381), .A2(new_n252), .B1(new_n250), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n360), .B1(new_n383), .B2(new_n244), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n284), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n244), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n378), .B(new_n388), .C1(new_n272), .C2(new_n279), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n352), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n284), .A2(KEYINPUT79), .A3(new_n378), .A4(new_n384), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n341), .B1(new_n269), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n347), .A2(new_n341), .B1(new_n393), .B2(new_n319), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT77), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n293), .A2(new_n250), .ZN(new_n397));
  INV_X1    g0197(.A(G159), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n302), .A2(KEYINPUT77), .A3(G159), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n399), .A2(new_n400), .B1(new_n401), .B2(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(G20), .B1(new_n249), .B2(new_n251), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n294), .A2(new_n296), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n406), .A2(new_n356), .A3(KEYINPUT7), .ZN(new_n407));
  OAI211_X1 g0207(.A(KEYINPUT16), .B(new_n402), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n408), .A2(new_n307), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT78), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n248), .A3(G33), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n413), .A3(new_n251), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n404), .B1(new_n356), .B2(G20), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n303), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n399), .A2(new_n400), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n401), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n410), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n395), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT18), .B1(new_n392), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n284), .A2(new_n378), .A3(new_n384), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(KEYINPUT79), .B1(new_n352), .B2(new_n389), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n411), .A2(new_n413), .A3(new_n251), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n416), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n420), .B1(new_n429), .B2(G68), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n307), .B(new_n408), .C1(new_n430), .C2(KEYINPUT16), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n394), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n425), .A2(new_n426), .A3(new_n432), .A4(new_n387), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n389), .A2(G200), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n284), .A2(G190), .A3(new_n378), .A4(new_n388), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n431), .A3(new_n394), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n434), .A4(new_n435), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n423), .A2(new_n433), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n356), .A2(G238), .A3(G1698), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n356), .A2(G232), .A3(new_n380), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n356), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n244), .B1(G244), .B2(new_n261), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n284), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n319), .B(G77), .C1(G1), .C2(new_n293), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n342), .A2(new_n302), .B1(new_n406), .B2(G77), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT15), .B(G87), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n297), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G77), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n307), .B1(new_n453), .B2(new_n347), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n446), .A2(G190), .A3(new_n284), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n448), .A2(new_n449), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n352), .ZN(new_n457));
  INV_X1    g0257(.A(new_n360), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n446), .A2(new_n284), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n449), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT73), .ZN(new_n463));
  AND4_X1   g0263(.A1(new_n340), .A2(new_n377), .A3(new_n441), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n306), .A2(new_n215), .B1(G20), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(G33), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n406), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n466), .B(KEYINPUT20), .C1(new_n406), .C2(new_n469), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n472), .A2(new_n473), .B1(new_n465), .B2(new_n347), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n250), .A2(G1), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n307), .C1(new_n314), .C2(new_n315), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT84), .B1(new_n476), .B2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(new_n475), .ZN(new_n478));
  AND4_X1   g0278(.A1(KEYINPUT84), .A2(new_n319), .A3(G116), .A4(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n474), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n269), .B(G45), .C1(new_n482), .C2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n275), .B2(new_n276), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n484), .A2(new_n485), .B1(new_n258), .B2(new_n260), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n266), .A2(new_n267), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n486), .A2(G270), .B1(new_n488), .B2(new_n274), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n249), .A2(new_n251), .A3(G264), .A4(G1698), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n249), .A2(new_n251), .A3(G257), .A4(new_n380), .ZN(new_n491));
  INV_X1    g0291(.A(G303), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n492), .C2(new_n356), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n244), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n481), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n480), .A2(G169), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n480), .A2(KEYINPUT85), .A3(G169), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n489), .A2(new_n494), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n480), .A2(G169), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n489), .A2(G179), .A3(new_n494), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n502), .A2(new_n481), .B1(new_n480), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n480), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(G200), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(new_n290), .C2(new_n501), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n500), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n302), .A2(G77), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n468), .A2(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n468), .A2(new_n444), .A3(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g0313(.A(KEYINPUT80), .B(G107), .Z(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT80), .B(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n512), .A3(new_n511), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n406), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n444), .B1(new_n415), .B2(new_n416), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n510), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n429), .A2(G107), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n307), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n476), .A2(new_n468), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n347), .A2(G97), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(G1698), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n249), .A2(new_n251), .A3(G244), .A4(new_n380), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n467), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n244), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n486), .A2(G257), .B1(new_n488), .B2(new_n274), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n524), .A2(new_n528), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n519), .A2(new_n520), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n518), .A2(new_n510), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n527), .B1(new_n545), .B2(new_n307), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n534), .A2(new_n535), .A3(new_n360), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n352), .B1(new_n534), .B2(new_n535), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n541), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n538), .A2(G169), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n534), .A2(new_n535), .A3(new_n360), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n307), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n518), .A2(new_n510), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(KEYINPUT81), .B2(new_n522), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n554), .B1(new_n556), .B2(new_n543), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n553), .B(KEYINPUT82), .C1(new_n557), .C2(new_n527), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n540), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n319), .A2(G107), .A3(new_n478), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT86), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(KEYINPUT25), .C1(new_n316), .C2(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT86), .B(KEYINPUT25), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n314), .A2(new_n563), .A3(new_n444), .A4(new_n315), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n565), .A2(KEYINPUT87), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(new_n562), .A3(new_n567), .A4(new_n564), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(KEYINPUT23), .A2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n406), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n250), .A2(new_n465), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n293), .B1(new_n572), .B2(KEYINPUT23), .ZN(new_n573));
  NAND2_X1  g0373(.A1(KEYINPUT23), .A2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n214), .A2(new_n356), .A3(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT22), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n214), .A2(new_n356), .A3(new_n578), .A4(G87), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n307), .B1(new_n580), .B2(KEYINPUT24), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(new_n579), .ZN(new_n582));
  INV_X1    g0382(.A(new_n575), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(KEYINPUT24), .A3(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n566), .A2(new_n569), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n486), .A2(G264), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n249), .A2(new_n251), .A3(G257), .A4(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(new_n380), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n244), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n488), .A2(new_n274), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G169), .ZN(new_n594));
  INV_X1    g0394(.A(G179), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(KEYINPUT88), .C1(new_n595), .C2(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT88), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n593), .A2(new_n595), .ZN(new_n598));
  AOI22_X1  g0398(.A1(G264), .A2(new_n486), .B1(new_n590), .B2(new_n244), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n352), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n585), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n249), .A2(new_n251), .A3(G244), .A4(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n249), .A2(new_n251), .A3(G238), .A4(new_n380), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G116), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n255), .A2(G1), .A3(G274), .ZN(new_n607));
  AOI21_X1  g0407(.A(G250), .B1(new_n269), .B2(G45), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n606), .A2(new_n244), .B1(new_n265), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n458), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT83), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n613), .A3(new_n458), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n294), .A2(new_n296), .A3(G33), .A4(G97), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT19), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n214), .A2(new_n356), .A3(G68), .ZN(new_n618));
  NAND3_X1  g0418(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n294), .A2(new_n296), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n382), .A2(new_n468), .A3(new_n444), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n307), .ZN(new_n624));
  INV_X1    g0424(.A(new_n451), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n476), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n347), .A2(new_n451), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n606), .A2(new_n244), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n609), .A2(new_n265), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n352), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n612), .A2(new_n614), .A3(new_n628), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(G200), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n476), .A2(G87), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n610), .A2(G190), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n623), .A2(new_n307), .B1(new_n347), .B2(new_n451), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n593), .A2(new_n288), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(G190), .B2(new_n593), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n582), .A2(new_n583), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT24), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n307), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n565), .A2(KEYINPUT87), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n568), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n602), .A2(new_n639), .A3(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n464), .A2(new_n509), .A3(new_n559), .A4(new_n650), .ZN(G372));
  AND2_X1   g0451(.A1(new_n423), .A2(new_n433), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n292), .A2(new_n326), .ZN(new_n653));
  INV_X1    g0453(.A(new_n461), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n338), .A2(new_n339), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n438), .A2(new_n439), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n372), .B2(new_n376), .ZN(new_n659));
  OAI211_X1 g0459(.A(KEYINPUT90), .B(new_n652), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n363), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n550), .A2(new_n558), .A3(KEYINPUT26), .A4(new_n639), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n547), .B2(new_n548), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n551), .A2(KEYINPUT89), .A3(new_n552), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n524), .A2(new_n528), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n628), .A2(new_n632), .A3(new_n611), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n638), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n585), .B1(new_n600), .B2(new_n598), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n500), .A2(new_n674), .A3(new_n505), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n524), .A2(new_n528), .A3(new_n537), .A4(new_n539), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n676), .A2(new_n649), .A3(new_n669), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n550), .A2(new_n558), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n673), .A2(new_n679), .A3(new_n668), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n464), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n661), .A2(new_n681), .ZN(G369));
  NAND3_X1  g0482(.A1(new_n214), .A2(new_n269), .A3(G13), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n480), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n500), .A2(new_n505), .A3(new_n508), .A4(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n500), .A2(new_n505), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n602), .A2(new_n649), .ZN(new_n695));
  INV_X1    g0495(.A(new_n688), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n646), .B2(new_n648), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n695), .A2(new_n697), .B1(new_n602), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n674), .A2(new_n688), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n688), .B1(new_n500), .B2(new_n505), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n602), .A2(new_n649), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  NAND2_X1  g0504(.A1(new_n277), .A2(new_n207), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n621), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n212), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND3_X1  g0509(.A1(new_n500), .A2(new_n602), .A3(new_n505), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n677), .A3(new_n678), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n668), .ZN(new_n712));
  AND4_X1   g0512(.A1(KEYINPUT26), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n550), .A2(new_n558), .A3(new_n639), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n671), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT29), .B(new_n696), .C1(new_n712), .C2(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n680), .A2(new_n696), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT91), .B(KEYINPUT31), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n696), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n599), .A2(new_n534), .A3(new_n535), .A4(new_n610), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n503), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n610), .A2(new_n360), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n538), .A2(new_n725), .A3(new_n501), .A4(new_n593), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT92), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n599), .A2(new_n610), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n504), .A2(new_n728), .A3(new_n536), .A4(KEYINPUT30), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n724), .A2(KEYINPUT92), .A3(new_n726), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n721), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n724), .A3(new_n726), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n688), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT93), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n735), .A2(new_n739), .A3(new_n736), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n733), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n509), .A2(new_n650), .A3(new_n559), .A4(new_n696), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n719), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n718), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n709), .B1(new_n745), .B2(new_n269), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT94), .Z(G364));
  INV_X1    g0547(.A(new_n692), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n719), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT95), .ZN(new_n750));
  INV_X1    g0550(.A(G13), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n406), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n269), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n705), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(KEYINPUT95), .A3(new_n705), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n749), .A2(new_n693), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT96), .Z(new_n760));
  INV_X1    g0560(.A(new_n758), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n356), .A2(new_n207), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n207), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n239), .A2(G45), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n252), .A2(new_n207), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n213), .B2(new_n255), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n215), .B1(G20), .B2(new_n352), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n761), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  INV_X1    g0576(.A(new_n771), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n692), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G58), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n458), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n214), .A2(new_n290), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n214), .A2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n779), .A2(new_n782), .B1(new_n784), .B2(new_n453), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n458), .A2(new_n288), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n781), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n783), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n202), .A2(new_n787), .B1(new_n788), .B2(new_n303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n288), .A2(G179), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(G20), .A3(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n214), .B1(G190), .B2(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n356), .B1(new_n382), .B2(new_n791), .C1(new_n793), .C2(new_n468), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n785), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  OR3_X1    g0595(.A1(new_n214), .A2(KEYINPUT98), .A3(G190), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT98), .B1(new_n214), .B2(G190), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n796), .A2(new_n797), .A3(new_n792), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n398), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n797), .A3(new_n790), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT99), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n795), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n798), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n802), .A2(G283), .B1(G329), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  INV_X1    g0607(.A(new_n782), .ZN(new_n808));
  INV_X1    g0608(.A(new_n787), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G322), .A2(new_n808), .B1(new_n809), .B2(G326), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT33), .B(G317), .Z(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n811), .B2(new_n793), .C1(new_n788), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n252), .B1(new_n492), .B2(new_n791), .C1(new_n784), .C2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n804), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n776), .B(new_n778), .C1(new_n817), .C2(new_n772), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n760), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  OR3_X1    g0620(.A1(new_n461), .A2(KEYINPUT102), .A3(new_n696), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT102), .B1(new_n461), .B2(new_n696), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n460), .A2(new_n688), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(new_n822), .B1(new_n462), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n717), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n824), .A2(new_n688), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n680), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n743), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT103), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n761), .B1(new_n831), .B2(new_n744), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n772), .ZN(new_n834));
  INV_X1    g0634(.A(new_n784), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G143), .A2(new_n808), .B1(new_n835), .B2(G159), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n837), .B2(new_n787), .C1(new_n838), .C2(new_n788), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT34), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n802), .A2(G68), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n356), .B1(new_n202), .B2(new_n791), .C1(new_n793), .C2(new_n779), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n805), .B2(G132), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n465), .A2(new_n784), .B1(new_n788), .B2(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n811), .A2(new_n782), .B1(new_n787), .B2(new_n492), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n252), .B1(new_n444), .B2(new_n791), .C1(new_n793), .C2(new_n468), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n802), .A2(G87), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(new_n814), .C2(new_n798), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n834), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n772), .A2(new_n769), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT101), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n758), .B(new_n854), .C1(new_n453), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n824), .A2(new_n769), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n833), .A2(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n752), .A2(new_n269), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n408), .A2(new_n307), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n252), .A2(new_n214), .A3(new_n404), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(G68), .C1(new_n404), .C2(new_n403), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT16), .B1(new_n866), .B2(new_n402), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n394), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n686), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n440), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n868), .A2(new_n387), .A3(new_n390), .A4(new_n391), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n436), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n425), .A2(new_n432), .A3(new_n387), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n432), .A2(new_n869), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n436), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n656), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT104), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n652), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n878), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n876), .A2(new_n436), .A3(new_n878), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n885), .A2(new_n886), .B1(new_n879), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n881), .B1(new_n889), .B2(KEYINPUT38), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n334), .B(KEYINPUT76), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n331), .A2(new_n333), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n339), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n323), .A2(new_n325), .A3(new_n688), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n653), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n338), .A2(new_n339), .A3(new_n688), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n824), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n735), .B2(new_n720), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n742), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n872), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n872), .B2(new_n880), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n897), .B(new_n900), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n890), .A2(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n906), .A2(new_n464), .A3(new_n900), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n464), .B2(new_n900), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n719), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT107), .Z(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n461), .A2(new_n688), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n828), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n895), .A2(new_n896), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n872), .A2(new_n880), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n881), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n652), .A2(new_n869), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n893), .A2(new_n688), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n440), .A2(new_n871), .B1(new_n875), .B2(new_n879), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT39), .B1(new_n926), .B2(KEYINPUT38), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n889), .B2(KEYINPUT38), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT39), .B1(new_n902), .B2(new_n903), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n923), .A2(new_n930), .A3(KEYINPUT105), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT105), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n326), .A2(new_n696), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n338), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n340), .B2(new_n894), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n828), .B2(new_n913), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n921), .B1(new_n936), .B2(new_n919), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n884), .A2(new_n423), .A3(new_n433), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT104), .B1(new_n438), .B2(new_n439), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n886), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n888), .A2(new_n879), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n881), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n918), .B2(new_n881), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n924), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n932), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n931), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n464), .B(new_n716), .C1(new_n717), .C2(KEYINPUT29), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n661), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n863), .B1(new_n911), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n911), .B2(new_n952), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n515), .A2(new_n517), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT35), .ZN(new_n957));
  OAI211_X1 g0757(.A(G116), .B(new_n216), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT36), .Z(new_n960));
  OAI21_X1  g0760(.A(G77), .B1(new_n779), .B2(new_n303), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n212), .A2(new_n961), .B1(G50), .B2(new_n303), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n751), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n960), .A3(new_n963), .ZN(G367));
  NAND2_X1  g0764(.A1(new_n637), .A2(new_n635), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n688), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n669), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n668), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n771), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n773), .B1(new_n207), .B2(new_n451), .C1(new_n234), .C2(new_n766), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n761), .A2(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n787), .A2(new_n814), .B1(new_n444), .B2(new_n793), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n791), .A2(new_n975), .A3(new_n465), .ZN(new_n976));
  INV_X1    g0776(.A(new_n791), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT46), .B1(new_n977), .B2(G116), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n976), .A2(new_n356), .A3(new_n978), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n847), .B2(new_n784), .C1(new_n492), .C2(new_n782), .ZN(new_n980));
  INV_X1    g0780(.A(new_n788), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n974), .B(new_n980), .C1(G294), .C2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G317), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n982), .B1(new_n468), .B2(new_n801), .C1(new_n983), .C2(new_n798), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n782), .A2(new_n838), .B1(new_n303), .B2(new_n793), .ZN(new_n985));
  INV_X1    g0785(.A(G143), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n985), .A2(KEYINPUT110), .B1(new_n986), .B2(new_n787), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(KEYINPUT110), .B2(new_n985), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT111), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n252), .B1(new_n977), .B2(G58), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n784), .B2(new_n202), .C1(new_n398), .C2(new_n788), .ZN(new_n991));
  INV_X1    g0791(.A(new_n801), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n991), .B1(G77), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n837), .B2(new_n798), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n984), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n834), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n995), .A2(new_n997), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n971), .B(new_n973), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n970), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n667), .A2(new_n688), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n559), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n546), .B1(new_n664), .B2(new_n665), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n688), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(new_n702), .A3(new_n701), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT42), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n559), .A2(new_n1005), .B1(new_n1007), .B2(new_n688), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(new_n602), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n688), .B1(new_n1013), .B2(new_n678), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1003), .B(new_n1004), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT42), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1010), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1014), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1017), .A2(new_n1018), .A3(new_n1002), .A4(new_n970), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n699), .A2(new_n1012), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1020), .B(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n718), .A2(new_n744), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT109), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n694), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n692), .B2(G330), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n701), .A2(new_n702), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n698), .B2(new_n701), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1026), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n703), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n1033), .B2(new_n1012), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1009), .A2(KEYINPUT45), .A3(new_n703), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT44), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1009), .B2(new_n703), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1012), .A3(KEYINPUT44), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n1040), .A3(new_n699), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n699), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1024), .A2(new_n1031), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1024), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n705), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n754), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1001), .B1(new_n1023), .B2(new_n1050), .ZN(G387));
  NAND2_X1  g0851(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n755), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT114), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT114), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1055), .A3(new_n755), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n1024), .C2(new_n1031), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT113), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n693), .A2(KEYINPUT109), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1030), .B(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1060), .B2(new_n753), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1031), .A2(KEYINPUT113), .A3(new_n754), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n698), .A2(new_n777), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n762), .A2(new_n706), .B1(G107), .B2(new_n207), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n231), .A2(new_n255), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n706), .ZN(new_n1066));
  AOI211_X1 g0866(.A(G45), .B(new_n1066), .C1(G68), .C2(G77), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n341), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n766), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1064), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n761), .B1(new_n1071), .B2(new_n774), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n356), .B1(new_n453), .B2(new_n791), .C1(new_n787), .C2(new_n398), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n202), .A2(new_n782), .B1(new_n788), .B2(new_n341), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n784), .A2(new_n303), .B1(new_n451), .B2(new_n793), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n802), .A2(G97), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n838), .C2(new_n798), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n793), .A2(new_n847), .B1(new_n811), .B2(new_n791), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G311), .A2(new_n981), .B1(new_n809), .B2(G322), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n492), .B2(new_n784), .C1(new_n983), .C2(new_n782), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT49), .Z(new_n1085));
  INV_X1    g0885(.A(G326), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n252), .B1(new_n801), .B2(new_n465), .C1(new_n1086), .C2(new_n798), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1078), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1072), .B1(new_n1088), .B2(new_n772), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1061), .A2(new_n1062), .B1(new_n1063), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1057), .A2(new_n1090), .ZN(G393));
  NAND3_X1  g0891(.A1(new_n1044), .A2(new_n754), .A3(new_n1041), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n242), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n773), .B1(new_n468), .B2(new_n207), .C1(new_n1093), .C2(new_n766), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n761), .A2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n788), .A2(new_n492), .B1(new_n465), .B2(new_n793), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n252), .B1(new_n847), .B2(new_n791), .C1(new_n784), .C2(new_n811), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(G322), .C2(new_n805), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n814), .A2(new_n782), .B1(new_n787), .B2(new_n983), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT52), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1100), .A3(new_n803), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n793), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n981), .A2(G50), .B1(G77), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n356), .C1(new_n341), .C2(new_n784), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n809), .B1(new_n808), .B2(G159), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n852), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n798), .A2(new_n986), .B1(new_n303), .B2(new_n791), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT116), .Z(new_n1111));
  OAI21_X1  g0911(.A(new_n1101), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1095), .B1(new_n777), .B2(new_n1009), .C1(new_n1113), .C2(new_n834), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1092), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1041), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n699), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1116), .A2(new_n1117), .B1(new_n1060), .B2(new_n745), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1045), .A3(new_n755), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT118), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT118), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1045), .A3(new_n1121), .A4(new_n755), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1115), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G390));
  AOI21_X1  g0924(.A(new_n719), .B1(new_n742), .B2(new_n899), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n464), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n661), .A2(new_n950), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n915), .B1(new_n743), .B2(new_n825), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n897), .A2(new_n1125), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n914), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1125), .A2(new_n825), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n935), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n743), .A2(new_n825), .A3(new_n915), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n696), .B(new_n825), .C1(new_n712), .C2(new_n715), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n913), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1127), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n913), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n915), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n940), .A2(new_n941), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n917), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n924), .B1(new_n1141), .B2(new_n881), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n912), .B1(new_n680), .B2(new_n827), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n925), .B1(new_n1144), .B2(new_n935), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n929), .A3(new_n928), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1129), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1134), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1137), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n945), .A2(new_n946), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1151), .A2(new_n1145), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1149), .B1(new_n1152), .B2(new_n1129), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n661), .A2(new_n950), .A3(new_n1126), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1157), .A3(new_n755), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1143), .A2(new_n1146), .A3(new_n1134), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n1147), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1151), .A2(new_n769), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n758), .B1(new_n341), .B2(new_n857), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT119), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n356), .B1(new_n977), .B2(G87), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n784), .A2(new_n468), .B1(KEYINPUT121), .B2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n981), .A2(G107), .B1(G77), .B2(new_n1102), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n465), .B2(new_n782), .C1(new_n847), .C2(new_n787), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(KEYINPUT121), .C2(new_n1164), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n842), .C1(new_n811), .C2(new_n798), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G128), .A2(new_n809), .B1(new_n808), .B2(G132), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n252), .B1(new_n1102), .B2(G159), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n791), .A2(new_n838), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n837), .A2(new_n788), .B1(new_n784), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT120), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G50), .A2(new_n992), .B1(new_n805), .B2(G125), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1169), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1163), .B1(new_n1180), .B2(new_n772), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1160), .A2(new_n754), .B1(new_n1161), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1158), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(G378));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n351), .A2(new_n686), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n377), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n377), .A2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n377), .A2(new_n1188), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n1189), .A3(new_n1185), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n906), .B2(G330), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n915), .A2(new_n900), .A3(new_n825), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n890), .A3(KEYINPUT40), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n915), .A2(new_n900), .A3(new_n825), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n902), .A2(new_n903), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n905), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AND4_X1   g1001(.A1(G330), .A2(new_n1195), .A3(new_n1198), .A4(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1196), .A2(new_n1202), .B1(new_n931), .B2(new_n948), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n1201), .A3(G330), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1195), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(KEYINPUT105), .B1(new_n923), .B2(new_n930), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n937), .A2(new_n947), .A3(new_n932), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1195), .A2(new_n1198), .A3(new_n1201), .A4(G330), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(new_n754), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G33), .A2(G41), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G50), .B(new_n1212), .C1(new_n252), .C2(new_n277), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G125), .A2(new_n809), .B1(new_n981), .B2(G132), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1175), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n808), .A2(G128), .B1(new_n977), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n835), .A2(G137), .B1(G150), .B2(new_n1102), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  XOR2_X1   g1019(.A(KEYINPUT123), .B(G124), .Z(new_n1220));
  OAI221_X1 g1020(.A(new_n1212), .B1(new_n801), .B2(new_n398), .C1(new_n798), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1218), .B2(KEYINPUT59), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1213), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n487), .B(new_n356), .C1(new_n977), .C2(G77), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n801), .B2(new_n779), .C1(new_n847), .C2(new_n798), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT122), .Z(new_n1226));
  OAI22_X1  g1026(.A1(new_n787), .A2(new_n465), .B1(new_n303), .B2(new_n793), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n468), .A2(new_n788), .B1(new_n784), .B2(new_n451), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G107), .C2(new_n808), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(KEYINPUT58), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1223), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT58), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n772), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n758), .B1(new_n202), .B2(new_n857), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n1195), .C2(new_n770), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1211), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1155), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1237), .A2(KEYINPUT57), .A3(new_n1210), .A4(new_n1203), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n755), .ZN(new_n1239));
  AND4_X1   g1039(.A1(new_n1208), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1209), .A2(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1237), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1236), .B1(new_n1239), .B2(new_n1243), .ZN(G375));
  INV_X1    g1044(.A(new_n1154), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1127), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1049), .A3(new_n1156), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n915), .A2(new_n770), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n252), .B1(new_n468), .B2(new_n791), .C1(new_n793), .C2(new_n451), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G107), .A2(new_n835), .B1(new_n981), .B2(G116), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n847), .B2(new_n782), .C1(new_n811), .C2(new_n787), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(G303), .C2(new_n805), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n802), .A2(G77), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n356), .B1(new_n791), .B2(new_n398), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G132), .A2(new_n809), .B1(new_n981), .B2(new_n1215), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n202), .B2(new_n793), .C1(new_n838), .C2(new_n784), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G137), .C2(new_n808), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G58), .A2(new_n992), .B1(new_n805), .B2(G128), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1252), .A2(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n761), .B1(G68), .B2(new_n856), .C1(new_n1259), .C2(new_n834), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1245), .A2(new_n753), .B1(new_n1248), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1247), .A2(new_n1262), .ZN(G381));
  OAI211_X1 g1063(.A(new_n1183), .B(new_n1236), .C1(new_n1239), .C2(new_n1243), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n860), .B1(new_n830), .B2(new_n832), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1001), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n753), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1020), .B(new_n1021), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1267), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1057), .A2(new_n819), .A3(new_n1090), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(G390), .A2(new_n1272), .A3(G381), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1265), .A2(new_n1266), .A3(new_n1271), .A4(new_n1273), .ZN(G407));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G343), .C2(new_n1264), .ZN(G409));
  NAND2_X1  g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1158), .A2(new_n1182), .A3(new_n1211), .A4(new_n1235), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1242), .A2(new_n1049), .A3(new_n1237), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1278), .A2(new_n1279), .B1(G213), .B2(new_n687), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(KEYINPUT60), .B2(new_n1156), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1127), .A2(new_n1131), .A3(KEYINPUT60), .A4(new_n1136), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n755), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G384), .B(new_n1262), .C1(new_n1282), .C2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1156), .A2(KEYINPUT60), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1284), .B1(new_n1286), .B2(new_n1246), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1266), .B1(new_n1287), .B2(new_n1261), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1276), .A2(new_n1280), .A3(new_n1290), .ZN(new_n1291));
  XOR2_X1   g1091(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1276), .A2(new_n1280), .A3(new_n1295), .A4(new_n1290), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n687), .A2(G213), .A3(G2897), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1285), .A2(new_n1288), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT57), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1127), .B1(new_n1160), .B2(new_n1137), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n755), .A3(new_n1238), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1183), .B1(new_n1305), .B2(new_n1236), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1279), .ZN(new_n1307));
  INV_X1    g1107(.A(G213), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1307), .A2(new_n1277), .B1(new_n1308), .B2(G343), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1300), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G393), .A2(G396), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1272), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1123), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(G387), .A2(new_n1123), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G390), .A2(new_n1271), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1318), .A2(new_n1272), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1311), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1317), .A2(new_n1294), .A3(new_n1319), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1306), .A2(new_n1309), .A3(new_n1289), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(KEYINPUT63), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT124), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1300), .B(new_n1325), .C1(new_n1306), .C2(new_n1309), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1291), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1310), .A2(KEYINPUT124), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1324), .A2(new_n1326), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1321), .A2(new_n1330), .ZN(G405));
  OAI21_X1  g1131(.A(new_n1289), .B1(new_n1265), .B2(new_n1306), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1276), .A2(new_n1264), .A3(new_n1290), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1320), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1320), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1334), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AOI211_X1 g1137(.A(KEYINPUT126), .B(new_n1320), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


