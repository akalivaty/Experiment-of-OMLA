//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987;
  AND2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G169gat), .B2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G183gat), .B(G190gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n204), .B(new_n210), .C1(new_n203), .C2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT28), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n219), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n202), .B1(KEYINPUT26), .B2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n221), .A2(new_n224), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n219), .A2(G183gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n215), .A2(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n232), .A2(new_n233), .A3(new_n210), .A4(new_n204), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G226gat), .A2(G233gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n235), .A2(KEYINPUT71), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT71), .B1(new_n235), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G197gat), .B(G204gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n245));
  INV_X1    g044(.A(G211gat), .ZN(new_n246));
  INV_X1    g045(.A(G218gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G211gat), .B(G218gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n240), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT72), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT37), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n239), .A2(new_n258), .A3(new_n251), .A4(new_n254), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G8gat), .B(G36gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT73), .ZN(new_n262));
  XNOR2_X1  g061(.A(G64gat), .B(G92gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n251), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n239), .A2(new_n252), .A3(new_n254), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT37), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT38), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n256), .A3(new_n259), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT37), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(KEYINPUT38), .A3(new_n264), .A4(new_n260), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT0), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT81), .ZN(new_n280));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT78), .B(G155gat), .Z(new_n282));
  INV_X1    g081(.A(G162gat), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT2), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G148gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(G141gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(KEYINPUT76), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294));
  AND2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n283), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT77), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n284), .A2(new_n293), .A3(new_n297), .A4(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n295), .B2(new_n296), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n304), .A3(new_n300), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(KEYINPUT2), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n292), .A2(G148gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n286), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n307), .B1(new_n306), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n302), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(G127gat), .A2(G134gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT65), .B(G134gat), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G113gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G120gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329));
  AND2_X1   g128(.A1(G127gat), .A2(G134gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n329), .C1(new_n314), .C2(new_n330), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n318), .A2(new_n320), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n330), .A2(new_n314), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n336), .A2(new_n326), .A3(new_n329), .A4(new_n328), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(KEYINPUT79), .C1(new_n320), .C2(new_n318), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n313), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n320), .ZN(new_n340));
  INV_X1    g139(.A(G134gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G134gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n314), .B1(new_n345), .B2(G127gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n329), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(new_n335), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n340), .A2(new_n346), .B1(new_n348), .B2(new_n326), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n349), .B(new_n302), .C1(new_n311), .C2(new_n312), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n281), .B1(new_n339), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n280), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT74), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n304), .B1(new_n299), .B2(new_n300), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n310), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT78), .B(G155gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(G162gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n297), .A2(new_n301), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n358), .A2(new_n359), .B1(new_n364), .B2(new_n293), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n350), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n281), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n334), .A2(new_n338), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n302), .B(new_n372), .C1(new_n311), .C2(new_n312), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n374), .A2(new_n281), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n365), .B2(new_n349), .ZN(new_n378));
  INV_X1    g177(.A(new_n350), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(KEYINPUT4), .B2(new_n379), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n353), .A2(new_n369), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n350), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n349), .A3(new_n377), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR4_X1   g185(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT5), .A4(new_n367), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n279), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(new_n281), .A3(new_n374), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT81), .B1(new_n368), .B2(KEYINPUT5), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n280), .B(new_n352), .C1(new_n366), .C2(new_n367), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n386), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n352), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n278), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n394), .ZN(new_n398));
  INV_X1    g197(.A(new_n396), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n279), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n271), .A2(new_n264), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n274), .A2(new_n397), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT39), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n367), .C1(new_n382), .C2(new_n386), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n281), .B1(new_n393), .B2(new_n374), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT39), .B1(new_n366), .B2(new_n367), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(new_n278), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT40), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n398), .A2(new_n279), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n271), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  INV_X1    g211(.A(new_n264), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n408), .A2(new_n409), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n271), .B2(new_n264), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n402), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n410), .A2(new_n414), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT3), .B1(new_n251), .B2(new_n236), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n420), .A2(new_n365), .ZN(new_n421));
  INV_X1    g220(.A(G228gat), .ZN(new_n422));
  INV_X1    g221(.A(G233gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n365), .B2(new_n372), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n421), .B(new_n424), .C1(new_n251), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G22gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n251), .B1(new_n373), .B2(new_n236), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n420), .A2(new_n365), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n428), .A2(new_n429), .B1(new_n422), .B2(new_n423), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G78gat), .B(G106gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT31), .B(G50gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n426), .A2(new_n430), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G22gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n439), .A2(KEYINPUT83), .A3(new_n431), .A4(new_n436), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n419), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n397), .A2(new_n400), .B1(new_n417), .B2(new_n414), .ZN(new_n445));
  AND4_X1   g244(.A1(KEYINPUT83), .A2(new_n439), .A3(new_n431), .A4(new_n436), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n433), .A2(new_n436), .B1(new_n439), .B2(new_n431), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n214), .A2(new_n234), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT67), .A3(new_n332), .A4(new_n229), .ZN(new_n454));
  INV_X1    g253(.A(G227gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n423), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n332), .A2(KEYINPUT67), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n337), .B(new_n458), .C1(new_n320), .C2(new_n318), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n235), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n461), .A2(new_n469), .A3(KEYINPUT32), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n465), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n464), .B1(new_n461), .B2(KEYINPUT32), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n468), .A2(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT34), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n460), .ZN(new_n475));
  INV_X1    g274(.A(new_n456), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g276(.A(KEYINPUT34), .B(new_n456), .C1(new_n454), .C2(new_n460), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n452), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(new_n470), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n479), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n479), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n480), .B1(new_n487), .B2(new_n452), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n451), .B1(new_n488), .B2(KEYINPUT36), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n481), .A2(new_n479), .A3(new_n482), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n452), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n480), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT36), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n490), .A2(new_n491), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT36), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n448), .B2(new_n487), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n443), .A2(new_n496), .A3(KEYINPUT84), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n445), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n445), .A3(new_n504), .A4(new_n443), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n450), .A2(new_n498), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n507));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT85), .B(G197gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT11), .B(G169gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT12), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(G1gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT16), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(G1gat), .B2(new_n516), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI221_X1 g322(.A(new_n519), .B1(new_n520), .B2(new_n515), .C1(G1gat), .C2(new_n516), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT90), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  INV_X1    g328(.A(G43gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n531));
  XOR2_X1   g330(.A(G43gat), .B(G50gat), .Z(new_n532));
  OAI211_X1 g331(.A(new_n529), .B(new_n531), .C1(new_n532), .C2(KEYINPUT87), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  INV_X1    g336(.A(G29gat), .ZN(new_n538));
  INV_X1    g337(.A(G36gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT88), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n533), .A2(new_n535), .A3(new_n536), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n536), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n535), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n546), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(new_n546), .B2(new_n553), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n526), .B(new_n528), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n546), .A2(new_n553), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n557), .A2(new_n525), .B1(G229gat), .B2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n514), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n558), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n557), .B(new_n525), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT13), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT18), .B1(new_n556), .B2(new_n558), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n514), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n513), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n562), .A2(new_n513), .A3(new_n566), .ZN(new_n574));
  AOI211_X1 g373(.A(KEYINPUT92), .B(KEYINPUT18), .C1(new_n556), .C2(new_n558), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n507), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n513), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n566), .B(new_n562), .C1(new_n569), .C2(new_n514), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n569), .A2(new_n514), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n574), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n569), .A2(new_n572), .ZN(new_n583));
  INV_X1    g382(.A(new_n575), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT93), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n506), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G57gat), .B(G64gat), .Z(new_n590));
  INV_X1    g389(.A(G71gat), .ZN(new_n591));
  INV_X1    g390(.A(G78gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n590), .B1(KEYINPUT9), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n594), .B(new_n595), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n525), .B1(KEYINPUT21), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n600), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT94), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n603), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n554), .B2(new_n555), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT95), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n624));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  OAI22_X1  g424(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n617), .B(new_n618), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n557), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n622), .A2(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n624), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n610), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n596), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n627), .A2(new_n601), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n640), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n650), .A3(new_n642), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n627), .A2(new_n601), .A3(KEYINPUT10), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n648), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n647), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n653), .B2(new_n643), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT98), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n659), .B(new_n656), .C1(new_n653), .C2(new_n643), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n655), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n639), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n589), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n397), .A2(new_n400), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT99), .B(G1gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1324gat));
  NAND2_X1  g467(.A1(new_n417), .A2(new_n414), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n515), .B2(new_n670), .ZN(new_n673));
  MUX2_X1   g472(.A(new_n672), .B(new_n673), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g473(.A1(new_n498), .A2(KEYINPUT100), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n494), .A2(KEYINPUT70), .B1(KEYINPUT36), .B2(new_n496), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n489), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n664), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n492), .A2(new_n493), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n664), .B2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n664), .A2(new_n443), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n610), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n661), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n638), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n589), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n665), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n538), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n506), .B2(new_n638), .ZN(new_n696));
  INV_X1    g495(.A(new_n638), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n444), .A2(new_n449), .B1(new_n676), .B2(new_n489), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n445), .A2(new_n504), .A3(new_n443), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n488), .A2(new_n699), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n697), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n581), .A2(new_n585), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n665), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n694), .A2(new_n707), .ZN(G1328gat));
  NOR3_X1   g507(.A1(new_n690), .A2(G36gat), .A3(new_n669), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT101), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G36gat), .B1(new_n706), .B2(new_n669), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(G1329gat));
  OAI21_X1  g516(.A(G43gat), .B1(new_n706), .B2(new_n498), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n690), .A2(G43gat), .A3(new_n681), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n679), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n702), .A2(new_n722), .A3(new_n705), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n719), .B1(new_n723), .B2(G43gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n721), .B1(new_n724), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n702), .A2(new_n448), .A3(new_n705), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n443), .A2(G50gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT103), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n726), .A2(G50gat), .B1(new_n691), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n450), .A2(new_n498), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n503), .A2(new_n505), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n639), .A2(new_n703), .A3(new_n661), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n692), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n737), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n741), .A2(new_n669), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743));
  INV_X1    g542(.A(new_n669), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT49), .B(G64gat), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n736), .A2(new_n744), .A3(new_n737), .A4(new_n745), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n742), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1333gat));
  NAND3_X1  g548(.A1(new_n738), .A2(new_n591), .A3(new_n488), .ZN(new_n750));
  OAI21_X1  g549(.A(G71gat), .B1(new_n741), .B2(new_n679), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1334gat));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n443), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(new_n592), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n610), .A2(new_n703), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n661), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n696), .A2(new_n701), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n696), .A2(KEYINPUT106), .A3(new_n701), .A4(new_n761), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n692), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n733), .A2(new_n697), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n760), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT107), .B1(new_n768), .B2(KEYINPUT51), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n760), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n506), .A2(new_n638), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(KEYINPUT107), .A3(KEYINPUT51), .A4(new_n759), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n692), .A2(new_n614), .A3(new_n662), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n766), .A2(new_n614), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI21_X1  g577(.A(G92gat), .B1(new_n762), .B2(new_n669), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n669), .A2(G92gat), .A3(new_n661), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n778), .B(new_n779), .C1(new_n775), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n744), .A3(new_n765), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n771), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n783), .A2(G92gat), .B1(new_n785), .B2(new_n780), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n786), .B2(new_n778), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n764), .A2(new_n722), .A3(new_n765), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G99gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n681), .A2(G99gat), .A3(new_n661), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n769), .B2(new_n774), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT108), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n789), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1338gat));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  OAI21_X1  g596(.A(G106gat), .B1(new_n762), .B2(new_n443), .ZN(new_n798));
  INV_X1    g597(.A(G106gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n448), .A2(new_n662), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n797), .B(new_n798), .C1(new_n775), .C2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n764), .A2(new_n448), .A3(new_n765), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n800), .B(KEYINPUT109), .Z(new_n803));
  AOI22_X1  g602(.A1(new_n802), .A2(G106gat), .B1(new_n785), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n797), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n744), .A2(new_n665), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n651), .A2(new_n652), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n640), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n651), .A2(new_n649), .A3(new_n652), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n812));
  AOI21_X1  g611(.A(new_n647), .B1(new_n653), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n655), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(new_n817), .A3(new_n703), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n557), .A2(new_n525), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n564), .B1(new_n556), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n563), .A2(new_n565), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n512), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n585), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n661), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n638), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n816), .A2(new_n814), .A3(new_n655), .ZN(new_n826));
  INV_X1    g625(.A(new_n823), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n697), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n610), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n639), .A2(new_n703), .A3(new_n662), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n831), .A2(KEYINPUT111), .A3(new_n448), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT111), .B1(new_n831), .B2(new_n448), .ZN(new_n833));
  AOI211_X1 g632(.A(new_n681), .B(new_n807), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n323), .B1(new_n834), .B2(new_n587), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n831), .A2(new_n807), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n500), .A2(new_n501), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n838), .A2(new_n323), .A3(new_n703), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n835), .A2(KEYINPUT112), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT112), .B1(new_n835), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1340gat));
  AOI21_X1  g641(.A(G120gat), .B1(new_n838), .B2(new_n662), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n661), .A2(new_n321), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n834), .B2(new_n844), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n317), .A3(new_n610), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n834), .A2(new_n610), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n317), .ZN(G1342gat));
  NAND3_X1  g647(.A1(new_n838), .A2(new_n316), .A3(new_n697), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT56), .Z(new_n850));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n697), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(G134gat), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT113), .B(new_n341), .C1(new_n834), .C2(new_n697), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n498), .A2(new_n806), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT114), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n824), .B1(new_n587), .B2(new_n826), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n828), .B1(new_n858), .B2(new_n697), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n830), .B1(new_n859), .B2(new_n687), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n860), .B2(new_n443), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n829), .A2(new_n830), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n448), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G141gat), .B1(new_n865), .B2(new_n588), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n836), .A2(new_n448), .A3(new_n679), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n588), .A2(G141gat), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT58), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n857), .A2(new_n703), .A3(new_n864), .A4(new_n861), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n871), .A2(G141gat), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT115), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n870), .B1(new_n875), .B2(new_n877), .ZN(G1344gat));
  NAND4_X1  g677(.A1(new_n867), .A2(new_n288), .A3(new_n290), .A4(new_n662), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT116), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n857), .A2(new_n662), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT93), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT93), .B1(new_n581), .B2(new_n585), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n826), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n824), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n697), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n828), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n687), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n663), .A2(new_n588), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n443), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT117), .B1(new_n890), .B2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n859), .A2(new_n687), .B1(new_n588), .B2(new_n663), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n892), .B(new_n863), .C1(new_n893), .C2(new_n443), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n448), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n285), .B1(new_n881), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT118), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n898), .B(new_n291), .C1(new_n865), .C2(new_n661), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n897), .A2(KEYINPUT118), .A3(new_n898), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n880), .B1(new_n901), .B2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(new_n361), .B1(new_n865), .B2(new_n687), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n867), .A2(new_n282), .A3(new_n610), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n867), .A2(new_n283), .A3(new_n697), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT119), .Z(new_n908));
  OAI21_X1  g707(.A(G162gat), .B1(new_n865), .B2(new_n638), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n831), .A2(new_n692), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n837), .A2(new_n744), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT120), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n206), .A3(new_n703), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n832), .A2(new_n833), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n692), .A2(new_n669), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n681), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n588), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n916), .B1(new_n922), .B2(new_n206), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT121), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n925), .B(new_n916), .C1(new_n922), .C2(new_n206), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1348gat));
  OAI21_X1  g726(.A(G176gat), .B1(new_n921), .B2(new_n661), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n915), .A2(new_n207), .A3(new_n662), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n921), .B2(new_n687), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n610), .A2(new_n222), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n915), .A2(new_n933), .B1(new_n934), .B2(KEYINPUT60), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(KEYINPUT60), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n936), .B(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n915), .A2(new_n219), .A3(new_n697), .ZN(new_n940));
  OAI21_X1  g739(.A(G190gat), .B1(new_n921), .B2(new_n638), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  INV_X1    g743(.A(new_n678), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n677), .B1(new_n676), .B2(new_n489), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n744), .B(new_n448), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n679), .A2(new_n949), .A3(new_n744), .A4(new_n448), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n948), .A2(new_n911), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n703), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n896), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT124), .A4(new_n895), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n722), .A2(new_n919), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n587), .A2(G197gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  INV_X1    g761(.A(G204gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n957), .A2(new_n662), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n661), .A2(G204gat), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n948), .A2(new_n950), .A3(new_n911), .A4(new_n967), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n962), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n968), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n964), .B1(new_n954), .B2(new_n955), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n972), .B(KEYINPUT125), .C1(new_n963), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n951), .A2(new_n246), .A3(new_n610), .ZN(new_n976));
  OAI21_X1  g775(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n722), .A2(new_n687), .A3(new_n919), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n896), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  AOI21_X1  g781(.A(G218gat), .B1(new_n951), .B2(new_n697), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n697), .A2(G218gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n958), .B2(KEYINPUT127), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n956), .A2(new_n986), .A3(new_n957), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n983), .B1(new_n985), .B2(new_n987), .ZN(G1355gat));
endmodule


