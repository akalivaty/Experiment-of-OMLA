//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G128), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n191), .C1(KEYINPUT1), .C2(new_n195), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT80), .A2(G104), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT80), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n203), .A2(KEYINPUT3), .A3(G107), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(KEYINPUT3), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n200), .A2(new_n201), .ZN(new_n209));
  AOI21_X1  g023(.A(G101), .B1(new_n209), .B2(G107), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n208), .A2(KEYINPUT81), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT81), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n197), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT10), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  INV_X1    g029(.A(new_n207), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT80), .A2(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT80), .A2(G104), .ZN(new_n218));
  AOI21_X1  g032(.A(G107), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(G107), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n198), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n215), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n208), .A2(KEYINPUT81), .A3(new_n210), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT10), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n197), .A4(new_n206), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n232), .A2(new_n234), .A3(new_n239), .A4(new_n235), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(KEYINPUT65), .A3(G131), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n216), .B(new_n222), .C1(new_n219), .C2(new_n220), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G101), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n211), .B2(new_n212), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n192), .A2(KEYINPUT64), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n249), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n198), .B1(new_n208), .B2(new_n222), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n244), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n248), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n248), .B1(new_n247), .B2(new_n258), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n229), .B(new_n243), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n264));
  INV_X1    g078(.A(new_n197), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n263), .B(new_n243), .C1(new_n266), .C2(new_n213), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n213), .ZN(new_n268));
  INV_X1    g082(.A(new_n243), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT12), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n262), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT77), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT78), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G227), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT79), .ZN(new_n278));
  INV_X1    g092(.A(new_n276), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n274), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT79), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n229), .B1(new_n260), .B2(new_n261), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n269), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n262), .A3(new_n280), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n262), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n247), .A2(new_n258), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT82), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n259), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n243), .B1(new_n294), .B2(new_n229), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n277), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n262), .A2(KEYINPUT84), .A3(new_n280), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n243), .B1(new_n266), .B2(new_n213), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT12), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT84), .B1(new_n262), .B2(new_n280), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n289), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n293), .A2(new_n259), .B1(new_n214), .B2(new_n228), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n277), .B1(new_n305), .B2(new_n243), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n271), .A2(new_n283), .B1(new_n306), .B2(new_n286), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT83), .B(G469), .C1(new_n307), .C2(G902), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n290), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  OAI21_X1  g124(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n316), .C1(G119), .C2(new_n195), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G110), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT71), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n321), .A3(G125), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n320), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n188), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(KEYINPUT16), .ZN(new_n334));
  OAI211_X1 g148(.A(G146), .B(new_n329), .C1(new_n334), .C2(new_n320), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(G119), .B(G128), .Z(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n319), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n328), .A2(new_n330), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT73), .A3(G146), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n188), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n338), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n317), .B2(G110), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n341), .A2(new_n343), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT74), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n339), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(KEYINPUT75), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n354));
  INV_X1    g168(.A(new_n350), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n349), .A2(new_n355), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n339), .B2(new_n347), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G217), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(G234), .B2(new_n303), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n364), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT25), .B1(new_n361), .B2(new_n303), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n339), .A2(new_n347), .ZN(new_n372));
  INV_X1    g186(.A(new_n359), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n351), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n374), .B(new_n303), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n303), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT76), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n367), .B1(new_n371), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(G237), .A2(G953), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G210), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT27), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT26), .B(G101), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n251), .A2(new_n255), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n241), .A3(new_n242), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n231), .A2(G137), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n233), .A2(G134), .ZN(new_n393));
  OAI21_X1  g207(.A(G131), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n240), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n197), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT2), .B(G113), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT67), .B1(new_n314), .B2(G116), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT67), .ZN(new_n400));
  INV_X1    g214(.A(G116), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(G119), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n401), .A2(G119), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT66), .B(new_n398), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n398), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n399), .B2(new_n402), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT66), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n397), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n391), .A2(new_n410), .A3(new_n396), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n389), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n389), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n388), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n387), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n197), .B2(new_n395), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n391), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n391), .A3(KEYINPUT68), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n410), .B1(new_n397), .B2(new_n419), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n418), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT31), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n417), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT68), .B1(new_n420), .B2(new_n391), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n420), .A2(new_n391), .A3(KEYINPUT68), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n418), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT69), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT69), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n436), .A3(new_n428), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n429), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G472), .A2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT70), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n433), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n391), .A2(new_n410), .A3(new_n396), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n410), .B1(new_n391), .B2(new_n396), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT28), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n415), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n443), .A2(KEYINPUT31), .B1(new_n447), .B2(new_n388), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n434), .A2(KEYINPUT69), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n436), .B1(new_n427), .B2(new_n428), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n439), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n441), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G472), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n387), .A3(new_n415), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n432), .A2(new_n413), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n456), .B(new_n457), .C1(new_n459), .C2(new_n387), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n456), .A2(new_n457), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G902), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n455), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n438), .A2(new_n440), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(KEYINPUT32), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n382), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n197), .A2(new_n323), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n323), .B2(new_n256), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n275), .A2(G224), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT87), .Z(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT88), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n469), .B(new_n472), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n257), .A2(new_n244), .B1(new_n405), .B2(new_n409), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n247), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n205), .B1(new_n224), .B2(new_n225), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g291(.A(G113), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT5), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n404), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n477), .A2(new_n480), .B1(new_n407), .B2(new_n406), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n247), .A2(new_n474), .B1(new_n476), .B2(new_n481), .ZN(new_n487));
  INV_X1    g301(.A(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT6), .ZN(new_n490));
  NOR4_X1   g304(.A1(new_n487), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n488), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n475), .B2(new_n482), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n473), .B(new_n490), .C1(new_n491), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n471), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n469), .B(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n488), .B2(new_n487), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n485), .B(KEYINPUT8), .Z(new_n501));
  INV_X1    g315(.A(new_n482), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n476), .A2(new_n481), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n496), .B2(new_n505), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n467), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n336), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n275), .A3(G214), .ZN(new_n515));
  NOR2_X1   g329(.A1(KEYINPUT89), .A2(G143), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n383), .B(G214), .C1(KEYINPUT89), .C2(G143), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n513), .B(new_n239), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n239), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n519), .B1(new_n523), .B2(KEYINPUT92), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n521), .A2(new_n525), .A3(new_n513), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n331), .A2(new_n335), .A3(KEYINPUT91), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n512), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n203), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT90), .B1(new_n333), .B2(new_n188), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n333), .A2(new_n188), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT18), .A2(G131), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n520), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n322), .A2(new_n324), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT19), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n521), .A2(new_n522), .B1(new_n542), .B2(new_n188), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n341), .A2(new_n343), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  INV_X1    g359(.A(new_n530), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n537), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G475), .A2(G902), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT93), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n510), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT20), .B(new_n550), .C1(new_n537), .C2(new_n547), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n528), .A2(new_n536), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n546), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n555), .B2(new_n537), .ZN(new_n556));
  INV_X1    g370(.A(G475), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n552), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n537), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n530), .B1(new_n528), .B2(new_n536), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n303), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G475), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n564), .B(KEYINPUT94), .C1(new_n552), .C2(new_n553), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n195), .A2(G143), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n190), .A2(G128), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n231), .ZN(new_n569));
  XNOR2_X1  g383(.A(G116), .B(G122), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G107), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n401), .A2(KEYINPUT14), .A3(G122), .ZN(new_n574));
  OAI211_X1 g388(.A(G107), .B(new_n574), .C1(new_n571), .C2(KEYINPUT14), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT13), .B1(new_n190), .B2(G128), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT95), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n567), .B1(KEYINPUT13), .B2(new_n566), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n231), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n231), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n570), .A2(new_n199), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n572), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n576), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n310), .A2(new_n363), .A3(G953), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n576), .B(new_n585), .C1(new_n580), .C2(new_n583), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(KEYINPUT96), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n303), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT15), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n589), .A2(new_n303), .A3(new_n591), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(G952), .A3(new_n275), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT21), .B(G898), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n595), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n560), .A2(new_n565), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n509), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n312), .A2(new_n466), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  OAI21_X1  g422(.A(G472), .B1(new_n438), .B2(G902), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n441), .A2(new_n609), .A3(new_n453), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n309), .A3(new_n381), .A4(new_n311), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n560), .A2(new_n565), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n589), .A2(new_n613), .A3(new_n591), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n587), .A2(KEYINPUT33), .A3(new_n588), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n593), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n592), .A2(new_n593), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n467), .B(new_n603), .C1(new_n507), .C2(new_n508), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n611), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  OR3_X1    g438(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT97), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT97), .B1(new_n552), .B2(new_n553), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n625), .A2(new_n626), .A3(new_n564), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n595), .A2(new_n597), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n611), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT35), .B(G107), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n359), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(new_n339), .A3(new_n347), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n637), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n372), .B1(new_n639), .B2(new_n635), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n380), .A2(new_n371), .B1(new_n641), .B2(new_n365), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n605), .A2(new_n509), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n312), .A2(new_n610), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  OAI21_X1  g460(.A(new_n599), .B1(new_n602), .B2(G900), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n629), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n467), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n496), .A2(new_n505), .ZN(new_n651));
  INV_X1    g465(.A(new_n506), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n642), .B1(new_n454), .B2(new_n465), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n312), .A2(new_n649), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XNOR2_X1  g472(.A(new_n647), .B(KEYINPUT39), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n312), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n638), .A2(new_n640), .A3(new_n365), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n378), .A2(KEYINPUT76), .A3(new_n379), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n364), .B1(new_n378), .B2(KEYINPUT76), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n458), .A2(new_n387), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n444), .A2(new_n445), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n668), .B2(new_n388), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n455), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n464), .B2(KEYINPUT32), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n666), .B1(new_n454), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n653), .A2(new_n654), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n612), .A2(new_n628), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n650), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n661), .A2(new_n662), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n190), .ZN(G45));
  NOR2_X1   g493(.A1(new_n620), .A2(new_n648), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n312), .A2(new_n655), .A3(new_n656), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  AOI21_X1  g496(.A(new_n280), .B1(new_n286), .B2(new_n262), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n270), .A2(new_n267), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n306), .B2(KEYINPUT84), .ZN(new_n685));
  INV_X1    g499(.A(new_n301), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(G469), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n311), .A3(new_n304), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n620), .A2(new_n621), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n688), .A2(KEYINPUT99), .A3(new_n311), .A4(new_n304), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n466), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n629), .A2(new_n621), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n691), .A2(new_n697), .A3(new_n466), .A4(new_n693), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NAND2_X1  g513(.A1(new_n454), .A2(new_n465), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n691), .A2(new_n700), .A3(new_n643), .A4(new_n693), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  AND2_X1   g516(.A1(new_n691), .A2(new_n693), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n435), .A2(new_n437), .ZN(new_n704));
  AOI21_X1  g518(.A(G902), .B1(new_n704), .B2(new_n448), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT100), .B1(new_n705), .B2(new_n455), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n707), .B(G472), .C1(new_n438), .C2(G902), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n451), .A2(new_n439), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n708), .A3(new_n709), .A4(new_n381), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n675), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n612), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n621), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n703), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AND4_X1   g532(.A1(new_n709), .A2(new_n706), .A3(new_n666), .A4(new_n708), .ZN(new_n719));
  INV_X1    g533(.A(new_n619), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n560), .B2(new_n565), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(new_n655), .A3(new_n647), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n691), .A2(new_n719), .A3(new_n722), .A4(new_n693), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  OAI21_X1  g538(.A(G469), .B1(new_n307), .B2(G902), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n304), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n311), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n650), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n507), .A2(new_n508), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n466), .A2(new_n731), .A3(new_n680), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n709), .A2(new_n442), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n733), .B(new_n382), .C1(new_n465), .C2(new_n734), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n721), .A2(new_n726), .A3(new_n730), .A4(new_n647), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n732), .A2(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n239), .ZN(G33));
  AND3_X1   g552(.A1(new_n649), .A2(new_n466), .A3(new_n731), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n231), .ZN(G36));
  AND3_X1   g554(.A1(new_n617), .A2(KEYINPUT104), .A3(new_n618), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT104), .B1(new_n617), .B2(new_n618), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n560), .A3(new_n565), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(KEYINPUT105), .A3(new_n745), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n612), .A2(new_n720), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT43), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n746), .A2(new_n747), .B1(new_n750), .B2(KEYINPUT43), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n610), .A2(new_n642), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n507), .A2(new_n508), .A3(new_n650), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n289), .A2(new_n303), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT103), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n284), .A2(new_n287), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n307), .A2(KEYINPUT103), .A3(KEYINPUT45), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n307), .B2(KEYINPUT45), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT46), .B(new_n764), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(new_n763), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n775), .A3(new_n304), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n311), .A3(new_n659), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n311), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n311), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n680), .A2(new_n382), .A3(new_n762), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n700), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NOR2_X1   g603(.A1(G952), .A2(G953), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n700), .A2(new_n381), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n606), .A2(new_n311), .A3(new_n309), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n610), .A2(new_n311), .A3(new_n309), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n606), .A2(new_n666), .ZN(new_n796));
  OAI22_X1  g610(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n560), .A2(new_n565), .A3(new_n628), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n620), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n621), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n611), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n792), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n621), .B1(new_n620), .B2(new_n798), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n312), .A2(new_n381), .A3(new_n804), .A4(new_n610), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n607), .A3(new_n644), .A4(KEYINPUT107), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n791), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n731), .A2(new_n719), .A3(new_n680), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n700), .A2(new_n311), .A3(new_n309), .A4(new_n666), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n628), .A2(new_n648), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n627), .A2(new_n762), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n653), .A2(new_n467), .A3(new_n654), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n625), .A2(new_n564), .A3(new_n626), .A4(new_n811), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT108), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n808), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n737), .A2(new_n817), .A3(new_n739), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n807), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n714), .A2(new_n715), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n691), .A3(new_n800), .A4(new_n693), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n710), .B(KEYINPUT101), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n698), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n694), .A2(new_n701), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n694), .A2(new_n701), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n717), .A3(KEYINPUT112), .A4(new_n698), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n727), .B(new_n648), .C1(new_n304), .C2(new_n725), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n821), .A2(new_n655), .A3(new_n672), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n657), .A2(new_n831), .A3(new_n681), .A4(new_n723), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT109), .B1(new_n832), .B2(new_n834), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n831), .A2(new_n681), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n657), .A2(new_n723), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT109), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n819), .B(new_n829), .C1(new_n837), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n832), .B(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n803), .A2(new_n806), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n824), .A2(new_n825), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n818), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n791), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  XOR2_X1   g663(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n837), .A2(new_n843), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n791), .B1(new_n853), .B2(new_n848), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n846), .A2(new_n847), .A3(new_n818), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n832), .B(new_n834), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT111), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n852), .B1(new_n861), .B2(KEYINPUT54), .ZN(new_n862));
  INV_X1    g676(.A(new_n599), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n752), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n691), .A2(new_n693), .A3(new_n762), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n382), .B1(new_n465), .B2(new_n734), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT48), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n864), .A2(new_n823), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n655), .A3(new_n703), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n275), .A2(G952), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n454), .A2(new_n671), .A3(new_n381), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n863), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n873), .B1(new_n876), .B2(new_n721), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n866), .A2(KEYINPUT48), .A3(new_n867), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n870), .A2(new_n872), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n688), .A2(new_n727), .A3(new_n304), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT115), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n783), .A2(new_n784), .A3(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n864), .A2(new_n823), .A3(new_n813), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n674), .A2(new_n467), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n871), .A2(new_n885), .A3(new_n703), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n599), .B1(new_n755), .B2(new_n749), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n703), .A3(new_n712), .A4(new_n886), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT50), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n612), .A2(new_n619), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n866), .A2(new_n719), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n884), .A2(new_n887), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n879), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n887), .A3(new_n890), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n892), .A2(new_n887), .A3(KEYINPUT116), .A4(new_n890), .ZN(new_n899));
  INV_X1    g713(.A(new_n880), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n883), .B1(new_n785), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(KEYINPUT51), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n895), .A2(new_n902), .A3(KEYINPUT117), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT117), .B1(new_n895), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n790), .B1(new_n862), .B2(new_n905), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n674), .A2(new_n612), .A3(new_n720), .A4(new_n729), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n688), .A2(new_n304), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT49), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n909), .A3(new_n874), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT118), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n858), .A2(new_n860), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n835), .A2(new_n836), .ZN(new_n914));
  INV_X1    g728(.A(new_n843), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n916), .B2(new_n855), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT54), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n895), .A2(new_n902), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n895), .A2(new_n902), .A3(KEYINPUT117), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n918), .A2(new_n851), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n790), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n910), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n912), .A2(new_n927), .ZN(G75));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n829), .A2(new_n818), .A3(new_n807), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n849), .B1(new_n853), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(G210), .A3(G902), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT119), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n490), .B1(new_n491), .B2(new_n495), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n473), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(KEYINPUT56), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n932), .B2(KEYINPUT119), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n929), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n932), .A2(KEYINPUT119), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(KEYINPUT120), .A3(new_n933), .A4(new_n938), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n275), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n932), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n937), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n940), .A2(new_n942), .A3(new_n946), .ZN(G51));
  NAND2_X1  g761(.A1(new_n931), .A2(G902), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n948), .A2(new_n770), .A3(new_n771), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n930), .B1(new_n914), .B2(new_n915), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n849), .A2(new_n850), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT121), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n850), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n931), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n844), .A2(new_n955), .A3(new_n849), .A4(new_n850), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n763), .B(KEYINPUT57), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n687), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n949), .B1(new_n959), .B2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  INV_X1    g775(.A(new_n958), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n851), .A2(KEYINPUT121), .B1(new_n931), .B2(new_n953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n956), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(new_n687), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n943), .B1(new_n960), .B2(new_n965), .ZN(G54));
  INV_X1    g780(.A(new_n948), .ZN(new_n967));
  AND2_X1   g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n967), .A2(new_n548), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n548), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n943), .ZN(G60));
  NAND2_X1  g785(.A1(new_n614), .A2(new_n615), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT59), .Z(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n862), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n972), .A2(new_n974), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n943), .B1(new_n957), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(G63));
  INV_X1    g792(.A(new_n931), .ZN(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n641), .ZN(new_n983));
  INV_X1    g797(.A(new_n943), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n361), .B(KEYINPUT123), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n979), .B2(new_n981), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G66));
  AOI21_X1  g803(.A(new_n275), .B1(new_n601), .B2(G224), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n846), .A2(new_n847), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n275), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT125), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n935), .B1(G898), .B2(new_n275), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(G69));
  NAND2_X1  g810(.A1(new_n840), .A2(new_n681), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n678), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n466), .A2(new_n762), .A3(new_n799), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n660), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n785), .B2(new_n787), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT62), .B1(new_n678), .B2(new_n997), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n998), .A2(new_n779), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n275), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n397), .A2(new_n419), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n425), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(new_n542), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(G900), .B2(G953), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n997), .A2(new_n737), .A3(new_n739), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n778), .A2(new_n655), .A3(new_n821), .A4(new_n867), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n779), .A2(new_n1010), .A3(new_n788), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1009), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT126), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1008), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G72));
  INV_X1    g834(.A(new_n861), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n459), .A2(new_n388), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  NAND3_X1  g838(.A1(new_n1022), .A2(new_n667), .A3(new_n1024), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1012), .A2(new_n992), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n1026), .A2(new_n1024), .ZN(new_n1027));
  OAI221_X1 g841(.A(new_n984), .B1(new_n1021), .B2(new_n1025), .C1(new_n1027), .C2(new_n1022), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1024), .B1(new_n1003), .B2(new_n992), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n387), .A3(new_n458), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT127), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1028), .A2(new_n1031), .ZN(G57));
endmodule


