

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U324 ( .A1(n500), .A2(n499), .ZN(n501) );
  NOR2_X1 U325 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U326 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n292) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U328 ( .A(n413), .B(n293), .ZN(n414) );
  XNOR2_X1 U329 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U330 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U331 ( .A(n423), .B(n422), .ZN(n425) );
  NOR2_X1 U332 ( .A1(n569), .A2(n561), .ZN(n553) );
  XNOR2_X1 U333 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n447) );
  XOR2_X1 U334 ( .A(G1GAT), .B(KEYINPUT34), .Z(n445) );
  XOR2_X1 U335 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n295) );
  XNOR2_X1 U336 ( .A(G197GAT), .B(G218GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(KEYINPUT21), .B(n296), .Z(n339) );
  XOR2_X1 U339 ( .A(G22GAT), .B(G155GAT), .Z(n382) );
  XOR2_X1 U340 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n298) );
  XNOR2_X1 U341 ( .A(G141GAT), .B(KEYINPUT86), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n366) );
  XOR2_X1 U343 ( .A(n382), .B(n366), .Z(n300) );
  NAND2_X1 U344 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n339), .B(n301), .ZN(n314) );
  XOR2_X1 U347 ( .A(KEYINPUT23), .B(KEYINPUT82), .Z(n303) );
  XNOR2_X1 U348 ( .A(G204GAT), .B(G211GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U350 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n305) );
  XNOR2_X1 U351 ( .A(KEYINPUT24), .B(KEYINPUT83), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n307), .B(n306), .Z(n312) );
  XOR2_X1 U354 ( .A(G78GAT), .B(KEYINPUT71), .Z(n309) );
  XNOR2_X1 U355 ( .A(G148GAT), .B(G106GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n417) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G162GAT), .Z(n310) );
  XOR2_X1 U358 ( .A(KEYINPUT75), .B(n310), .Z(n396) );
  XNOR2_X1 U359 ( .A(n417), .B(n396), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n548) );
  XOR2_X1 U362 ( .A(G71GAT), .B(G176GAT), .Z(n316) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G99GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U365 ( .A(n317), .B(G190GAT), .Z(n319) );
  XOR2_X1 U366 ( .A(G15GAT), .B(G127GAT), .Z(n391) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(n391), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U369 ( .A(KEYINPUT65), .B(KEYINPUT80), .Z(n321) );
  XNOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT81), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(n323), .B(n322), .Z(n328) );
  XOR2_X1 U373 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n325) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n345) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(G120GAT), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n326), .B(KEYINPUT0), .ZN(n363) );
  XNOR2_X1 U378 ( .A(n345), .B(n363), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U380 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n330) );
  NAND2_X1 U381 ( .A1(G227GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(KEYINPUT79), .B(n331), .Z(n332) );
  XOR2_X1 U384 ( .A(n333), .B(n332), .Z(n513) );
  NAND2_X1 U385 ( .A1(n548), .A2(n513), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n334), .B(KEYINPUT94), .ZN(n335) );
  XOR2_X1 U387 ( .A(KEYINPUT26), .B(n335), .Z(n527) );
  XOR2_X1 U388 ( .A(G92GAT), .B(G64GAT), .Z(n337) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(KEYINPUT73), .B(n338), .Z(n424) );
  XNOR2_X1 U392 ( .A(n424), .B(n339), .ZN(n349) );
  XOR2_X1 U393 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n341) );
  NAND2_X1 U394 ( .A1(G226GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n342), .B(G211GAT), .ZN(n387) );
  XOR2_X1 U398 ( .A(n343), .B(n387), .Z(n347) );
  XNOR2_X1 U399 ( .A(G36GAT), .B(G190GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n344), .B(KEYINPUT77), .ZN(n397) );
  XNOR2_X1 U401 ( .A(n345), .B(n397), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U403 ( .A(n349), .B(n348), .Z(n541) );
  XNOR2_X1 U404 ( .A(n541), .B(KEYINPUT27), .ZN(n376) );
  NAND2_X1 U405 ( .A1(n527), .A2(n376), .ZN(n354) );
  INV_X1 U406 ( .A(n513), .ZN(n551) );
  AND2_X1 U407 ( .A1(n551), .A2(n541), .ZN(n350) );
  NOR2_X1 U408 ( .A1(n548), .A2(n350), .ZN(n351) );
  XOR2_X1 U409 ( .A(n351), .B(KEYINPUT95), .Z(n352) );
  XNOR2_X1 U410 ( .A(KEYINPUT25), .B(n352), .ZN(n353) );
  NAND2_X1 U411 ( .A1(n354), .A2(n353), .ZN(n375) );
  XOR2_X1 U412 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n356) );
  XNOR2_X1 U413 ( .A(KEYINPUT91), .B(KEYINPUT1), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n374) );
  XOR2_X1 U415 ( .A(G57GAT), .B(G148GAT), .Z(n358) );
  XNOR2_X1 U416 ( .A(G127GAT), .B(G85GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n360) );
  XNOR2_X1 U419 ( .A(G155GAT), .B(KEYINPUT4), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U421 ( .A(n362), .B(n361), .Z(n372) );
  XOR2_X1 U422 ( .A(KEYINPUT89), .B(n363), .Z(n365) );
  NAND2_X1 U423 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U425 ( .A(n366), .B(G162GAT), .Z(n368) );
  XOR2_X1 U426 ( .A(G113GAT), .B(G1GAT), .Z(n426) );
  XNOR2_X1 U427 ( .A(G29GAT), .B(n426), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n487) );
  INV_X1 U432 ( .A(n487), .ZN(n545) );
  NAND2_X1 U433 ( .A1(n375), .A2(n545), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n548), .B(KEYINPUT28), .ZN(n494) );
  INV_X1 U435 ( .A(n494), .ZN(n515) );
  NAND2_X1 U436 ( .A1(n376), .A2(n487), .ZN(n511) );
  NOR2_X1 U437 ( .A1(n551), .A2(n511), .ZN(n377) );
  NAND2_X1 U438 ( .A1(n515), .A2(n377), .ZN(n378) );
  NAND2_X1 U439 ( .A1(n379), .A2(n378), .ZN(n454) );
  XOR2_X1 U440 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n381) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n385) );
  XNOR2_X1 U443 ( .A(G64GAT), .B(G78GAT), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U445 ( .A(n385), .B(n384), .Z(n389) );
  XNOR2_X1 U446 ( .A(G71GAT), .B(G57GAT), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n292), .B(n386), .ZN(n415) );
  XNOR2_X1 U448 ( .A(n415), .B(n387), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U451 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XOR2_X1 U452 ( .A(n393), .B(n392), .Z(n578) );
  INV_X1 U453 ( .A(n578), .ZN(n536) );
  XOR2_X1 U454 ( .A(G29GAT), .B(G43GAT), .Z(n395) );
  XNOR2_X1 U455 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n427) );
  XNOR2_X1 U457 ( .A(n427), .B(n396), .ZN(n410) );
  XOR2_X1 U458 ( .A(n397), .B(G218GAT), .Z(n399) );
  XOR2_X1 U459 ( .A(G99GAT), .B(G85GAT), .Z(n413) );
  XNOR2_X1 U460 ( .A(G134GAT), .B(n413), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n401) );
  NAND2_X1 U463 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U465 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U466 ( .A(KEYINPUT66), .B(KEYINPUT76), .Z(n405) );
  XNOR2_X1 U467 ( .A(G92GAT), .B(G106GAT), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n406), .B(KEYINPUT10), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n538) );
  INV_X1 U472 ( .A(n538), .ZN(n562) );
  NAND2_X1 U473 ( .A1(n536), .A2(n562), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT16), .B(n411), .Z(n412) );
  AND2_X1 U475 ( .A1(n454), .A2(n412), .ZN(n474) );
  XOR2_X1 U476 ( .A(n416), .B(KEYINPUT31), .Z(n423) );
  XNOR2_X1 U477 ( .A(n417), .B(KEYINPUT32), .ZN(n421) );
  XOR2_X1 U478 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n419) );
  XNOR2_X1 U479 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n471) );
  INV_X1 U482 ( .A(n471), .ZN(n504) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U484 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U486 ( .A(G8GAT), .B(KEYINPUT30), .Z(n431) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(KEYINPUT67), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n435) );
  XNOR2_X1 U491 ( .A(G50GAT), .B(G36GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U493 ( .A(G15GAT), .B(G22GAT), .Z(n437) );
  XNOR2_X1 U494 ( .A(G197GAT), .B(G141GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n529) );
  INV_X1 U498 ( .A(n529), .ZN(n569) );
  NOR2_X1 U499 ( .A1(n504), .A2(n569), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n442), .B(KEYINPUT74), .ZN(n459) );
  NAND2_X1 U501 ( .A1(n474), .A2(n459), .ZN(n443) );
  XOR2_X1 U502 ( .A(KEYINPUT96), .B(n443), .Z(n452) );
  NAND2_X1 U503 ( .A1(n452), .A2(n487), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(G1324GAT) );
  NAND2_X1 U506 ( .A1(n452), .A2(n541), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n448), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U508 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n450) );
  NAND2_X1 U509 ( .A1(n452), .A2(n551), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U511 ( .A(G15GAT), .B(n451), .Z(G1326GAT) );
  NAND2_X1 U512 ( .A1(n452), .A2(n494), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT101), .B(KEYINPUT37), .Z(n458) );
  NAND2_X1 U515 ( .A1(n578), .A2(n454), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT100), .B(n455), .Z(n456) );
  XNOR2_X1 U517 ( .A(KEYINPUT36), .B(n538), .ZN(n581) );
  NAND2_X1 U518 ( .A1(n456), .A2(n581), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n484) );
  NAND2_X1 U520 ( .A1(n459), .A2(n484), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT38), .B(n460), .Z(n468) );
  NAND2_X1 U522 ( .A1(n468), .A2(n487), .ZN(n463) );
  XOR2_X1 U523 ( .A(G29GAT), .B(KEYINPUT39), .Z(n461) );
  XNOR2_X1 U524 ( .A(KEYINPUT102), .B(n461), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n463), .B(n462), .ZN(G1328GAT) );
  NAND2_X1 U526 ( .A1(n468), .A2(n541), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n464), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U528 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n466) );
  NAND2_X1 U529 ( .A1(n468), .A2(n551), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U531 ( .A(G43GAT), .B(n467), .ZN(G1330GAT) );
  XNOR2_X1 U532 ( .A(G50GAT), .B(KEYINPUT104), .ZN(n470) );
  NAND2_X1 U533 ( .A1(n494), .A2(n468), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(G1331GAT) );
  XNOR2_X1 U535 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n477) );
  INV_X1 U536 ( .A(KEYINPUT41), .ZN(n472) );
  XNOR2_X1 U537 ( .A(n472), .B(n471), .ZN(n497) );
  XOR2_X1 U538 ( .A(n497), .B(KEYINPUT105), .Z(n555) );
  NOR2_X1 U539 ( .A1(n529), .A2(n555), .ZN(n473) );
  XNOR2_X1 U540 ( .A(n473), .B(KEYINPUT106), .ZN(n485) );
  NAND2_X1 U541 ( .A1(n485), .A2(n474), .ZN(n475) );
  XNOR2_X1 U542 ( .A(n475), .B(KEYINPUT107), .ZN(n480) );
  NAND2_X1 U543 ( .A1(n480), .A2(n487), .ZN(n476) );
  XNOR2_X1 U544 ( .A(n477), .B(n476), .ZN(G1332GAT) );
  NAND2_X1 U545 ( .A1(n541), .A2(n480), .ZN(n478) );
  XNOR2_X1 U546 ( .A(n478), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U547 ( .A1(n551), .A2(n480), .ZN(n479) );
  XNOR2_X1 U548 ( .A(n479), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n482) );
  NAND2_X1 U550 ( .A1(n480), .A2(n494), .ZN(n481) );
  XNOR2_X1 U551 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U552 ( .A(G78GAT), .B(n483), .ZN(G1335GAT) );
  NAND2_X1 U553 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n486), .B(KEYINPUT109), .ZN(n493) );
  NAND2_X1 U555 ( .A1(n493), .A2(n487), .ZN(n488) );
  XNOR2_X1 U556 ( .A(G85GAT), .B(n488), .ZN(G1336GAT) );
  NAND2_X1 U557 ( .A1(n541), .A2(n493), .ZN(n489) );
  XNOR2_X1 U558 ( .A(n489), .B(KEYINPUT110), .ZN(n490) );
  XNOR2_X1 U559 ( .A(G92GAT), .B(n490), .ZN(G1337GAT) );
  XOR2_X1 U560 ( .A(G99GAT), .B(KEYINPUT111), .Z(n492) );
  NAND2_X1 U561 ( .A1(n493), .A2(n551), .ZN(n491) );
  XNOR2_X1 U562 ( .A(n492), .B(n491), .ZN(G1338GAT) );
  NAND2_X1 U563 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U564 ( .A(n495), .B(KEYINPUT44), .ZN(n496) );
  XNOR2_X1 U565 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  NOR2_X1 U566 ( .A1(n569), .A2(n497), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n498), .B(KEYINPUT46), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n578), .B(KEYINPUT112), .ZN(n559) );
  NAND2_X1 U569 ( .A1(n559), .A2(n562), .ZN(n499) );
  XNOR2_X1 U570 ( .A(n501), .B(KEYINPUT47), .ZN(n509) );
  XOR2_X1 U571 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n503) );
  NAND2_X1 U572 ( .A1(n536), .A2(n581), .ZN(n502) );
  XNOR2_X1 U573 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U575 ( .A(KEYINPUT114), .B(n506), .ZN(n507) );
  NAND2_X1 U576 ( .A1(n507), .A2(n569), .ZN(n508) );
  NAND2_X1 U577 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U578 ( .A(KEYINPUT48), .B(n510), .Z(n543) );
  NOR2_X1 U579 ( .A1(n511), .A2(n543), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(KEYINPUT115), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n513), .A2(n528), .ZN(n514) );
  XNOR2_X1 U582 ( .A(KEYINPUT116), .B(n514), .ZN(n516) );
  NAND2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n569), .A2(n523), .ZN(n517) );
  XOR2_X1 U585 ( .A(G113GAT), .B(n517), .Z(G1340GAT) );
  NOR2_X1 U586 ( .A1(n555), .A2(n523), .ZN(n519) );
  XNOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(G1341GAT) );
  NOR2_X1 U589 ( .A1(n559), .A2(n523), .ZN(n521) );
  XNOR2_X1 U590 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(n522), .ZN(G1342GAT) );
  NOR2_X1 U593 ( .A1(n562), .A2(n523), .ZN(n525) );
  XNOR2_X1 U594 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(n526), .ZN(G1343GAT) );
  INV_X1 U597 ( .A(n527), .ZN(n566) );
  NOR2_X1 U598 ( .A1(n566), .A2(n528), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n539), .A2(n529), .ZN(n530) );
  XNOR2_X1 U600 ( .A(G141GAT), .B(n530), .ZN(G1344GAT) );
  INV_X1 U601 ( .A(n539), .ZN(n531) );
  NOR2_X1 U602 ( .A1(n531), .A2(n497), .ZN(n535) );
  XOR2_X1 U603 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n533) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n532) );
  XNOR2_X1 U605 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(G1345GAT) );
  NAND2_X1 U607 ( .A1(n539), .A2(n536), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n537), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U609 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n540), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U611 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n550) );
  XOR2_X1 U612 ( .A(n541), .B(KEYINPUT120), .Z(n542) );
  XNOR2_X1 U613 ( .A(n544), .B(KEYINPUT54), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT64), .ZN(n567) );
  NOR2_X1 U616 ( .A1(n567), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n561) );
  XOR2_X1 U619 ( .A(G169GAT), .B(n553), .Z(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT122), .B(n554), .ZN(G1348GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n561), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n561), .ZN(n560) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT124), .B(n568), .ZN(n582) );
  INV_X1 U633 ( .A(n582), .ZN(n579) );
  NOR2_X1 U634 ( .A1(n579), .A2(n569), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n579), .A2(n471), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n575) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

