//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G104), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT71), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n191), .A2(new_n193), .A3(G214), .A4(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT71), .B(G953), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(G143), .A3(G214), .A4(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT18), .A3(G131), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(KEYINPUT75), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(G146), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT76), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND4_X1   g026(.A1(KEYINPUT76), .A2(new_n203), .A3(new_n205), .A4(new_n211), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT18), .A2(G131), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n197), .A2(new_n199), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n207), .B2(new_n208), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n211), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n220), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n202), .A2(KEYINPUT75), .A3(G140), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n210), .B2(new_n206), .ZN(new_n224));
  OAI211_X1 g038(.A(G146), .B(new_n222), .C1(new_n224), .C2(new_n218), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  AOI211_X1 g042(.A(new_n227), .B(new_n228), .C1(new_n197), .C2(new_n199), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n197), .A2(new_n199), .A3(new_n228), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n200), .A2(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT86), .A4(new_n228), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n227), .A4(new_n235), .ZN(new_n236));
  AOI221_X4 g050(.A(new_n189), .B1(new_n201), .B2(new_n217), .C1(new_n230), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n189), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n219), .A2(new_n211), .A3(new_n220), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n207), .A2(KEYINPUT19), .A3(new_n208), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT19), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n203), .A2(new_n205), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT87), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n210), .A2(new_n244), .A3(new_n241), .ZN(new_n245));
  AND4_X1   g059(.A1(new_n211), .A2(new_n240), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n239), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n233), .A2(new_n235), .A3(new_n234), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n240), .A2(new_n243), .A3(new_n211), .A4(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT88), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n217), .A2(new_n201), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n238), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n187), .B1(new_n237), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(G475), .A2(G902), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n233), .A2(new_n235), .A3(new_n234), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n244), .B1(new_n210), .B2(new_n241), .ZN(new_n258));
  AND4_X1   g072(.A1(new_n244), .A2(new_n203), .A3(new_n205), .A4(new_n241), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(new_n247), .A3(new_n211), .A4(new_n240), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n251), .A3(new_n225), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n253), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n189), .ZN(new_n264));
  INV_X1    g078(.A(new_n236), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n221), .B(new_n225), .C1(new_n234), .C2(new_n227), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n238), .B(new_n253), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(KEYINPUT89), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n256), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT20), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT90), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT90), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n272), .A3(KEYINPUT20), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n237), .A2(new_n254), .ZN(new_n274));
  INV_X1    g088(.A(new_n256), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n274), .A2(KEYINPUT20), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G107), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n280), .A2(G122), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n281), .B2(KEYINPUT14), .ZN(new_n282));
  XNOR2_X1  g096(.A(G116), .B(G122), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G128), .B(G143), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT91), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n284), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n287), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n196), .A2(G128), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT13), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(G128), .B2(new_n196), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  OAI21_X1  g110(.A(G134), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n283), .B(new_n279), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  INV_X1    g115(.A(G217), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n301), .A2(new_n302), .A3(G953), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n300), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  INV_X1    g120(.A(G478), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT15), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n305), .B2(new_n306), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n190), .A2(G952), .ZN(new_n314));
  INV_X1    g128(.A(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n194), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n306), .B(new_n198), .C1(G234), .C2(G237), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT21), .B(G898), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n230), .A2(new_n236), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n238), .B1(new_n322), .B2(new_n253), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n306), .B1(new_n237), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G475), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n278), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT92), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n278), .A2(new_n321), .A3(new_n328), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n280), .B2(G119), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT68), .A3(G116), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n280), .A2(G119), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G113), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT2), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G113), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n340), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n343), .A2(new_n334), .A3(new_n335), .A4(new_n332), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT69), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT69), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(KEYINPUT0), .A2(G128), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n211), .A2(G143), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT64), .B1(new_n196), .B2(G146), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n349), .B(new_n350), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n196), .A2(G146), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(KEYINPUT0), .A2(G128), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n348), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n360));
  INV_X1    g174(.A(G137), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT11), .A3(G134), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n287), .A2(G137), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT11), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n287), .B2(G137), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT65), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT65), .B(new_n365), .C1(new_n287), .C2(G137), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n360), .B(new_n364), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n360), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n369), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n362), .A2(new_n363), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n359), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G128), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT1), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n350), .B(new_n377), .C1(new_n352), .C2(new_n353), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n196), .A2(G146), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT1), .ZN(new_n380));
  OAI21_X1  g194(.A(G128), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n356), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n369), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n361), .A2(G134), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT65), .B1(new_n385), .B2(new_n365), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n373), .B(new_n228), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n363), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G131), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(G131), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT67), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n383), .A2(new_n387), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n347), .A2(new_n375), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n347), .A2(new_n375), .A3(KEYINPUT70), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n342), .A2(new_n344), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AND4_X1   g214(.A1(new_n383), .A2(new_n387), .A3(new_n390), .A4(new_n392), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n354), .A2(new_n358), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n373), .B1(new_n384), .B2(new_n386), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n360), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n372), .A2(new_n373), .A3(new_n371), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT30), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n375), .A2(new_n408), .A3(new_n393), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n400), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n198), .A2(G210), .A3(new_n194), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT27), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT26), .B(G101), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT31), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT31), .ZN(new_n417));
  INV_X1    g231(.A(new_n415), .ZN(new_n418));
  NOR4_X1   g232(.A1(new_n398), .A2(new_n410), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n394), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n399), .B1(new_n401), .B2(new_n406), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n375), .A2(new_n393), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n399), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n396), .A3(new_n397), .A4(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI22_X1  g243(.A1(new_n416), .A2(new_n419), .B1(new_n429), .B2(new_n415), .ZN(new_n430));
  INV_X1    g244(.A(G472), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n306), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n430), .A2(KEYINPUT32), .A3(new_n431), .A4(new_n306), .ZN(new_n435));
  OAI22_X1  g249(.A1(new_n401), .A2(new_n406), .B1(new_n346), .B2(new_n345), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n396), .A2(new_n397), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n421), .B1(new_n437), .B2(KEYINPUT28), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT29), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n418), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n418), .B(new_n421), .C1(new_n427), .C2(new_n428), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n411), .B2(new_n415), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G472), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n434), .A2(new_n435), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT24), .B(G110), .Z(new_n447));
  XNOR2_X1  g261(.A(G119), .B(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT74), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n333), .B2(G128), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n376), .A2(KEYINPUT23), .A3(G119), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n452), .B(new_n453), .C1(G119), .C2(new_n376), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G110), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n226), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  OAI22_X1  g270(.A1(new_n454), .A2(G110), .B1(new_n448), .B2(new_n447), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n225), .B(new_n457), .C1(new_n212), .C2(new_n213), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G137), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT77), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n460), .B(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT78), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n198), .A2(G221), .A3(G234), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n464), .A2(new_n465), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n456), .A3(new_n458), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n302), .B1(G234), .B2(new_n306), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G902), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n476), .B2(new_n306), .ZN(new_n484));
  AOI211_X1 g298(.A(G902), .B(new_n482), .C1(new_n473), .C2(new_n475), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n484), .A2(new_n485), .B1(KEYINPUT79), .B2(KEYINPUT25), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n479), .B1(new_n486), .B2(new_n477), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n446), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n198), .A2(G227), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G140), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n353), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n379), .B1(new_n493), .B2(new_n351), .ZN(new_n494));
  INV_X1    g308(.A(new_n381), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n378), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT80), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n279), .A4(G104), .ZN(new_n500));
  INV_X1    g314(.A(G104), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n501), .A2(KEYINPUT80), .A3(G107), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT3), .B1(new_n501), .B2(G107), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n497), .B(new_n500), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n501), .A2(G107), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n279), .A2(G104), .ZN(new_n506));
  OAI21_X1  g320(.A(G101), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n504), .A2(new_n507), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n504), .A2(KEYINPUT81), .A3(new_n507), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(KEYINPUT10), .A3(new_n383), .A4(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G101), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n520), .A3(G101), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n359), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n511), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n370), .A2(new_n374), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT84), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n511), .A2(new_n516), .A3(new_n524), .A4(new_n522), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n492), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n512), .A2(new_n382), .A3(new_n378), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT82), .B1(new_n509), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT83), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n509), .A2(KEYINPUT83), .A3(new_n533), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n524), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n534), .B2(new_n525), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n492), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n489), .B(new_n306), .C1(new_n532), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n541), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n530), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n531), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n539), .A2(new_n546), .A3(new_n540), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(G469), .C1(new_n547), .C2(new_n492), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n489), .A2(new_n306), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(G110), .B(G122), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n514), .A2(new_n515), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT5), .B1(new_n333), .B2(G116), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n336), .B2(KEYINPUT5), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n344), .B1(new_n558), .B2(new_n337), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n519), .A2(new_n399), .A3(new_n521), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n555), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n554), .C1(new_n556), .C2(new_n559), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n555), .C1(new_n560), .C2(new_n562), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n202), .B1(new_n354), .B2(new_n358), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n378), .A2(new_n382), .A3(new_n202), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G224), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G953), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n571), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n554), .B(KEYINPUT8), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n559), .B(new_n512), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n570), .B1(new_n568), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n578), .B2(new_n570), .ZN(new_n580));
  INV_X1    g394(.A(new_n573), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT7), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n576), .A2(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n569), .A2(KEYINPUT7), .A3(new_n570), .A4(new_n581), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n564), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G210), .B1(G237), .B2(G902), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n575), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n575), .B2(new_n586), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G214), .B1(G237), .B2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n553), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n330), .A2(new_n488), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND2_X1  g409(.A1(new_n427), .A2(new_n428), .ZN(new_n596));
  INV_X1    g410(.A(new_n421), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n375), .A2(new_n408), .A3(new_n393), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n408), .B1(new_n375), .B2(new_n393), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n399), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(new_n415), .A3(new_n396), .A4(new_n397), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n417), .ZN(new_n603));
  INV_X1    g417(.A(new_n398), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT31), .A3(new_n415), .A4(new_n601), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n598), .A2(new_n418), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n606), .B2(G902), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n432), .A3(new_n487), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n608), .A2(new_n553), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n278), .A2(new_n325), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n305), .A2(new_n307), .A3(new_n306), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n305), .B(KEYINPUT33), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n306), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n613), .B2(G478), .ZN(new_n614));
  INV_X1    g428(.A(new_n320), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(new_n591), .C1(new_n588), .C2(new_n589), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n610), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  OR2_X1    g435(.A1(new_n269), .A2(KEYINPUT20), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n271), .A2(new_n273), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n325), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n312), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n623), .A2(new_n617), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NAND2_X1  g444(.A1(new_n607), .A2(new_n432), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n474), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n459), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n486), .A2(new_n477), .B1(new_n478), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n330), .A2(new_n593), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  INV_X1    g452(.A(new_n553), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n592), .A2(new_n634), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n446), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n317), .B1(new_n318), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n623), .A2(new_n625), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  INV_X1    g461(.A(new_n602), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n437), .A2(new_n418), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n306), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G472), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n434), .A2(new_n435), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT93), .B(KEYINPUT38), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n590), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n313), .A2(new_n591), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n278), .B2(new_n325), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n634), .A2(new_n652), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n643), .B(KEYINPUT39), .Z(new_n658));
  NAND3_X1  g472(.A1(new_n551), .A2(new_n552), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT94), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n551), .A2(KEYINPUT94), .A3(new_n552), .A4(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n665), .A3(new_n662), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n657), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n610), .A2(new_n669), .A3(new_n614), .A4(new_n644), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n269), .A2(new_n272), .A3(KEYINPUT20), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n272), .B1(new_n269), .B2(KEYINPUT20), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n671), .A2(new_n672), .A3(new_n276), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n614), .B(new_n644), .C1(new_n673), .C2(new_n624), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT95), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n641), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n610), .A2(new_n614), .A3(new_n617), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n532), .A2(new_n542), .ZN(new_n680));
  OAI21_X1  g494(.A(G469), .B1(new_n680), .B2(G902), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n681), .A2(new_n552), .A3(new_n543), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n488), .A2(new_n678), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n446), .A2(new_n487), .A3(new_n682), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT96), .B1(new_n684), .B2(new_n618), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT97), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n626), .A2(new_n446), .A3(new_n487), .A4(new_n682), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  NAND3_X1  g505(.A1(new_n446), .A2(new_n640), .A3(new_n682), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n329), .B2(new_n327), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n333), .ZN(G21));
  NAND2_X1  g508(.A1(new_n437), .A2(KEYINPUT28), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n597), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n603), .A2(new_n605), .B1(new_n696), .B2(new_n418), .ZN(new_n697));
  NOR2_X1   g511(.A1(G472), .A2(G902), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT98), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n416), .A2(new_n419), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n438), .A2(new_n415), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n701), .B(new_n698), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n487), .A2(new_n607), .A3(new_n700), .A4(new_n704), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n615), .A2(new_n681), .A3(new_n552), .A4(new_n543), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n590), .A3(new_n656), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT99), .B(G122), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G24));
  NAND3_X1  g523(.A1(new_n682), .A2(new_n591), .A3(new_n590), .ZN(new_n710));
  INV_X1    g524(.A(new_n634), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n607), .A3(new_n700), .A4(new_n704), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n670), .A3(new_n675), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n675), .A2(new_n670), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n588), .A2(new_n589), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n552), .A3(new_n591), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n548), .B(KEYINPUT100), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n543), .A2(new_n550), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n446), .A3(new_n487), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n716), .B1(new_n717), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n487), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n435), .A2(new_n445), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n434), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n432), .A2(KEYINPUT101), .A3(new_n433), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n719), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n548), .B(KEYINPUT100), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n721), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n716), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n670), .A3(new_n735), .A4(new_n675), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n725), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NAND4_X1  g552(.A1(new_n723), .A2(new_n446), .A3(new_n487), .A4(new_n645), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NOR2_X1   g554(.A1(new_n547), .A2(new_n492), .ZN(new_n741));
  INV_X1    g555(.A(new_n545), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT45), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n545), .B(new_n744), .C1(new_n547), .C2(new_n492), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n550), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(G469), .C1(new_n746), .C2(G902), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n543), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n552), .A3(new_n658), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n718), .A2(new_n591), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n631), .A2(new_n711), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n278), .A2(new_n614), .A3(new_n325), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT43), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(KEYINPUT102), .A3(new_n759), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n755), .B1(new_n764), .B2(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(KEYINPUT44), .B2(new_n764), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OR3_X1    g581(.A1(new_n446), .A2(new_n487), .A3(new_n753), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n751), .A2(new_n552), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n552), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n717), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NAND2_X1  g590(.A1(new_n707), .A2(new_n690), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n693), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n312), .A2(new_n325), .A3(new_n644), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n634), .A2(new_n753), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n446), .A2(new_n780), .A3(new_n639), .A4(new_n623), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n739), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n737), .A2(new_n686), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n734), .A2(new_n712), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n675), .A3(new_n670), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT104), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n675), .A3(new_n787), .A4(new_n670), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n610), .A2(new_n614), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n610), .B2(new_n312), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n608), .A2(new_n553), .A3(new_n616), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n594), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n636), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT105), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n594), .A2(new_n636), .A3(new_n793), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n788), .B2(new_n786), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n778), .A2(new_n686), .A3(new_n782), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT105), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n737), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n656), .A2(new_n590), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n720), .A2(new_n722), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n634), .A2(new_n552), .A3(new_n644), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n652), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n714), .A2(new_n676), .A3(new_n805), .A4(new_n646), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n796), .A2(new_n801), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n796), .A2(new_n801), .A3(new_n808), .A4(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT54), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n783), .A2(new_n795), .A3(new_n810), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n809), .A2(new_n810), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n760), .A2(new_n316), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n681), .A2(new_n543), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n732), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n822), .A2(new_n726), .A3(new_n316), .ZN(new_n825));
  INV_X1    g639(.A(new_n652), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n610), .A2(new_n614), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n824), .A2(new_n712), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n820), .A2(new_n705), .ZN(new_n830));
  INV_X1    g644(.A(new_n682), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n654), .A3(new_n591), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n820), .A2(new_n705), .ZN(new_n835));
  INV_X1    g649(.A(new_n832), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n829), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n821), .B(KEYINPUT106), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n771), .B(new_n772), .C1(new_n552), .C2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n830), .A2(new_n840), .A3(new_n754), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT51), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n731), .A3(new_n823), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(KEYINPUT109), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT48), .B1(new_n843), .B2(KEYINPUT109), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  OAI221_X1 g662(.A(new_n314), .B1(new_n790), .B2(new_n827), .C1(new_n835), .C2(new_n710), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n842), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT108), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n838), .A2(KEYINPUT107), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n841), .A2(KEYINPUT51), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n838), .B2(KEYINPUT107), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n851), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n838), .A2(KEYINPUT107), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT108), .A3(new_n852), .A4(new_n854), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n819), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n487), .A2(new_n552), .A3(new_n591), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT103), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n821), .B(KEYINPUT49), .Z(new_n864));
  OR4_X1    g678(.A1(new_n652), .A2(new_n863), .A3(new_n654), .A4(new_n864), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n860), .A2(new_n861), .B1(new_n757), .B2(new_n865), .ZN(G75));
  NOR2_X1   g680(.A1(new_n198), .A2(G952), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(G210), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n816), .A2(new_n869), .A3(new_n306), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n565), .A2(new_n567), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n574), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT112), .B(KEYINPUT56), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n868), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n815), .A2(new_n808), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n306), .B1(new_n811), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT111), .B1(new_n880), .B2(new_n874), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT111), .ZN(new_n882));
  INV_X1    g696(.A(new_n874), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n882), .B(new_n883), .C1(new_n870), .C2(KEYINPUT56), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n877), .B1(new_n881), .B2(new_n884), .ZN(G51));
  XNOR2_X1  g699(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n549), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n811), .A2(new_n817), .A3(new_n878), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n817), .B1(new_n811), .B2(new_n878), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n680), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n879), .A2(G469), .A3(new_n746), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n867), .B1(new_n892), .B2(new_n893), .ZN(G54));
  NAND2_X1  g708(.A1(new_n811), .A2(new_n878), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n255), .A2(new_n268), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n895), .A2(G902), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n868), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n897), .B1(new_n879), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT114), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n895), .A2(G902), .A3(new_n898), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n896), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n868), .A4(new_n899), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n906), .ZN(G60));
  NOR2_X1   g721(.A1(new_n888), .A2(new_n889), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n612), .B(KEYINPUT115), .ZN(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n910));
  NAND2_X1  g724(.A1(G478), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n868), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n909), .B1(new_n819), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n895), .A2(new_n633), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n918), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n475), .B(new_n473), .C1(new_n816), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n922), .A3(new_n868), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n920), .A2(new_n922), .A3(KEYINPUT61), .A4(new_n868), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G66));
  OAI21_X1  g741(.A(G953), .B1(new_n319), .B2(new_n572), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT117), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n778), .A2(new_n686), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n797), .ZN(new_n931));
  INV_X1    g745(.A(new_n198), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n871), .B1(G898), .B2(new_n198), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  NOR2_X1   g749(.A1(new_n599), .A2(new_n600), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n260), .A2(new_n240), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n936), .B(new_n937), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n659), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n488), .A2(new_n791), .A3(new_n940), .A4(new_n754), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n773), .B2(new_n774), .ZN(new_n942));
  INV_X1    g756(.A(new_n755), .ZN(new_n943));
  INV_X1    g757(.A(new_n756), .ZN(new_n944));
  INV_X1    g758(.A(new_n763), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT102), .B1(new_n758), .B2(new_n759), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT44), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n764), .A2(KEYINPUT44), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n667), .A2(new_n676), .A3(new_n646), .A4(new_n714), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT118), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n952), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n766), .A2(new_n956), .A3(new_n957), .A4(new_n942), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n939), .B1(new_n959), .B2(new_n198), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT119), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n198), .B1(G227), .B2(G900), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT120), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n737), .A2(new_n739), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT121), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n714), .A2(new_n646), .A3(new_n676), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n752), .A2(new_n802), .A3(new_n731), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n775), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n766), .A3(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(new_n932), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n938), .B1(G900), .B2(new_n932), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n960), .A2(KEYINPUT119), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n961), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n970), .A2(new_n971), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n962), .B1(new_n975), .B2(new_n960), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G72));
  NOR2_X1   g791(.A1(new_n411), .A2(new_n418), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n954), .A2(new_n958), .A3(new_n931), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT122), .B(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT123), .Z(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n931), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n984), .B1(new_n969), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n411), .A2(new_n418), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT125), .Z(new_n991));
  AOI21_X1  g805(.A(new_n867), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n411), .B(new_n415), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n983), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n813), .A2(KEYINPUT126), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT126), .B1(new_n813), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n987), .A2(new_n997), .ZN(G57));
endmodule


