//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n538, new_n539, new_n540, new_n541, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(G220));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G137), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n460), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n475), .B2(G2105), .ZN(G160));
  NAND2_X1  g051(.A1(new_n467), .A2(new_n469), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n461), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n460), .A2(new_n493), .A3(G138), .A4(new_n461), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT71), .A3(G543), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(new_n500), .B1(KEYINPUT5), .B2(new_n497), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OR3_X1    g078(.A1(new_n502), .A2(KEYINPUT72), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT72), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(G88), .B1(new_n509), .B2(G50), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  NAND2_X1  g087(.A1(new_n507), .A2(G89), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT7), .Z(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(G51), .B2(new_n509), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G168));
  AOI22_X1  g094(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n503), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n501), .A2(new_n506), .ZN(new_n522));
  INV_X1    g097(.A(G90), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT73), .B(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n522), .A2(new_n523), .B1(new_n508), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(G171));
  AOI22_X1  g101(.A1(new_n507), .A2(G81), .B1(new_n509), .B2(G43), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT75), .Z(G153));
  AND3_X1   g110(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G36), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT76), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT8), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT77), .Z(G188));
  NAND2_X1  g117(.A1(G78), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(new_n501), .ZN(new_n544));
  INV_X1    g119(.A(G65), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  OR3_X1    g123(.A1(new_n508), .A2(KEYINPUT9), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT9), .B1(new_n508), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n507), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n522), .A2(KEYINPUT78), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n561));
  NAND2_X1  g136(.A1(G168), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(G286));
  NAND2_X1  g139(.A1(new_n555), .A2(new_n556), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G87), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n501), .A2(G74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(G49), .B2(new_n509), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n565), .A2(G86), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n565), .A2(KEYINPUT80), .A3(G86), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n503), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(G48), .B2(new_n509), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n503), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n522), .A2(new_n580), .B1(new_n508), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n579), .A2(new_n582), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G171), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n544), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n565), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT81), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(KEYINPUT81), .B2(new_n585), .ZN(G284));
  OAI21_X1  g174(.A(new_n598), .B1(KEYINPUT81), .B2(new_n585), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n558), .B2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(KEYINPUT82), .B2(new_n601), .ZN(G297));
  XNOR2_X1  g180(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n532), .A2(new_n584), .ZN(new_n609));
  INV_X1    g184(.A(new_n595), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT10), .B1(new_n565), .B2(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n590), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n609), .B1(new_n613), .B2(new_n584), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n460), .A2(new_n464), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n478), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n480), .A2(G135), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n622), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n618), .A2(G2100), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n619), .A2(new_n625), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT85), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT84), .B(G2438), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT16), .B(G1341), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n635), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(KEYINPUT17), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n654), .C1(new_n655), .C2(new_n651), .ZN(new_n656));
  OR3_X1    g231(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n650), .ZN(new_n657));
  OAI21_X1  g232(.A(KEYINPUT18), .B1(new_n654), .B2(new_n650), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2096), .B(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n668), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1991), .ZN(new_n675));
  INV_X1    g250(.A(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n683), .B1(new_n680), .B2(new_n681), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G6), .ZN(new_n689));
  INV_X1    g264(.A(G305), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(G288), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(G166), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G22), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT89), .B(G1971), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n698), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n693), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT34), .ZN(new_n706));
  MUX2_X1   g281(.A(G24), .B(G290), .S(G16), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1986), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n478), .A2(G119), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n480), .A2(G131), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n461), .A2(G107), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT87), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n708), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n706), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT36), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT36), .ZN(new_n725));
  AOI22_X1  g300(.A1(G128), .A2(new_n478), .B1(new_n480), .B2(G140), .ZN(new_n726));
  NOR3_X1   g301(.A1(KEYINPUT91), .A2(G104), .A3(G2105), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT91), .B1(G104), .B2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n715), .A2(G26), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT92), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2067), .ZN(new_n737));
  OR2_X1    g312(.A1(G29), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n464), .A2(G103), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT25), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G139), .B2(new_n480), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n461), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n715), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n478), .A2(G129), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n480), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n464), .A2(G105), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  NAND4_X1  g326(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G32), .B(new_n752), .S(G29), .Z(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n624), .A2(new_n715), .ZN(new_n756));
  INV_X1    g331(.A(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND4_X1   g337(.A1(new_n746), .A2(new_n755), .A3(new_n756), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G27), .A2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n737), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G21), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G168), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT98), .B(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n688), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n596), .B2(new_n688), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT90), .B(G1348), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n768), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n688), .A2(G20), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT23), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT23), .B1(new_n558), .B2(new_n688), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n779), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT101), .B(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n776), .B2(new_n775), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n715), .A2(G35), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT99), .Z(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n715), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G1961), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(G1961), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n793), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n688), .A2(G19), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n533), .B2(new_n688), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1341), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n744), .A2(new_n745), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT94), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n805));
  INV_X1    g380(.A(G34), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n715), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT96), .Z(new_n809));
  INV_X1    g384(.A(G160), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n715), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G2084), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n799), .A2(new_n802), .A3(new_n804), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n778), .A2(new_n786), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n724), .A2(new_n725), .B1(new_n816), .B2(new_n817), .ZN(G311));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n816), .ZN(new_n819));
  INV_X1    g394(.A(new_n725), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n723), .A2(KEYINPUT36), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G150));
  AOI22_X1  g397(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n503), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n522), .A2(new_n825), .B1(new_n508), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n596), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n533), .A2(new_n829), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n532), .A2(new_n828), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n833), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT104), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n838), .A2(new_n839), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT103), .B1(new_n837), .B2(KEYINPUT39), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(KEYINPUT104), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n831), .B1(new_n843), .B2(new_n847), .ZN(G145));
  NAND2_X1  g423(.A1(new_n492), .A2(new_n494), .ZN(new_n849));
  INV_X1    g424(.A(new_n490), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n752), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n730), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n478), .A2(G130), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n480), .A2(G142), .ZN(new_n860));
  OR2_X1    g435(.A1(G106), .A2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n617), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n713), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT107), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n858), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(G160), .B(KEYINPUT105), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n484), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n624), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n858), .B2(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n856), .A2(new_n857), .A3(new_n865), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n874), .A2(KEYINPUT108), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(KEYINPUT108), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g453(.A(G288), .B(G290), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(G303), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n690), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT111), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n880), .B(G305), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n596), .A2(G299), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT109), .B1(new_n612), .B2(new_n558), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT109), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n596), .A2(new_n890), .A3(G299), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n596), .B2(G299), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n612), .A2(KEYINPUT110), .A3(new_n558), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n889), .A2(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n894), .B1(KEYINPUT41), .B2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n613), .B(new_n836), .Z(new_n900));
  MUX2_X1   g475(.A(new_n893), .B(new_n899), .S(new_n900), .Z(new_n901));
  AND2_X1   g476(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n887), .A2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n828), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n828), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n892), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G301), .B1(new_n562), .B2(new_n563), .ZN(new_n910));
  NOR2_X1   g485(.A1(G171), .A2(new_n518), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n836), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n834), .B(new_n835), .C1(new_n910), .C2(new_n911), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n909), .B(new_n915), .C1(new_n898), .C2(new_n908), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n915), .B2(new_n892), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n914), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n893), .A2(KEYINPUT112), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n881), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n899), .A2(new_n915), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n915), .A2(new_n892), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n884), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n907), .B1(new_n928), .B2(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n924), .B1(new_n899), .B2(new_n915), .ZN(new_n930));
  AOI21_X1  g505(.A(G37), .B1(new_n930), .B2(new_n884), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n889), .A2(new_n891), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n896), .A2(new_n897), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n908), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n919), .B1(new_n936), .B2(new_n894), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n881), .B1(new_n937), .B2(new_n924), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n931), .A2(KEYINPUT113), .A3(new_n932), .A4(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n926), .A2(new_n938), .A3(new_n932), .A4(new_n927), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT113), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n929), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n931), .A2(new_n932), .A3(new_n922), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n932), .B1(new_n931), .B2(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n907), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(G397));
  INV_X1    g522(.A(KEYINPUT114), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(G160), .B2(G40), .ZN(new_n949));
  INV_X1    g524(.A(new_n474), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n470), .B2(KEYINPUT70), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n461), .B1(new_n951), .B2(new_n473), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  NOR4_X1   g528(.A1(new_n952), .A2(KEYINPUT114), .A3(new_n953), .A4(new_n466), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G164), .B2(G1384), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(KEYINPUT115), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(KEYINPUT115), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n730), .B(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n752), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(KEYINPUT46), .A3(new_n676), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n961), .B2(G1996), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n752), .B(G1996), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n713), .A2(new_n720), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(G2067), .B2(new_n730), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n962), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n962), .A2(KEYINPUT48), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n980));
  INV_X1    g555(.A(new_n978), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n961), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n713), .B(new_n720), .Z(new_n983));
  NAND2_X1  g558(.A1(new_n973), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n979), .B(new_n982), .C1(new_n961), .C2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n971), .A2(new_n977), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G303), .A2(G8), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT55), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1971), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n851), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n957), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n955), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G164), .B2(G1384), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n851), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n949), .B2(new_n954), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n995), .B1(G2090), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n990), .A2(G8), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G164), .A2(G1384), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n475), .A2(G2105), .ZN(new_n1006));
  INV_X1    g581(.A(new_n466), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(G40), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT114), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G160), .A2(new_n948), .A3(G40), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1005), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n572), .A2(new_n1014), .A3(new_n573), .A4(new_n576), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n1016));
  INV_X1    g591(.A(G86), .ZN(new_n1017));
  INV_X1    g592(.A(G48), .ZN(new_n1018));
  OAI22_X1  g593(.A1(new_n522), .A2(new_n1017), .B1(new_n508), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(G1981), .B1(new_n575), .B2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1016), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1013), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1013), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1013), .B(new_n1028), .C1(new_n1025), .C2(G288), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1003), .A2(new_n1023), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n998), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n949), .A2(new_n954), .B1(new_n1004), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g609(.A(KEYINPUT118), .B1(new_n1004), .B2(new_n1031), .C1(new_n949), .C2(new_n954), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1004), .A2(new_n996), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n995), .B1(new_n1037), .B2(G2090), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n990), .B1(new_n1038), .B2(G8), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1000), .B(new_n812), .C1(new_n949), .C2(new_n954), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT119), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n772), .B1(new_n955), .B2(new_n994), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n812), .A4(new_n1000), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1047), .A2(G286), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1030), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1023), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1002), .A2(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n989), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(KEYINPUT63), .A3(new_n1003), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1049), .A2(KEYINPUT63), .B1(new_n1053), .B2(new_n1048), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n695), .A2(new_n1025), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT117), .ZN(new_n1056));
  OR3_X1    g631(.A1(new_n1056), .A2(new_n1022), .A3(new_n1021), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1024), .B1(new_n1057), .B2(new_n1015), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1003), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1050), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  INV_X1    g637(.A(new_n557), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n546), .A2(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n552), .A2(new_n557), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1037), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n994), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT120), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1043), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1068), .B(new_n1075), .C1(new_n1037), .C2(new_n1070), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1062), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1032), .A2(new_n1033), .B1(new_n996), .B2(new_n1004), .ZN(new_n1080));
  AOI21_X1  g655(.A(G1956), .B1(new_n1080), .B2(new_n1035), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1068), .B1(new_n1081), .B2(new_n1075), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1071), .A2(new_n1069), .A3(new_n1076), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT61), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(G1341), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT122), .B1(new_n1011), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1004), .B1(new_n949), .B2(new_n954), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1086), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1043), .A2(new_n1072), .A3(new_n676), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n533), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT59), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(new_n533), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n776), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n963), .A2(new_n1011), .B1(new_n1001), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n612), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1089), .A2(G2067), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n776), .B1(new_n1043), .B2(new_n1000), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n596), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1105), .A2(KEYINPUT60), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1079), .A2(new_n1084), .A3(new_n1098), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1104), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1083), .B1(new_n1077), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1043), .A2(new_n1072), .A3(new_n766), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n1001), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT53), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n955), .A2(new_n994), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT125), .B1(new_n1118), .B2(new_n766), .ZN(new_n1119));
  OAI211_X1 g694(.A(G301), .B(new_n1115), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT127), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(KEYINPUT125), .A3(new_n766), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT53), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(G301), .A4(new_n1115), .ZN(new_n1126));
  OR4_X1    g701(.A1(new_n1113), .A2(new_n994), .A3(G2078), .A4(new_n1008), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1115), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1121), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT54), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1115), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G171), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1128), .A2(G171), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT54), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1132), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1131), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1111), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1047), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1046), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G168), .A2(new_n1012), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(KEYINPUT51), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1144), .A2(KEYINPUT124), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1047), .B1(new_n1012), .B2(G168), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT51), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1046), .A2(new_n1146), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1142), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1141), .A2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1030), .A2(new_n1039), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1148), .A2(new_n1149), .B1(KEYINPUT51), .B2(new_n1152), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1159), .A2(new_n1151), .B1(new_n1146), .B2(new_n1046), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT62), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1158), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1061), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(G290), .B(G1986), .Z(new_n1165));
  AOI21_X1  g740(.A(new_n961), .B1(new_n985), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n987), .B1(new_n1164), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g742(.A(G319), .B(new_n661), .C1(new_n642), .C2(new_n643), .ZN(new_n1169));
  NOR3_X1   g743(.A1(new_n685), .A2(new_n686), .A3(new_n1169), .ZN(new_n1170));
  OAI211_X1 g744(.A(new_n1170), .B(new_n877), .C1(new_n944), .C2(new_n945), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


