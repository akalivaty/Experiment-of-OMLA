//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT4), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G104), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT3), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n190), .B(G101), .C1(new_n198), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G116), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT2), .B(G113), .Z(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n206), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT2), .B(G113), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n209), .A2(KEYINPUT66), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT66), .B1(new_n209), .B2(new_n212), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n202), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT79), .B(G101), .C1(new_n198), .C2(new_n201), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT78), .B(G107), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n196), .B1(new_n218), .B2(G104), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n200), .C1(new_n219), .C2(KEYINPUT3), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n198), .B2(new_n201), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n215), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n218), .A2(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n199), .A2(G107), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n229), .B(G113), .C1(new_n230), .C2(new_n210), .ZN(new_n231));
  AND4_X1   g045(.A1(new_n209), .A2(new_n220), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n189), .B1(new_n225), .B2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n216), .A4(new_n220), .ZN(new_n234));
  INV_X1    g048(.A(new_n215), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n232), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n188), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n238), .A3(KEYINPUT6), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n240));
  OR3_X1    g054(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n188), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n244), .A2(new_n246), .A3(KEYINPUT0), .A4(G128), .ZN(new_n247));
  XNOR2_X1  g061(.A(G143), .B(G146), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n242), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(KEYINPUT80), .A3(G125), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n245), .A2(G146), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n243), .A2(G143), .ZN(new_n257));
  OAI211_X1 g071(.A(G128), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n244), .B(new_n246), .C1(KEYINPUT1), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n252), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(new_n254), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G224), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n239), .A2(new_n241), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT7), .B1(new_n264), .B2(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n253), .A2(new_n254), .A3(new_n262), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n240), .B2(new_n188), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n188), .B(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n220), .A2(new_n228), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n231), .A2(new_n209), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G210), .B1(G237), .B2(G902), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n267), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n283), .B(KEYINPUT82), .Z(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n267), .B2(new_n282), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT83), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n267), .A2(new_n282), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n285), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n267), .A2(new_n282), .A3(new_n283), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n187), .ZN(new_n295));
  INV_X1    g109(.A(G953), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(G952), .ZN(new_n297));
  NAND2_X1  g111(.A1(G234), .A2(G237), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT21), .B(G898), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(G902), .A3(G953), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n289), .A2(new_n295), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G137), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n296), .A2(G221), .A3(G234), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT71), .A2(G125), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G140), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT72), .B1(new_n312), .B2(G125), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT71), .A3(G125), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT16), .B1(new_n312), .B2(G125), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT73), .A2(G146), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(KEYINPUT73), .A2(G146), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT70), .B1(new_n259), .B2(G119), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n203), .A3(G128), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n259), .A2(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT24), .B(G110), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n203), .A2(G128), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n332), .B1(G110), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n317), .B1(new_n315), .B2(KEYINPUT16), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT73), .A3(G146), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n324), .A2(new_n325), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n319), .A2(G146), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n312), .A2(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n252), .A2(G140), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n343), .A2(new_n344), .A3(new_n243), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n330), .A2(new_n331), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT75), .B(G110), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT76), .B1(new_n342), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n341), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n324), .A2(new_n340), .A3(new_n338), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n308), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G902), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n342), .A2(new_n349), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n341), .A4(new_n307), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n355), .A2(new_n356), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n363), .A4(new_n356), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G217), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(G234), .B2(new_n356), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n355), .A2(new_n363), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n372), .A2(G902), .A3(new_n370), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(KEYINPUT77), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n376));
  INV_X1    g190(.A(new_n370), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n366), .B2(new_n367), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n378), .B2(new_n373), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G137), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT11), .A3(G134), .ZN(new_n382));
  INV_X1    g196(.A(G134), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G137), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT64), .ZN(new_n386));
  INV_X1    g200(.A(G131), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT11), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n383), .B2(G137), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n382), .A3(new_n387), .A4(new_n384), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT64), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n383), .A2(G137), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n381), .A2(G134), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n258), .A2(new_n396), .A3(new_n260), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(new_n382), .A3(new_n384), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n390), .A2(new_n392), .B1(G131), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n402), .A3(new_n250), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(G131), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n391), .A2(KEYINPUT64), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n391), .A2(KEYINPUT64), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT65), .B1(new_n407), .B2(new_n251), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n399), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n399), .B(KEYINPUT30), .C1(new_n401), .C2(new_n250), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT67), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n407), .A2(new_n251), .B1(new_n393), .B2(new_n398), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT30), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n213), .A2(new_n214), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT31), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT26), .B(G101), .Z(new_n422));
  NOR2_X1   g236(.A1(G237), .A2(G953), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G210), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n422), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n418), .B2(new_n414), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n420), .A2(new_n421), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n421), .B1(new_n420), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n414), .A2(new_n418), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT28), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n397), .B1(new_n390), .B2(new_n392), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n402), .B1(new_n401), .B2(new_n250), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n407), .A2(KEYINPUT65), .A3(new_n251), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n418), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n427), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n430), .A2(new_n431), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(G472), .A2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT32), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n415), .B1(new_n414), .B2(KEYINPUT30), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n250), .B1(new_n393), .B2(new_n404), .ZN(new_n446));
  NOR4_X1   g260(.A1(new_n446), .A2(new_n434), .A3(KEYINPUT67), .A4(new_n410), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n445), .A2(new_n447), .B1(new_n437), .B2(KEYINPUT30), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n429), .B1(new_n448), .B2(new_n418), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT31), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT28), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n432), .B(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n428), .B1(new_n452), .B2(new_n438), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n420), .A2(new_n421), .A3(new_n429), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT32), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n442), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n444), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n420), .A2(new_n428), .A3(new_n432), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n427), .B1(new_n452), .B2(new_n438), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT29), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n432), .A2(new_n451), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n419), .B1(new_n434), .B2(new_n446), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n432), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT28), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n427), .A2(KEYINPUT29), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n356), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G472), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n380), .B1(new_n458), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G237), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n296), .A3(G214), .ZN(new_n474));
  NOR2_X1   g288(.A1(KEYINPUT84), .A2(G143), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n423), .B(G214), .C1(KEYINPUT84), .C2(G143), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT17), .A3(G131), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n478), .A2(KEYINPUT87), .A3(KEYINPUT17), .A4(G131), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n324), .A2(new_n340), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(G131), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n476), .A2(new_n477), .A3(new_n387), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n484), .A2(KEYINPUT88), .A3(new_n485), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G113), .B(G122), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(G104), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n345), .B1(G146), .B2(new_n315), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT18), .A2(G131), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n478), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n492), .A2(new_n495), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n495), .B1(new_n492), .B2(new_n502), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n356), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G475), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n315), .A2(KEYINPUT19), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT19), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n343), .A2(new_n344), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n243), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n511), .B(KEYINPUT86), .C1(new_n243), .C2(new_n339), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n484), .A2(new_n486), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT86), .B1(new_n342), .B2(new_n511), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n502), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n494), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n492), .A2(new_n495), .A3(new_n502), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n507), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  AOI211_X1 g336(.A(KEYINPUT20), .B(new_n522), .C1(new_n517), .C2(new_n518), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n506), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT89), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n506), .B(new_n526), .C1(new_n521), .C2(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G221), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT9), .B(G234), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n532), .B2(new_n356), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n202), .A2(new_n251), .ZN(new_n535));
  INV_X1    g349(.A(new_n224), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n261), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n220), .A2(new_n539), .A3(new_n228), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT10), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT10), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n220), .A2(new_n539), .A3(new_n542), .A4(new_n228), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n544), .A3(new_n401), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n276), .A2(new_n261), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n540), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT12), .B1(new_n547), .B2(new_n407), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n549));
  AOI211_X1 g363(.A(new_n549), .B(new_n401), .C1(new_n546), .C2(new_n540), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G110), .B(G140), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n296), .A2(G227), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n552), .B(new_n553), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n234), .A2(new_n535), .B1(new_n541), .B2(new_n543), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n556), .B2(new_n401), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n401), .B1(new_n538), .B2(new_n544), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(G469), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(G469), .A2(G902), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n538), .A2(new_n544), .A3(new_n401), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n554), .B1(new_n564), .B2(new_n558), .ZN(new_n565));
  INV_X1    g379(.A(new_n554), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n545), .B(new_n566), .C1(new_n548), .C2(new_n550), .ZN(new_n567));
  AOI211_X1 g381(.A(G469), .B(G902), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n534), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  XNOR2_X1  g385(.A(G116), .B(G122), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n218), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n245), .A2(G128), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n259), .A2(G143), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G134), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n383), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n205), .A2(KEYINPUT14), .A3(G122), .ZN(new_n582));
  XOR2_X1   g396(.A(G116), .B(G122), .Z(new_n583));
  OAI211_X1 g397(.A(G107), .B(new_n582), .C1(new_n583), .C2(KEYINPUT14), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n218), .A2(new_n572), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT90), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n575), .A2(new_n581), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n259), .B2(G143), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n577), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n576), .A2(new_n588), .ZN(new_n591));
  OAI21_X1  g405(.A(G134), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n218), .A2(new_n572), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n592), .B(new_n580), .C1(new_n573), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n531), .A2(new_n369), .A3(G953), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n595), .B(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT91), .B1(new_n598), .B2(new_n356), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n595), .A2(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n587), .B2(new_n594), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT91), .B(new_n356), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n571), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n356), .B1(new_n600), .B2(new_n601), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n571), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n529), .A2(new_n569), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n304), .A2(new_n472), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  AOI22_X1  g427(.A1(new_n551), .A2(new_n554), .B1(new_n557), .B2(new_n559), .ZN(new_n614));
  OAI21_X1  g428(.A(G469), .B1(new_n614), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n565), .A2(new_n567), .ZN(new_n616));
  INV_X1    g430(.A(G469), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n356), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n533), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n455), .A2(new_n442), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT77), .B1(new_n371), .B2(new_n374), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n378), .A2(new_n376), .A3(new_n373), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n441), .B2(G902), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n621), .A2(new_n624), .A3(KEYINPUT92), .A4(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n620), .A3(new_n619), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n380), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n605), .A2(new_n570), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT95), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n356), .A2(G478), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n525), .A2(new_n527), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n283), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n290), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT93), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n292), .ZN(new_n641));
  INV_X1    g455(.A(new_n187), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n283), .B1(new_n267), .B2(new_n282), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(KEYINPUT93), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n637), .A2(new_n303), .A3(new_n641), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n630), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT34), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  OAI211_X1 g462(.A(new_n610), .B(new_n506), .C1(new_n521), .C2(new_n523), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n303), .A2(new_n641), .A3(new_n650), .A4(new_n644), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n626), .A2(new_n629), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n370), .A2(G902), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n352), .A2(new_n354), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n308), .A2(KEYINPUT36), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n656), .B(new_n657), .Z(new_n658));
  AOI21_X1  g472(.A(new_n378), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n625), .A2(new_n620), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n304), .A2(new_n611), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  XOR2_X1   g478(.A(new_n299), .B(KEYINPUT96), .Z(new_n665));
  NOR2_X1   g479(.A1(new_n302), .A2(G900), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT98), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n659), .B1(new_n458), .B2(new_n471), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n290), .A2(KEYINPUT93), .A3(new_n638), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n292), .A2(new_n640), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n187), .B(new_n672), .C1(new_n673), .C2(new_n643), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n670), .A2(new_n671), .A3(new_n619), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT99), .B(G128), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G30));
  XOR2_X1   g492(.A(new_n668), .B(KEYINPUT39), .Z(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n569), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n420), .A2(new_n432), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n427), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n465), .A2(new_n432), .A3(new_n428), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(KEYINPUT101), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n356), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT101), .B1(new_n684), .B2(new_n685), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n458), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n293), .B(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n525), .A2(new_n527), .A3(new_n610), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n660), .A2(new_n693), .A3(new_n642), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n682), .A2(new_n690), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  INV_X1    g510(.A(new_n668), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n525), .A2(new_n527), .A3(new_n636), .A4(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n671), .A2(new_n619), .A3(new_n675), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n455), .A2(new_n456), .A3(new_n442), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n456), .B1(new_n455), .B2(new_n442), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n471), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n616), .A2(new_n356), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n534), .A3(new_n618), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n624), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n702), .B1(new_n710), .B2(new_n645), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n525), .A2(new_n527), .A3(new_n636), .ZN(new_n712));
  INV_X1    g526(.A(new_n303), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n674), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n472), .A2(new_n714), .A3(KEYINPUT102), .A4(new_n709), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n651), .A2(new_n705), .A3(new_n624), .A4(new_n709), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR2_X1   g534(.A1(new_n674), .A2(new_n708), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n713), .B(new_n610), .C1(new_n525), .C2(new_n527), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n705), .A3(new_n660), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NOR2_X1   g538(.A1(new_n674), .A2(new_n713), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n693), .A2(new_n708), .ZN(new_n726));
  INV_X1    g540(.A(G472), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n455), .B2(new_n356), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n430), .A2(new_n431), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n468), .A2(new_n428), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n443), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n371), .A2(KEYINPUT103), .A3(new_n374), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n378), .B2(new_n373), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n725), .A2(new_n726), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n659), .A2(new_n728), .A3(new_n731), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(new_n721), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NAND3_X1  g558(.A1(new_n291), .A2(new_n187), .A3(new_n292), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n569), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n472), .A2(new_n740), .A3(new_n741), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n284), .A2(new_n287), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n619), .A2(new_n750), .A3(KEYINPUT42), .A4(new_n187), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n749), .A2(new_n739), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n705), .ZN(new_n753));
  INV_X1    g567(.A(new_n736), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n747), .A2(new_n748), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n387), .ZN(G33));
  NAND3_X1  g571(.A1(new_n670), .A2(new_n472), .A3(new_n746), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(new_n745), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n528), .A2(new_n636), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n659), .B1(new_n625), .B2(new_n620), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT107), .B(new_n760), .C1(new_n766), .C2(new_n767), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n614), .A2(KEYINPUT45), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n614), .A2(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(G469), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n562), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n618), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n777), .A2(KEYINPUT105), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(KEYINPUT105), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n534), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n680), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n766), .A2(new_n767), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n770), .A2(new_n771), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NOR4_X1   g598(.A1(new_n705), .A2(new_n624), .A3(new_n698), .A4(new_n745), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n779), .A2(new_n534), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n786), .B1(new_n779), .B2(new_n534), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND2_X1  g604(.A1(new_n707), .A2(new_n618), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n642), .B(new_n533), .C1(new_n791), .C2(KEYINPUT49), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n736), .A3(new_n761), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT109), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n791), .A2(KEYINPUT49), .ZN(new_n795));
  OR4_X1    g609(.A1(new_n690), .A2(new_n794), .A3(new_n692), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n764), .A2(new_n665), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n732), .A2(new_n736), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n799), .A2(new_n187), .A3(new_n692), .A4(new_n708), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT50), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n787), .A2(new_n788), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n534), .B2(new_n791), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n798), .A3(new_n760), .A4(new_n797), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n760), .A2(new_n709), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT117), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n690), .A2(new_n380), .A3(new_n299), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n529), .A2(new_n636), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n797), .A2(new_n806), .ZN(new_n811));
  INV_X1    g625(.A(new_n742), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n801), .A2(new_n804), .A3(KEYINPUT51), .A4(new_n814), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n797), .A2(new_n755), .A3(new_n806), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT119), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT48), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n637), .ZN(new_n823));
  INV_X1    g637(.A(new_n721), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n297), .B(new_n823), .C1(new_n799), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT118), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n820), .A2(new_n821), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n822), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(new_n818), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n740), .A2(new_n742), .A3(new_n741), .A4(new_n746), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  INV_X1    g646(.A(new_n609), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n608), .B1(new_n607), .B2(new_n602), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n834), .A3(new_n668), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n506), .C1(new_n521), .C2(new_n523), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n745), .A2(new_n569), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n832), .B1(new_n671), .B2(new_n837), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n832), .A2(new_n837), .A3(new_n705), .A4(new_n660), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n758), .B(new_n831), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n756), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  INV_X1    g656(.A(new_n610), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n525), .B2(new_n527), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n295), .A2(new_n289), .A3(new_n303), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n626), .A3(new_n629), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n842), .B1(new_n846), .B2(new_n662), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n304), .A2(new_n637), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n612), .B1(new_n630), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n846), .A2(new_n842), .A3(new_n662), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n841), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n711), .A2(new_n715), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n719), .A2(new_n723), .A3(new_n737), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT110), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n719), .A2(new_n723), .A3(new_n737), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT110), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n716), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n830), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n857), .A2(new_n716), .A3(new_n858), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n857), .B2(new_n716), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n851), .A2(new_n847), .A3(new_n849), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(KEYINPUT113), .A3(new_n865), .A4(new_n841), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n659), .A2(new_n619), .A3(new_n697), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT114), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n674), .A2(new_n693), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n690), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n676), .A3(new_n743), .A4(new_n700), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n676), .A2(new_n743), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(KEYINPUT52), .A3(new_n700), .A4(new_n870), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n861), .A2(new_n866), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n857), .A2(new_n716), .A3(KEYINPUT53), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n853), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n875), .A3(KEYINPUT115), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n871), .A2(new_n883), .A3(new_n872), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n882), .A2(new_n884), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n861), .A3(new_n878), .A4(new_n866), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(KEYINPUT54), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT116), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n890), .A2(new_n895), .A3(new_n892), .A4(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n829), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n796), .B1(new_n897), .B2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n296), .A2(G952), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n239), .A2(new_n241), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n266), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n879), .A2(new_n887), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(G210), .A3(G902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(G902), .A3(new_n285), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n903), .A2(new_n906), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n900), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(G51));
  NAND2_X1  g724(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n889), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n562), .B(KEYINPUT57), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n616), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n886), .B1(new_n878), .B2(new_n877), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n916), .A2(new_n356), .A3(new_n774), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n900), .B1(new_n915), .B2(new_n917), .ZN(G54));
  AND4_X1   g732(.A1(KEYINPUT58), .A2(new_n904), .A3(G475), .A4(G902), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n919), .A2(new_n920), .A3(new_n519), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n919), .B2(new_n519), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n900), .B1(new_n919), .B2(new_n519), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n894), .A2(new_n896), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n634), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n634), .A2(new_n926), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n900), .B1(new_n912), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n937));
  OR2_X1    g751(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n658), .A4(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n372), .B1(new_n916), .B2(new_n940), .ZN(new_n943));
  INV_X1    g757(.A(new_n900), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n916), .A2(new_n940), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT122), .B1(new_n946), .B2(new_n658), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n937), .B(new_n938), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NOR4_X1   g763(.A1(new_n945), .A2(new_n947), .A3(KEYINPUT123), .A4(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  AOI21_X1  g765(.A(new_n296), .B1(new_n301), .B2(G224), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n864), .A2(new_n865), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n296), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n901), .B1(G898), .B2(new_n296), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(new_n955), .Z(G69));
  AOI21_X1  g770(.A(new_n296), .B1(G227), .B2(G900), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n448), .B(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n508), .A2(new_n510), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(new_n960));
  NOR2_X1   g774(.A1(new_n296), .A2(G900), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n874), .A2(new_n700), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n755), .A2(new_n869), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n781), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n758), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n756), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n783), .A2(new_n789), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n961), .B1(new_n967), .B2(new_n296), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n970), .B(new_n961), .C1(new_n967), .C2(new_n296), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n960), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n957), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n874), .A2(new_n695), .A3(new_n700), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT62), .Z(new_n976));
  INV_X1    g790(.A(new_n844), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n680), .B1(new_n977), .B2(new_n712), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n472), .A3(new_n746), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n783), .A2(new_n976), .A3(new_n789), .A4(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n980), .A2(new_n296), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(new_n960), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n972), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n974), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n972), .B(new_n982), .C1(new_n973), .C2(new_n957), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n967), .B2(new_n953), .ZN(new_n989));
  INV_X1    g803(.A(new_n459), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n900), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n988), .B1(new_n980), .B2(new_n953), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n427), .A3(new_n683), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n684), .A2(new_n459), .A3(new_n988), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n890), .A2(new_n892), .A3(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(G57));
endmodule


