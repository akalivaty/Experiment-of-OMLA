//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0002(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI221_X1 g0007(.A(new_n203), .B1(new_n204), .B2(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G50), .B2(G226), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n219), .A2(new_n220), .ZN(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT86), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n252), .B1(G226), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G223), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n204), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n262), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n266), .B2(G232), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(G169), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n230), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G58), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n212), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G58), .A2(G68), .ZN(new_n279));
  OAI21_X1  g0079(.A(G20), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G159), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT79), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT7), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n252), .B2(G20), .ZN(new_n292));
  AOI21_X1  g0092(.A(G20), .B1(new_n284), .B2(new_n286), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(KEYINPUT79), .A3(KEYINPUT7), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n283), .B1(new_n295), .B2(G68), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n276), .B1(new_n296), .B2(KEYINPUT16), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT16), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT80), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n293), .B2(KEYINPUT7), .ZN(new_n300));
  OAI211_X1 g0100(.A(KEYINPUT80), .B(new_n291), .C1(new_n252), .C2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT81), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n284), .B1(new_n286), .B2(new_n303), .ZN(new_n306));
  OAI211_X1 g0106(.A(KEYINPUT7), .B(new_n220), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n212), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n298), .B1(new_n308), .B2(new_n283), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT84), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n276), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  INV_X1    g0114(.A(new_n312), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n275), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT71), .B1(new_n220), .B2(G1), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n219), .A3(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT82), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT8), .B(G58), .Z(new_n325));
  INV_X1    g0125(.A(KEYINPUT82), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n319), .A4(new_n321), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n314), .A2(new_n318), .A3(new_n324), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n323), .A2(new_n315), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT83), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT83), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n328), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n310), .A2(new_n311), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n311), .B1(new_n310), .B2(new_n334), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n272), .B(new_n273), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n268), .A2(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n269), .A2(G190), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n310), .A2(new_n334), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n297), .A2(new_n309), .B1(new_n331), .B2(new_n333), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n343), .A2(KEYINPUT17), .A3(new_n338), .A4(new_n339), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n295), .A2(G68), .ZN(new_n346));
  INV_X1    g0146(.A(new_n283), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n275), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n302), .A2(new_n307), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G68), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT16), .B1(new_n351), .B2(new_n347), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n334), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT84), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n343), .A2(new_n311), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n354), .A2(new_n355), .B1(new_n271), .B2(new_n270), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n251), .B1(new_n345), .B2(new_n359), .ZN(new_n360));
  MUX2_X1   g0160(.A(G222), .B(G223), .S(G1698), .Z(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n252), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n216), .B2(new_n252), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n260), .ZN(new_n365));
  INV_X1    g0165(.A(new_n264), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n266), .A2(G226), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n319), .A2(new_n321), .A3(G50), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT72), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(new_n314), .A3(new_n318), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G50), .B2(new_n312), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n256), .A2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n323), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G150), .ZN(new_n378));
  INV_X1    g0178(.A(new_n281), .ZN(new_n379));
  NOR3_X1   g0179(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n378), .A2(new_n379), .B1(new_n380), .B2(new_n220), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n275), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT69), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n374), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n386));
  INV_X1    g0186(.A(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n370), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n370), .A2(KEYINPUT73), .A3(new_n385), .A4(new_n388), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G238), .A2(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(G232), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n252), .B(new_n393), .C1(new_n394), .C2(G1698), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(new_n260), .C1(G107), .C2(new_n252), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n366), .C1(new_n217), .C2(new_n265), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n387), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G179), .B2(new_n397), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n325), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(new_n376), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n275), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n313), .A2(new_n322), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G77), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n315), .A2(new_n216), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n399), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n391), .A2(new_n392), .A3(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n368), .A2(G190), .B1(new_n384), .B2(KEYINPUT9), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n384), .A2(KEYINPUT9), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n386), .A2(G200), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT10), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n272), .B1(new_n335), .B2(new_n336), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n357), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n342), .A2(new_n344), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT86), .A4(new_n337), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n360), .A2(new_n414), .A3(new_n419), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n266), .A2(G238), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n287), .A2(new_n394), .A3(new_n253), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n252), .A2(G226), .A3(new_n253), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n252), .A2(KEYINPUT75), .A3(G226), .A4(new_n253), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n429), .B(new_n430), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n427), .B(new_n366), .C1(new_n435), .C2(new_n259), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n428), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n260), .ZN(new_n441));
  INV_X1    g0241(.A(new_n437), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n427), .A4(new_n366), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n426), .B1(new_n444), .B2(G169), .ZN(new_n445));
  AOI211_X1 g0245(.A(KEYINPUT14), .B(new_n387), .C1(new_n438), .C2(new_n443), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G179), .A3(new_n443), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OR3_X1    g0249(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n376), .A2(new_n216), .B1(new_n220), .B2(G68), .ZN(new_n451));
  INV_X1    g0251(.A(G50), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n379), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n275), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT11), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n454), .A2(new_n455), .B1(new_n408), .B2(G68), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n315), .A2(new_n212), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n458), .C1(new_n455), .C2(new_n454), .ZN(new_n459));
  XOR2_X1   g0259(.A(new_n459), .B(KEYINPUT78), .Z(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n460), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n444), .A2(G200), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n447), .A2(G190), .A3(new_n443), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT77), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT77), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n447), .A2(new_n443), .A3(new_n466), .A4(G190), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n462), .A2(new_n463), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n397), .A2(G200), .ZN(new_n469));
  INV_X1    g0269(.A(G190), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n411), .B(new_n469), .C1(new_n470), .C2(new_n397), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n461), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n425), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n478), .A2(G264), .A3(new_n259), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n205), .A2(new_n253), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n207), .A2(G1698), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n284), .A2(new_n480), .A3(new_n286), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G294), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n259), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n475), .B(G274), .C1(new_n477), .C2(new_n476), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n479), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G169), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(G179), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n252), .A2(new_n220), .A3(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT22), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT22), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n252), .A2(new_n495), .A3(new_n220), .A4(G87), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT94), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n498), .C1(new_n220), .C2(G107), .ZN(new_n499));
  INV_X1    g0299(.A(G107), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(G20), .C1(KEYINPUT94), .C2(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT88), .A2(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT88), .A2(G116), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n375), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT94), .A2(KEYINPUT23), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT95), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT95), .A4(new_n506), .ZN(new_n510));
  AOI221_X4 g0310(.A(KEYINPUT24), .B1(new_n494), .B2(new_n496), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n494), .A2(new_n496), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n275), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n219), .A2(G33), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n312), .A2(new_n517), .A3(new_n230), .A4(new_n274), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G107), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n315), .A2(new_n500), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT25), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n516), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT96), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n516), .A2(KEYINPUT96), .A3(new_n520), .A4(new_n523), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n492), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G200), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n487), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n487), .A2(G190), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n524), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n315), .A2(new_n206), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n518), .B2(new_n206), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n500), .B1(new_n302), .B2(new_n307), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n206), .A2(new_n500), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n500), .A2(KEYINPUT6), .A3(G97), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n220), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n379), .A2(new_n216), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n538), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n537), .B1(new_n547), .B2(new_n276), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n284), .A2(new_n286), .A3(G244), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(new_n284), .A3(new_n286), .A4(G244), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n284), .A2(new_n286), .A3(G250), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n253), .B1(new_n556), .B2(KEYINPUT4), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n260), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n478), .A2(G257), .A3(new_n259), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n485), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n387), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n558), .A2(new_n369), .A3(new_n485), .A4(new_n559), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n548), .A2(new_n561), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n544), .A2(new_n220), .ZN(new_n567));
  INV_X1    g0367(.A(new_n546), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n285), .A2(G33), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(KEYINPUT81), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(new_n571), .B2(new_n304), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(KEYINPUT7), .B1(new_n300), .B2(new_n301), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n567), .B(new_n568), .C1(new_n573), .C2(new_n500), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n536), .B1(new_n574), .B2(new_n275), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n560), .A2(G200), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n470), .C2(new_n560), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n284), .A2(new_n286), .A3(new_n220), .A4(G68), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT91), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n252), .A2(KEYINPUT91), .A3(new_n220), .A4(G68), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n376), .B2(new_n206), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n220), .B1(new_n428), .B2(new_n583), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n541), .A2(new_n204), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT90), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n275), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n213), .A2(new_n253), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n217), .A2(G1698), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n284), .A2(new_n594), .A3(new_n286), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n503), .A2(G33), .A3(new_n504), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n259), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n475), .A2(new_n263), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n205), .B1(new_n474), .B2(G1), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n599), .A2(new_n259), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n405), .A2(new_n315), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n518), .A2(new_n204), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n593), .A2(new_n602), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n598), .A2(new_n601), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n470), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n403), .A2(new_n404), .A3(new_n519), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n593), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n387), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n598), .A2(new_n601), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n369), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT89), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT89), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n617), .A3(new_n369), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n612), .A2(new_n613), .A3(new_n616), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(KEYINPUT88), .A2(G116), .ZN(new_n622));
  NOR2_X1   g0422(.A1(KEYINPUT88), .A2(G116), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n312), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n518), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G20), .B1(new_n622), .B2(new_n623), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n552), .B(new_n220), .C1(G33), .C2(new_n206), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n275), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n628), .A2(KEYINPUT20), .A3(new_n275), .A4(new_n629), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n625), .B(new_n627), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G303), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n569), .B2(new_n570), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n253), .A2(G257), .ZN(new_n637));
  NAND2_X1  g0437(.A1(G264), .A2(G1698), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n284), .A2(new_n286), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n639), .A3(new_n260), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n478), .A2(G270), .A3(new_n259), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n485), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G169), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT92), .B1(new_n634), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n632), .A2(new_n633), .ZN(new_n645));
  INV_X1    g0445(.A(new_n625), .ZN(new_n646));
  INV_X1    g0446(.A(new_n627), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(G169), .A4(new_n642), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n644), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT93), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT93), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n644), .A2(new_n650), .A3(new_n654), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n640), .A2(G179), .A3(new_n485), .A4(new_n641), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n643), .B2(new_n651), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n648), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n642), .A2(G200), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n634), .B(new_n660), .C1(new_n470), .C2(new_n642), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n621), .A2(new_n656), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n473), .A2(new_n534), .A3(new_n578), .A4(new_n662), .ZN(G372));
  NAND2_X1  g0463(.A1(new_n353), .A2(new_n272), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n460), .B1(G200), .B2(new_n444), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n465), .A2(new_n467), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n461), .A2(new_n413), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n670), .B2(new_n423), .ZN(new_n671));
  INV_X1    g0471(.A(new_n419), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n391), .B(new_n392), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n419), .A2(new_n424), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n461), .A2(new_n468), .A3(new_n471), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n414), .A4(new_n360), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n524), .A2(new_n491), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n656), .A2(new_n659), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n516), .A2(new_n520), .ZN(new_n680));
  INV_X1    g0480(.A(new_n530), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n523), .A3(new_n681), .A4(new_n531), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n609), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n679), .A2(new_n578), .A3(new_n682), .A4(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT26), .B1(new_n566), .B2(new_n620), .ZN(new_n687));
  INV_X1    g0487(.A(new_n561), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n575), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n562), .B(KEYINPUT87), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n685), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n692), .A3(new_n683), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT97), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT97), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n689), .A2(new_n691), .A3(new_n610), .A4(new_n619), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n684), .B1(new_n696), .B2(KEYINPUT26), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(new_n692), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n686), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n674), .B1(new_n677), .B2(new_n700), .ZN(G369));
  NAND2_X1  g0501(.A1(new_n656), .A2(new_n659), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n224), .A2(G20), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n219), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n648), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n703), .A2(new_n661), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n703), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n526), .A2(new_n527), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n710), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n534), .A2(new_n717), .B1(new_n528), .B2(new_n710), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n703), .B2(new_n710), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n710), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n534), .A2(new_n702), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n524), .A2(new_n491), .A3(new_n721), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(G399));
  NOR2_X1   g0525(.A1(new_n225), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n587), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n229), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  INV_X1    g0532(.A(new_n685), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n733), .B2(new_n566), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n566), .A2(new_n620), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n684), .B1(new_n735), .B2(new_n690), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n528), .A2(new_n702), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n682), .A2(new_n566), .A3(new_n577), .A4(new_n610), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n734), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n732), .B1(new_n739), .B2(new_n721), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n693), .A2(KEYINPUT97), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n697), .A2(new_n695), .A3(new_n692), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n710), .B1(new_n743), .B2(new_n686), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n740), .B1(new_n732), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n534), .A2(new_n662), .A3(new_n578), .A4(new_n721), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT98), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n487), .A2(new_n558), .A3(new_n559), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n640), .A2(new_n641), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n614), .A3(G179), .A4(new_n485), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT99), .B(KEYINPUT30), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n607), .A2(new_n657), .ZN(new_n753));
  INV_X1    g0553(.A(new_n559), .ZN(new_n754));
  INV_X1    g0554(.A(new_n552), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n549), .B2(new_n550), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n550), .B1(new_n252), .B2(G250), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n554), .C1(new_n253), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n758), .B2(new_n260), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n753), .A2(new_n759), .A3(KEYINPUT98), .A4(new_n487), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n751), .A2(new_n752), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n753), .A2(new_n759), .A3(KEYINPUT30), .A4(new_n487), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT100), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n479), .A2(new_n484), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n763), .B(new_n485), .C1(new_n759), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n560), .A2(KEYINPUT100), .A3(new_n488), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n607), .A2(new_n369), .A3(new_n642), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n761), .A2(new_n762), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n710), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT31), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n746), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G330), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n745), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n731), .B1(new_n776), .B2(new_n219), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT101), .Z(G364));
  NOR3_X1   g0578(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n712), .B(new_n779), .C1(new_n703), .C2(new_n711), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n230), .B1(G20), .B2(new_n387), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n220), .A2(new_n470), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(G179), .A3(new_n529), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n369), .A2(new_n529), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n784), .A2(G322), .B1(new_n787), .B2(G326), .ZN(new_n788));
  INV_X1    g0588(.A(G294), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n220), .B1(new_n790), .B2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n529), .A2(G179), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT103), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT103), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n788), .B1(new_n789), .B2(new_n791), .C1(new_n797), .C2(new_n635), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n220), .A2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n800), .A2(new_n369), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(new_n792), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n799), .A2(new_n790), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n252), .B1(new_n809), .B2(G329), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n785), .A2(new_n799), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT33), .B(G317), .Z(new_n812));
  OAI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n798), .A2(new_n804), .A3(new_n807), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n796), .A2(G87), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n783), .B(KEYINPUT102), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n277), .B2(new_n817), .C1(new_n500), .C2(new_n805), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n801), .A2(G77), .B1(new_n787), .B2(G50), .ZN(new_n819));
  INV_X1    g0619(.A(new_n811), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G68), .ZN(new_n821));
  INV_X1    g0621(.A(new_n791), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G97), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n819), .A2(new_n252), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n809), .A2(G159), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT32), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n818), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n781), .B1(new_n814), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n229), .A2(G45), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n225), .A2(new_n252), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(new_n249), .C2(new_n474), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n226), .A2(G355), .A3(new_n252), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(G116), .C2(new_n226), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n781), .A2(new_n779), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n704), .A2(G45), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n727), .A2(G1), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n780), .A2(new_n828), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n714), .A2(new_n837), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n713), .A2(G330), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(G396));
  NAND3_X1  g0642(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n710), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n471), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n413), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n412), .A2(new_n721), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT105), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n699), .A2(new_n721), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT106), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n849), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n852), .B2(new_n744), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(new_n775), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n775), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n837), .A3(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n783), .A2(new_n789), .B1(new_n805), .B2(new_n204), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n823), .B1(new_n635), .B2(new_n786), .C1(new_n797), .C2(new_n500), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(G283), .C2(new_n820), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n252), .B1(new_n809), .B2(G311), .ZN(new_n860));
  INV_X1    g0660(.A(new_n624), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n802), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT104), .Z(new_n863));
  NAND2_X1  g0663(.A1(new_n816), .A2(G143), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G137), .A2(new_n787), .B1(new_n820), .B2(G150), .ZN(new_n865));
  INV_X1    g0665(.A(G159), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n802), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT34), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n867), .A2(new_n868), .B1(G132), .B2(new_n809), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n287), .B1(new_n822), .B2(G58), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n805), .A2(new_n212), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G50), .B2(new_n796), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n781), .B1(new_n863), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n849), .ZN(new_n877));
  NOR2_X1   g0677(.A1(G13), .A2(G33), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n837), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n781), .A2(new_n878), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n876), .B(new_n879), .C1(G77), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n856), .A2(new_n882), .ZN(G384));
  NAND3_X1  g0683(.A1(new_n450), .A2(new_n460), .A3(new_n710), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n460), .A2(new_n710), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n468), .B(new_n885), .C1(new_n886), .C2(new_n462), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n850), .B2(new_n847), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n329), .B(new_n328), .C1(new_n349), .C2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n708), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n422), .B1(new_n356), .B2(new_n273), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n421), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n335), .A2(new_n336), .B1(new_n272), .B2(new_n894), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n340), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n272), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n895), .A3(new_n340), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n891), .B1(new_n897), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n421), .A2(new_n423), .A3(new_n337), .ZN(new_n907));
  INV_X1    g0707(.A(new_n895), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n890), .A2(new_n911), .B1(new_n667), .B2(new_n708), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n708), .B1(new_n354), .B2(new_n355), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n664), .A2(new_n340), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT37), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT108), .B(KEYINPUT37), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n900), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n914), .B1(new_n667), .B2(new_n422), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI221_X4 g0722(.A(new_n891), .B1(new_n900), .B2(new_n903), .C1(new_n907), .C2(new_n908), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n913), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n461), .A2(new_n710), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n906), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n912), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT109), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n745), .B2(new_n677), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n699), .A2(new_n732), .A3(new_n721), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n739), .A2(new_n721), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT29), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT109), .A3(new_n473), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n673), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n928), .B(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n772), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n770), .A2(KEYINPUT110), .A3(new_n771), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n746), .A2(new_n941), .A3(new_n773), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT111), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n746), .A2(new_n941), .A3(KEYINPUT111), .A4(new_n773), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n888), .A2(new_n849), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n911), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n920), .A2(new_n921), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n891), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n910), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n947), .B1(new_n944), .B2(new_n945), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT40), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(G330), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n946), .A2(G330), .A3(new_n473), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n951), .A2(new_n946), .A3(new_n956), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n677), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n937), .B(new_n961), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n219), .B2(new_n704), .ZN(new_n963));
  OAI21_X1  g0763(.A(G77), .B1(new_n277), .B2(new_n212), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n964), .A2(new_n229), .B1(G50), .B2(new_n212), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(G1), .A3(new_n224), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT35), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n220), .B(new_n230), .C1(new_n544), .C2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n968), .B(G116), .C1(new_n967), .C2(new_n544), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT107), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT36), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n963), .A2(new_n966), .A3(new_n971), .ZN(G367));
  INV_X1    g0772(.A(KEYINPUT113), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n578), .B1(new_n575), .B2(new_n721), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n566), .B2(new_n721), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT112), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n722), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT42), .ZN(new_n978));
  INV_X1    g0778(.A(new_n528), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n566), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n721), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n593), .A2(new_n603), .A3(new_n605), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n710), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n683), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n685), .B2(new_n983), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n978), .A2(new_n981), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT43), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n978), .A2(new_n981), .A3(new_n991), .A4(new_n985), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n720), .A2(new_n976), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n973), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n836), .A2(G1), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n976), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n722), .A2(new_n724), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n715), .A2(new_n719), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n723), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n776), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n776), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n726), .B(KEYINPUT41), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n999), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n990), .A2(new_n992), .A3(KEYINPUT113), .A4(new_n994), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n996), .A2(new_n997), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n811), .A2(new_n866), .B1(new_n805), .B2(new_n216), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n784), .A2(G150), .B1(new_n787), .B2(G143), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n452), .B2(new_n802), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1017), .B(new_n1019), .C1(G137), .C2(new_n809), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n822), .A2(G68), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n796), .A2(G58), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1020), .A2(new_n252), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(G317), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n808), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n287), .B1(new_n805), .B2(new_n206), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n861), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT46), .B1(new_n797), .B2(new_n626), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1025), .B(new_n1026), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n822), .A2(G107), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n816), .A2(G303), .B1(G294), .B2(new_n820), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n801), .A2(G283), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n786), .A2(new_n803), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n781), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n985), .A2(new_n779), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n830), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n834), .B1(new_n226), .B2(new_n405), .C1(new_n241), .C2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n838), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1016), .A2(new_n1041), .ZN(G387));
  AOI22_X1  g0842(.A1(G322), .A2(new_n787), .B1(new_n820), .B2(G311), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n635), .B2(new_n802), .C1(new_n817), .C2(new_n1024), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT48), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n806), .B2(new_n791), .C1(new_n789), .C2(new_n797), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT49), .Z(new_n1047));
  AOI21_X1  g0847(.A(new_n252), .B1(new_n809), .B2(G326), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n861), .B2(new_n805), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n802), .A2(new_n212), .B1(new_n783), .B2(new_n452), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n405), .A2(new_n791), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n811), .A2(new_n323), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n786), .A2(new_n866), .B1(new_n805), .B2(new_n206), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n796), .A2(G77), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n287), .B(new_n1057), .C1(G150), .C2(new_n809), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n781), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n325), .A2(new_n452), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT50), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n212), .A2(new_n216), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n728), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1061), .A2(G45), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n830), .B1(new_n237), .B2(new_n474), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n226), .A3(new_n252), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n226), .A2(G107), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n834), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n837), .B1(new_n718), .B2(new_n779), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1059), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1009), .A2(new_n776), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n726), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1071), .B1(new_n999), .B2(new_n1009), .C1(new_n1073), .C2(new_n1010), .ZN(G393));
  NAND2_X1  g0874(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1007), .B(new_n720), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n726), .B(new_n1075), .C1(new_n1076), .C2(new_n1010), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n976), .A2(new_n779), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n834), .B1(new_n206), .B2(new_n226), .C1(new_n246), .C2(new_n1039), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n783), .A2(new_n803), .B1(new_n786), .B2(new_n1024), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G303), .B2(new_n820), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n802), .A2(new_n789), .B1(new_n500), .B2(new_n805), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n252), .B(new_n1083), .C1(G322), .C2(new_n809), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(new_n806), .C2(new_n797), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n624), .B2(new_n822), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n801), .A2(new_n325), .B1(new_n820), .B2(G50), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT115), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G68), .B2(new_n796), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n822), .A2(G77), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n805), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G87), .A2(new_n1091), .B1(new_n809), .B2(G143), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n783), .A2(new_n866), .B1(new_n786), .B2(new_n378), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  NOR3_X1   g0895(.A1(new_n1093), .A2(new_n287), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n781), .B1(new_n1086), .B2(new_n1096), .ZN(new_n1097));
  AND4_X1   g0897(.A1(new_n838), .A2(new_n1078), .A3(new_n1079), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1076), .B2(new_n998), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1077), .A2(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n850), .A2(new_n847), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n888), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n925), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n924), .B2(new_n926), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n922), .A2(new_n923), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n849), .A2(new_n739), .A3(new_n721), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n889), .B1(new_n1106), .B2(new_n847), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1105), .A2(new_n1107), .A3(new_n925), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n774), .A2(new_n888), .A3(G330), .A4(new_n849), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G330), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n944), .B2(new_n945), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n948), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT39), .B1(new_n953), .B2(new_n910), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n926), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n890), .B2(new_n925), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1106), .A2(new_n847), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n954), .B(new_n1103), .C1(new_n889), .C2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1114), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1110), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n958), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1112), .A2(KEYINPUT116), .A3(new_n473), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1101), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n774), .A2(G330), .A3(new_n849), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n889), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1118), .A2(new_n1109), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n946), .A2(new_n852), .A3(G330), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n889), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1125), .B(new_n936), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1112), .A2(new_n948), .B1(new_n889), .B2(new_n1127), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n888), .B1(new_n1112), .B2(new_n852), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1136), .A2(new_n1126), .B1(new_n1137), .B2(new_n1130), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1138), .A2(KEYINPUT117), .A3(new_n936), .A4(new_n1125), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1135), .A2(KEYINPUT119), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT119), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1121), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1121), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(KEYINPUT118), .A3(new_n726), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT118), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1121), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n727), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1142), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1144), .A2(new_n998), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  AOI21_X1  g0952(.A(new_n287), .B1(new_n801), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n784), .A2(G132), .B1(new_n822), .B2(G159), .ZN(new_n1154));
  INV_X1    g0954(.A(G125), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1153), .B(new_n1154), .C1(new_n1155), .C2(new_n808), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n796), .A2(G150), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT53), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G50), .C2(new_n1091), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1160), .B2(new_n786), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G137), .B2(new_n820), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n815), .B1(new_n626), .B2(new_n783), .C1(new_n806), .C2(new_n786), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G294), .B2(new_n809), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1090), .B1(new_n500), .B2(new_n811), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n872), .B(new_n1165), .C1(G97), .C2(new_n801), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n287), .A3(new_n1166), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT120), .Z(new_n1168));
  OAI21_X1  g0968(.A(new_n781), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n838), .C1(new_n325), .C2(new_n881), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT121), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n878), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1150), .A2(new_n1151), .A3(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n419), .A2(new_n389), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n384), .A2(new_n708), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1175), .B(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n957), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n951), .A2(G330), .A3(new_n956), .A4(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1180), .A2(new_n928), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n928), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1125), .A2(new_n936), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1148), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1185), .B(KEYINPUT57), .C1(new_n1148), .C2(new_n1186), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n726), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n405), .A2(new_n802), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1091), .A2(G58), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n820), .A2(G97), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n809), .B2(G283), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1056), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1192), .B(new_n1196), .C1(G107), .C2(new_n784), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n787), .A2(G116), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n287), .A3(new_n1021), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n258), .B1(new_n285), .B2(new_n256), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1199), .A2(new_n1200), .B1(new_n452), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT122), .ZN(new_n1203));
  INV_X1    g1003(.A(G132), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n811), .A2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n783), .A2(new_n1160), .B1(new_n791), .B2(new_n378), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n796), .C2(new_n1152), .ZN(new_n1207));
  INV_X1    g1007(.A(G137), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1207), .B1(new_n1155), .B2(new_n786), .C1(new_n1208), .C2(new_n802), .ZN(new_n1209));
  XOR2_X1   g1009(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1210));
  XOR2_X1   g1010(.A(new_n1209), .B(new_n1210), .Z(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n866), .B2(new_n805), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1211), .A2(new_n1213), .B1(new_n1200), .B2(new_n1199), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n781), .B1(new_n1203), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n838), .C1(G50), .C2(new_n881), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n878), .B2(new_n1181), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT124), .Z(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1185), .B2(new_n998), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1191), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1138), .A2(new_n998), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n889), .A2(new_n878), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n880), .A2(new_n212), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n786), .A2(new_n789), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n796), .A2(G97), .B1(G303), .B2(new_n809), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT125), .Z(new_n1226));
  AOI211_X1 g1026(.A(new_n252), .B(new_n1052), .C1(G77), .C2(new_n1091), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n801), .A2(G107), .B1(new_n820), .B2(new_n624), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1224), .B(new_n1229), .C1(G283), .C2(new_n784), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n287), .B1(new_n820), .B2(new_n1152), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n1208), .B2(new_n817), .C1(new_n797), .C2(new_n866), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n808), .A2(new_n1160), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n802), .A2(new_n378), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1193), .B1(new_n452), .B2(new_n791), .C1(new_n1204), .C2(new_n786), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n781), .B1(new_n1230), .B2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1222), .A2(new_n838), .A3(new_n1223), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1221), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1186), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1240), .B1(new_n1243), .B2(new_n1013), .ZN(G381));
  OR2_X1    g1044(.A1(G375), .A2(G378), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1245), .A2(G384), .A3(G381), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1016), .A2(new_n1041), .A3(new_n1099), .A4(new_n1077), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1247), .A2(G396), .A3(G393), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND2_X1  g1050(.A1(G375), .A2(G378), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1012), .B1(new_n1148), .B2(new_n1186), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n999), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1217), .B1(new_n1253), .B2(new_n1185), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1254), .A2(new_n1151), .A3(new_n1150), .A4(new_n1173), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1186), .A2(new_n1241), .A3(KEYINPUT60), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1135), .A2(KEYINPUT60), .A3(new_n1139), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n727), .B(new_n1256), .C1(new_n1257), .C2(new_n1242), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n882), .B(new_n856), .C1(new_n1258), .C2(new_n1239), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1256), .B1(new_n1257), .B2(new_n1242), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n726), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(G384), .A3(new_n1240), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n709), .A2(G213), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1251), .A2(new_n1255), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1251), .A2(new_n1264), .A3(new_n1255), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n709), .A2(G213), .A3(G2897), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT126), .Z(new_n1269));
  AND3_X1   g1069(.A1(new_n1259), .A2(new_n1262), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G375), .A2(G378), .B1(G213), .B2(new_n709), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1263), .A4(new_n1255), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1266), .A2(new_n1273), .A3(new_n1274), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(G390), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1247), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G393), .B(G396), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1281), .A3(new_n1247), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1273), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1285), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1267), .A2(new_n1272), .A3(KEYINPUT127), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1288), .A2(new_n1274), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1265), .B(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1291), .B2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1285), .A2(new_n1245), .A3(new_n1251), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1263), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1263), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(G402));
endmodule


