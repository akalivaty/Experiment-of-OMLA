//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n461), .A2(new_n462), .ZN(new_n465));
  AOI211_X1 g040(.A(new_n464), .B(new_n465), .C1(new_n456), .C2(G2106), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  NAND2_X1  g054(.A1(G101), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n473), .A2(new_n481), .ZN(G160));
  AOI21_X1  g057(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G138), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  AOI22_X1  g067(.A1(G126), .A2(new_n483), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n485), .A2(KEYINPUT4), .A3(G138), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT69), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT70), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n499), .A2(KEYINPUT70), .A3(new_n501), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n493), .B(new_n494), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT71), .A3(G543), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(new_n510), .B1(KEYINPUT5), .B2(new_n507), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR3_X1    g089(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(new_n517), .A2(G89), .ZN(new_n523));
  AND3_X1   g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n518), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G51), .Z(new_n526));
  OAI221_X1 g101(.A(new_n523), .B1(KEYINPUT7), .B2(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n511), .A2(G63), .ZN(new_n528));
  NAND3_X1  g103(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n514), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n517), .A2(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n525), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n514), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(new_n517), .A2(G81), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT74), .B(G43), .Z(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n514), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT75), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT76), .ZN(G188));
  NAND2_X1  g125(.A1(new_n518), .A2(G53), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT9), .Z(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n508), .A2(new_n510), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT78), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n511), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT79), .B(G65), .Z(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n514), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n511), .A2(G91), .A3(new_n516), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT77), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n553), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  OAI21_X1  g144(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n518), .A2(G49), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n511), .A2(G87), .A3(new_n516), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n511), .A2(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n514), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n518), .A2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n511), .A2(G86), .A3(new_n516), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n517), .A2(G85), .B1(G47), .B2(new_n518), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n514), .B2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n557), .A2(G66), .A3(new_n559), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT80), .Z(new_n589));
  AOI21_X1  g164(.A(new_n514), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(G54), .B2(new_n518), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n517), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  AND2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n586), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT81), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g182(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT82), .Z(new_n613));
  AOI22_X1  g188(.A1(G123), .A2(new_n483), .B1(new_n485), .B2(G135), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n616), .B(new_n617), .C1(G111), .C2(new_n467), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n610), .A2(new_n611), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n613), .A2(new_n620), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2438), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G14), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XOR2_X1   g213(.A(G2067), .B(G2678), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(new_n611), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  AOI21_X1  g222(.A(KEYINPUT18), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(G227));
  XOR2_X1   g224(.A(G1956), .B(G2474), .Z(new_n650));
  XOR2_X1   g225(.A(G1961), .B(G1966), .Z(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n651), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n661), .C1(new_n659), .C2(new_n658), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G1986), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1991), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT22), .B(G1981), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G229));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n670));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G23), .ZN(new_n672));
  INV_X1    g247(.A(G288), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n673), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT33), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT87), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(G6), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n581), .B2(new_n671), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT32), .B(G1981), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G16), .A2(G22), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G166), .B2(G16), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT88), .B(G1971), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n682), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n682), .B2(new_n686), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n691));
  MUX2_X1   g266(.A(G24), .B(G290), .S(G16), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G1986), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(G1986), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G119), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n485), .A2(G131), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n698));
  NOR2_X1   g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT85), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n694), .A2(new_n695), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n690), .A2(new_n691), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n691), .B1(new_n690), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n670), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(KEYINPUT36), .A3(new_n709), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(KEYINPUT98), .B1(G29), .B2(G32), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT96), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n483), .A2(G129), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n718), .B(new_n719), .C1(G141), .C2(new_n485), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(new_n716), .B(KEYINPUT98), .S(new_n726), .Z(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  OR2_X1    g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n725), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n619), .B2(new_n725), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT99), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(G29), .A2(G33), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT25), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n485), .A2(G139), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n467), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n725), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n737), .B(new_n746), .C1(new_n727), .C2(new_n729), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G19), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n543), .B2(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G1341), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n725), .A2(G26), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n483), .A2(G128), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n485), .A2(G140), .ZN(new_n753));
  NOR2_X1   g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n756), .B2(G29), .ZN(new_n757));
  MUX2_X1   g332(.A(new_n751), .B(new_n757), .S(KEYINPUT28), .Z(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT91), .B(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G168), .A2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G16), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NOR2_X1   g338(.A1(G5), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G171), .B2(G16), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(G1961), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n747), .A2(new_n750), .A3(new_n760), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(G164), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G27), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n771), .B1(G1341), .B2(new_n749), .C1(G1961), .C2(new_n765), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n735), .A2(new_n736), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n744), .A2(new_n745), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n773), .B1(new_n774), .B2(new_n775), .C1(new_n762), .C2(new_n763), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n767), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n774), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n769), .A2(new_n770), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(KEYINPUT24), .A2(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g359(.A1(G160), .A2(G29), .B1(KEYINPUT92), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(KEYINPUT92), .B2(new_n784), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT93), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2084), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT94), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n671), .A2(KEYINPUT23), .A3(G20), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n791));
  INV_X1    g366(.A(G20), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G16), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n793), .C1(new_n598), .C2(new_n671), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n671), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n594), .B2(new_n671), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT90), .B(G1348), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n789), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n780), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n787), .A2(G2084), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n715), .A2(new_n730), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n725), .A2(G35), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n725), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT29), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(KEYINPUT29), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n807), .A2(new_n808), .B1(KEYINPUT100), .B2(G2090), .ZN(new_n809));
  NAND2_X1  g384(.A1(KEYINPUT100), .A2(G2090), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n804), .A2(new_n811), .ZN(G311));
  OR2_X1    g387(.A1(new_n804), .A2(new_n811), .ZN(G150));
  AOI22_X1  g388(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(G651), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT102), .B(G93), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n517), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n518), .A2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(G860), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n591), .A2(new_n593), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n601), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT39), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT103), .B1(new_n817), .B2(new_n821), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n816), .A2(G651), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n830), .A2(new_n831), .A3(new_n820), .A4(new_n819), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n832), .C1(new_n542), .C2(new_n540), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n817), .A2(new_n821), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n831), .A3(new_n543), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n828), .B(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n823), .B1(new_n837), .B2(G860), .ZN(G145));
  XNOR2_X1  g413(.A(new_n724), .B(new_n701), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n485), .A2(G142), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT105), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n483), .A2(G130), .ZN(new_n842));
  OR2_X1    g417(.A1(G106), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(KEYINPUT105), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n841), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n839), .B(new_n846), .Z(new_n847));
  XNOR2_X1  g422(.A(G160), .B(new_n619), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n489), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n743), .B(new_n756), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n847), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n504), .B(new_n609), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(new_n855), .A3(new_n853), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(G395));
  XNOR2_X1  g442(.A(new_n836), .B(new_n603), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n594), .A2(new_n598), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n824), .A2(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT107), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n869), .A2(KEYINPUT41), .A3(new_n870), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT41), .B1(new_n869), .B2(new_n870), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n868), .A2(new_n879), .A3(new_n872), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(G305), .B(G288), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G290), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G166), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n874), .A2(new_n878), .A3(new_n887), .A4(new_n880), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n882), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n882), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g467(.A(new_n891), .B1(G868), .B2(new_n834), .ZN(G331));
  XNOR2_X1  g468(.A(G168), .B(G171), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n836), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n833), .A2(new_n835), .A3(new_n894), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n896), .B(new_n897), .C1(new_n875), .C2(new_n876), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n894), .B1(new_n833), .B2(new_n835), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n871), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n886), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n901), .A3(new_n885), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n858), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n903), .A2(new_n904), .A3(new_n907), .A4(new_n858), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(KEYINPUT108), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT44), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n908), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(G397));
  INV_X1    g490(.A(KEYINPUT125), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT117), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n570), .A2(new_n571), .A3(G1976), .A4(new_n573), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT114), .ZN(new_n919));
  AND2_X1   g494(.A1(KEYINPUT109), .A2(G40), .ZN(new_n920));
  NOR2_X1   g495(.A1(KEYINPUT109), .A2(G40), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n473), .A2(new_n481), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n504), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n919), .A2(G8), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT115), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n673), .A2(G1976), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n926), .B(new_n927), .C1(KEYINPUT52), .C2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(G8), .A3(new_n925), .A4(new_n919), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n919), .A2(new_n927), .A3(G8), .A4(new_n925), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT49), .ZN(new_n935));
  INV_X1    g510(.A(new_n577), .ZN(new_n936));
  INV_X1    g511(.A(G1981), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n579), .A4(new_n578), .ZN(new_n938));
  OAI21_X1  g513(.A(G1981), .B1(new_n577), .B2(new_n580), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n940), .B2(KEYINPUT116), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT116), .ZN(new_n942));
  AOI211_X1 g517(.A(new_n942), .B(KEYINPUT49), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n925), .A2(G8), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n917), .B1(new_n934), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n929), .B2(new_n933), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT117), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n504), .A2(new_n924), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n923), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1971), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n504), .A2(new_n956), .A3(new_n924), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n957), .A2(new_n923), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n504), .B2(new_n924), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT111), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n961), .B(new_n956), .C1(new_n504), .C2(new_n924), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT112), .B(G2090), .Z(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G303), .A2(G8), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n968), .A3(G8), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n946), .A2(new_n948), .A3(new_n970), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n945), .A2(G1976), .A3(G288), .ZN(new_n972));
  NOR2_X1   g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  OAI211_X1 g548(.A(G8), .B(new_n925), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT63), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n953), .A2(new_n763), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT118), .B(G2084), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n963), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(G8), .A3(G168), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n970), .A2(new_n976), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n965), .A2(G8), .ZN(new_n983));
  INV_X1    g558(.A(new_n968), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n982), .A2(new_n946), .A3(new_n948), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n957), .A2(new_n923), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n987), .A2(new_n959), .A3(new_n964), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n954), .B2(new_n953), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n947), .A2(new_n991), .A3(new_n969), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n976), .B1(new_n992), .B2(new_n981), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n975), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n795), .B1(new_n987), .B2(new_n959), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT119), .B(new_n795), .C1(new_n987), .C2(new_n959), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n504), .B2(new_n924), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT56), .B(G2072), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n923), .A4(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n951), .A2(new_n923), .A3(new_n952), .A4(new_n1004), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT120), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n553), .B2(new_n566), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n552), .A2(new_n563), .A3(new_n565), .A4(KEYINPUT57), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n999), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n925), .A2(G2067), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n961), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n959), .A2(KEYINPUT111), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n987), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1019), .B2(G1348), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1013), .A2(new_n594), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n999), .A2(new_n1008), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT60), .B(new_n1015), .C1(new_n1019), .C2(G1348), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1348), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1014), .B1(new_n963), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n594), .B1(new_n1030), .B2(KEYINPUT60), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT61), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n999), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1012), .B1(new_n999), .B2(new_n1008), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(G1996), .ZN(new_n1040));
  INV_X1    g615(.A(new_n925), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT58), .B(G1341), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n953), .A2(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n543), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT59), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1035), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT122), .B1(new_n1048), .B2(KEYINPUT61), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1024), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n1013), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1025), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n980), .B2(G286), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n977), .B(G168), .C1(new_n963), .C2(new_n979), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1054), .B1(new_n1056), .B2(G8), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT124), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n953), .B2(G2078), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1002), .A2(KEYINPUT53), .A3(new_n770), .A4(new_n923), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1062), .B(new_n1063), .C1(new_n1019), .C2(G1961), .ZN(new_n1064));
  XOR2_X1   g639(.A(G171), .B(KEYINPUT54), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AND4_X1   g641(.A1(new_n1066), .A2(new_n947), .A3(new_n991), .A4(new_n969), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1068), .B(new_n1069), .C1(new_n1057), .C2(new_n1055), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n770), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n473), .A2(new_n481), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1065), .B1(new_n1002), .B2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1062), .C1(G1961), .C2(new_n1019), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1060), .A2(new_n1067), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n916), .B(new_n994), .C1(new_n1053), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1044), .B(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1024), .A2(new_n1013), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1036), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n1013), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n824), .B1(new_n1020), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT123), .B1(new_n1030), .B2(KEYINPUT60), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1080), .A2(new_n1083), .A3(new_n1090), .A4(new_n1050), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1025), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1075), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n986), .A2(new_n993), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n971), .A2(new_n974), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT125), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1060), .A2(KEYINPUT62), .A3(new_n1070), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT62), .B1(new_n1060), .B2(new_n1070), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n992), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(G171), .A3(new_n1064), .A4(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1076), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1001), .A2(new_n923), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT110), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2067), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n756), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(G1996), .B2(new_n724), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1104), .ZN(new_n1111));
  INV_X1    g686(.A(G1996), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1106), .A2(new_n1110), .B1(new_n724), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n701), .B(new_n703), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n1105), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(G290), .B(G1986), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1103), .A2(new_n1119), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1114), .A2(new_n701), .A3(new_n703), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n756), .A2(G2067), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1106), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1113), .B(KEYINPUT46), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1105), .B1(new_n724), .B2(new_n1109), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT126), .Z(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT47), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1104), .A2(G1986), .A3(G290), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT48), .Z(new_n1130));
  AOI211_X1 g705(.A(new_n1123), .B(new_n1128), .C1(new_n1116), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1120), .A2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g707(.A(G319), .ZN(new_n1134));
  NOR2_X1   g708(.A1(G227), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g709(.A1(new_n668), .A2(new_n636), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n1137));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g712(.A(new_n1138), .B1(new_n908), .B2(new_n906), .ZN(new_n1139));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n860), .A3(new_n1140), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


