//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n221), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  AND2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  OAI211_X1 g0049(.A(G222), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  OAI211_X1 g0050(.A(G223), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OR2_X1    g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n250), .B(new_n251), .C1(new_n252), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n258), .A3(G274), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n260), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(KEYINPUT70), .A3(G200), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n258), .A2(new_n265), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n264), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n259), .B2(new_n256), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT10), .B1(new_n274), .B2(G190), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n269), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT9), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n220), .A2(KEYINPUT8), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT8), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT66), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n207), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(new_n207), .A3(G33), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n284), .A2(new_n287), .A3(new_n289), .A4(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n216), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G50), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n206), .B2(G20), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(G50), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n279), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n297), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n292), .B2(new_n294), .ZN(new_n305));
  INV_X1    g0105(.A(new_n302), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT9), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT69), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n298), .A2(new_n279), .A3(new_n302), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT9), .B1(new_n305), .B2(new_n306), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT69), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n278), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n278), .A2(new_n308), .A3(KEYINPUT71), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n274), .A2(G190), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n317), .B1(new_n275), .B2(new_n274), .C1(new_n303), .C2(new_n307), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n315), .A2(new_n316), .B1(KEYINPUT10), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n305), .A2(new_n306), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n268), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n274), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT72), .B1(new_n299), .B2(G68), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT12), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(G68), .B2(new_n301), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n289), .A2(G77), .A3(new_n291), .ZN(new_n330));
  INV_X1    g0130(.A(G68), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n293), .A2(G50), .B1(G20), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n304), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n255), .A2(G232), .A3(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  OAI211_X1 g0140(.A(G226), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n259), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n258), .A2(G274), .ZN(new_n344));
  AOI22_X1  g0144(.A1(G238), .A2(new_n266), .B1(new_n344), .B2(new_n263), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n343), .B2(new_n345), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n338), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n345), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G179), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n338), .B1(new_n355), .B2(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n337), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G200), .B1(new_n347), .B2(new_n348), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n351), .A2(G190), .A3(new_n352), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n358), .A2(new_n359), .A3(new_n336), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n253), .A2(new_n207), .A3(new_n254), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n254), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n331), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n220), .A2(new_n331), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n201), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n293), .A2(G159), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n363), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n248), .A2(new_n249), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n374), .B2(new_n207), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n248), .A2(new_n249), .A3(new_n365), .A4(G20), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n372), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n379), .A3(new_n297), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n285), .A2(new_n286), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n301), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n299), .B1(new_n381), .B2(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(G223), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n389));
  OAI211_X1 g0189(.A(G226), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n259), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n258), .A2(G232), .A3(new_n265), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n264), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n393), .A2(new_n323), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n259), .B2(new_n392), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(G169), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n388), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT18), .ZN(new_n402));
  INV_X1    g0202(.A(G190), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n393), .A2(new_n403), .A3(new_n396), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G200), .B2(new_n398), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n380), .A2(new_n405), .A3(new_n387), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n399), .B1(new_n380), .B2(new_n387), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n380), .A2(new_n405), .A3(new_n387), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n402), .A2(new_n407), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n266), .A2(G244), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n264), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT68), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n255), .A2(G232), .A3(new_n247), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n255), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n259), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT68), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n423), .A3(new_n264), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n417), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n425), .A2(G200), .ZN(new_n426));
  INV_X1    g0226(.A(new_n299), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n252), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n384), .B2(new_n252), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(new_n288), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n283), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n304), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n425), .B2(new_n403), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n425), .A2(G179), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n425), .B2(new_n321), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n362), .A2(new_n414), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n326), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G264), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n444));
  OAI211_X1 g0244(.A(G257), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n253), .A2(G303), .A3(new_n254), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n259), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n261), .B2(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n262), .A2(G1), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n451), .B2(KEYINPUT77), .ZN(new_n454));
  OAI211_X1 g0254(.A(G270), .B(new_n258), .C1(new_n452), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n206), .A2(G45), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n449), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(new_n451), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n344), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n448), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G200), .ZN(new_n462));
  INV_X1    g0262(.A(G33), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT74), .B1(new_n463), .B2(G1), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n464), .A2(new_n299), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT74), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n206), .A3(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n304), .A3(G116), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n299), .A2(G116), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n296), .A2(new_n216), .B1(G20), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(new_n207), .C1(G33), .C2(new_n222), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT20), .B1(new_n472), .B2(new_n474), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n468), .B(new_n470), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n448), .A2(new_n455), .A3(G190), .A4(new_n460), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n462), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT79), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n462), .A2(new_n479), .A3(new_n483), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n461), .A2(new_n478), .A3(KEYINPUT21), .A4(G169), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT78), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n464), .A2(new_n467), .A3(new_n299), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n297), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n469), .B1(new_n489), .B2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n472), .A2(new_n474), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n475), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n321), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT78), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT21), .A4(new_n461), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n461), .A2(new_n478), .A3(G169), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n448), .A2(new_n455), .A3(G179), .A4(new_n460), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(new_n499), .B1(new_n501), .B2(new_n478), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n485), .A2(new_n487), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n505), .B1(G33), .B2(G283), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(G1698), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(G244), .C1(new_n249), .C2(new_n248), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT75), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n255), .A2(KEYINPUT75), .A3(G244), .A4(new_n507), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G250), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT76), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT76), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n255), .A2(new_n515), .A3(G250), .A4(G1698), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n259), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n258), .B1(new_n452), .B2(new_n454), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n460), .B1(new_n519), .B2(new_n223), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n323), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n299), .A2(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n489), .B2(G97), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n420), .B1(new_n366), .B2(new_n367), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT73), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  AND2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n527), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(G97), .A4(new_n420), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n207), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n252), .A2(G20), .A3(G33), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n525), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n524), .B1(new_n538), .B2(new_n304), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n514), .A2(new_n516), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(new_n506), .A3(new_n510), .A4(new_n511), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n520), .B1(new_n541), .B2(new_n259), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n522), .B(new_n539), .C1(G169), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n518), .A2(G190), .A3(new_n521), .ZN(new_n544));
  INV_X1    g0344(.A(new_n524), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n532), .A2(new_n535), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n537), .B1(new_n546), .B2(G20), .ZN(new_n547));
  OAI21_X1  g0347(.A(G107), .B1(new_n375), .B2(new_n376), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n549), .B2(new_n297), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n544), .B(new_n550), .C1(new_n275), .C2(new_n542), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n553));
  OAI211_X1 g0353(.A(G238), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n259), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n258), .A2(G274), .A3(new_n453), .ZN(new_n558));
  INV_X1    g0358(.A(G250), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n206), .B2(G45), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n258), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n207), .B1(new_n340), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n530), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n207), .B(G68), .C1(new_n248), .C2(new_n249), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n288), .B2(new_n222), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n297), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n489), .A2(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n430), .A2(new_n427), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n562), .B1(new_n556), .B2(new_n259), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n565), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n323), .ZN(new_n581));
  INV_X1    g0381(.A(new_n430), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n489), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n574), .A2(new_n583), .A3(new_n576), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n581), .B(new_n584), .C1(G169), .C2(new_n578), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n259), .B1(new_n458), .B2(new_n459), .ZN(new_n587));
  OAI211_X1 g0387(.A(G257), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n587), .A2(G264), .B1(new_n591), .B2(new_n259), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(G179), .A3(new_n460), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n259), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(new_n258), .C1(new_n452), .C2(new_n454), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n460), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n207), .B(G87), .C1(new_n248), .C2(new_n249), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n255), .A2(new_n601), .A3(new_n207), .A4(G87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n207), .B2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n420), .A2(KEYINPUT23), .A3(G20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT24), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n603), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n304), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT25), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n299), .B2(G107), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n427), .A2(KEYINPUT25), .A3(new_n420), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n489), .A2(G107), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n598), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  AOI211_X1 g0421(.A(KEYINPUT24), .B(new_n609), .C1(new_n600), .C2(new_n602), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n613), .B1(new_n603), .B2(new_n610), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n297), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(G200), .B1(new_n592), .B2(new_n460), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n596), .A2(G190), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n624), .B(new_n619), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n586), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n503), .A2(new_n552), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n443), .A2(new_n629), .ZN(G372));
  AND4_X1   g0430(.A1(KEYINPUT80), .A2(new_n574), .A3(new_n575), .A4(new_n576), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n573), .A2(new_n297), .B1(new_n427), .B2(new_n430), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT80), .B1(new_n632), .B2(new_n575), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n565), .A2(new_n579), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n585), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n543), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  AOI211_X1 g0438(.A(G179), .B(new_n562), .C1(new_n259), .C2(new_n556), .ZN(new_n639));
  AOI21_X1  g0439(.A(G169), .B1(new_n557), .B2(new_n563), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n637), .A2(new_n638), .B1(new_n584), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n543), .A2(new_n551), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT80), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n632), .A2(KEYINPUT80), .A3(new_n575), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n578), .A2(new_n275), .ZN(new_n649));
  AOI211_X1 g0449(.A(new_n403), .B(new_n562), .C1(new_n259), .C2(new_n556), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n627), .A2(new_n585), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n621), .A2(new_n502), .A3(new_n487), .A4(new_n497), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n643), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n580), .A2(new_n585), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT26), .B1(new_n543), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n642), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n443), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n325), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n402), .A2(new_n410), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n411), .B(KEYINPUT17), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n663), .A2(new_n361), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n357), .A2(new_n440), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n660), .B1(new_n666), .B2(new_n319), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n659), .A2(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n498), .A2(new_n499), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n501), .A2(new_n478), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n487), .A2(new_n670), .A3(new_n671), .A4(new_n497), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n479), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n503), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT81), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n624), .A2(new_n619), .B1(new_n593), .B2(new_n597), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n678), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT82), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n678), .B1(new_n615), .B2(new_n620), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n621), .A2(new_n688), .A3(new_n627), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n672), .A2(new_n679), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n685), .B2(new_n679), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(KEYINPUT83), .ZN(new_n698));
  INV_X1    g0498(.A(new_n210), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(G41), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n210), .A2(KEYINPUT83), .A3(new_n261), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n569), .A2(G116), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n703), .A2(new_n206), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n214), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n703), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n592), .A2(new_n578), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n542), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT84), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n501), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n542), .A3(new_n711), .A4(new_n713), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n461), .A2(new_n323), .A3(new_n564), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n518), .A2(new_n521), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n596), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n678), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n629), .A2(new_n679), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n710), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT26), .B1(new_n636), .B2(new_n543), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n550), .B1(new_n321), .B2(new_n721), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n586), .A2(new_n730), .A3(new_n638), .A4(new_n522), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n585), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT85), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n648), .A2(new_n651), .B1(new_n641), .B2(new_n584), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n543), .A2(new_n734), .A3(new_n551), .A4(new_n627), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n732), .A2(new_n733), .B1(new_n654), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n729), .A2(new_n731), .A3(KEYINPUT85), .A4(new_n585), .ZN(new_n737));
  AOI211_X1 g0537(.A(KEYINPUT86), .B(new_n678), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT86), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n733), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n655), .A3(new_n737), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n741), .B2(new_n679), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT29), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n658), .A2(new_n679), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n728), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n709), .B1(new_n747), .B2(G1), .ZN(G364));
  AND2_X1   g0548(.A1(new_n207), .A2(G13), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n703), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n684), .B(new_n753), .C1(G330), .C2(new_n682), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n210), .A2(new_n255), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n210), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT87), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n245), .A2(G45), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT88), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n699), .A2(new_n255), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n215), .B2(new_n262), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n758), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n216), .B1(G20), .B2(new_n321), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n752), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n207), .A2(new_n323), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n275), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(KEYINPUT33), .A2(G317), .ZN(new_n776));
  AND2_X1   g0576(.A1(KEYINPUT33), .A2(G317), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n772), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n780), .A2(G311), .B1(G283), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n779), .A2(new_n403), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n403), .A2(new_n275), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n781), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n785), .A2(G322), .B1(G303), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n772), .A2(new_n786), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n255), .B1(new_n791), .B2(G326), .ZN(new_n792));
  AND4_X1   g0592(.A1(new_n778), .A2(new_n784), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n207), .ZN(new_n798));
  INV_X1    g0598(.A(G329), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(G20), .A3(new_n403), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT90), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n793), .B1(new_n794), .B2(new_n798), .C1(new_n799), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G159), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  INV_X1    g0608(.A(new_n780), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n809), .A2(new_n252), .B1(new_n202), .B2(new_n790), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G68), .B2(new_n775), .ZN(new_n811));
  INV_X1    g0611(.A(new_n798), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G97), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n782), .A2(new_n420), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n255), .B1(new_n787), .B2(new_n568), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G58), .C2(new_n785), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n811), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n805), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT91), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n768), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n771), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n767), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n682), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n754), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND3_X1  g0627(.A1(new_n438), .A2(KEYINPUT94), .A3(new_n439), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT94), .B1(new_n438), .B2(new_n439), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n829), .A2(new_n830), .A3(new_n436), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n734), .A2(new_n543), .A3(new_n551), .A4(new_n627), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n672), .A2(new_n685), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n734), .A2(new_n730), .A3(new_n638), .A4(new_n522), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n657), .A3(new_n585), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n679), .B(new_n831), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT95), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n658), .A2(KEYINPUT95), .A3(new_n679), .A4(new_n831), .ZN(new_n840));
  INV_X1    g0640(.A(new_n830), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n678), .B1(new_n429), .B2(new_n433), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(new_n437), .A3(new_n828), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n438), .A2(new_n439), .A3(new_n678), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n839), .A2(new_n840), .B1(new_n744), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n728), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT98), .Z(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n728), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT96), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT96), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n753), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n852), .B2(KEYINPUT97), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(KEYINPUT97), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n768), .A2(new_n765), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT92), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n752), .B1(G77), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G137), .A2(new_n791), .B1(new_n775), .B2(G150), .ZN(new_n858));
  INV_X1    g0658(.A(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G143), .ZN(new_n860));
  INV_X1    g0660(.A(new_n785), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n858), .B1(new_n809), .B2(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n255), .B1(new_n782), .B2(new_n331), .C1(new_n202), .C2(new_n787), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n812), .B2(G58), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n863), .B(new_n865), .C1(new_n866), .C2(new_n804), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n804), .A2(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n787), .A2(new_n420), .B1(new_n782), .B2(new_n568), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n374), .B1(new_n861), .B2(new_n794), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(G303), .C2(new_n791), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n780), .A2(G116), .B1(G283), .B2(new_n775), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT93), .Z(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n813), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n867), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n857), .B1(new_n876), .B2(new_n768), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n843), .A2(new_n844), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n766), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n854), .A2(new_n879), .ZN(G384));
  OR2_X1    g0680(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(G116), .A3(new_n217), .A4(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT36), .Z(new_n884));
  OR3_X1    g0684(.A1(new_n214), .A2(new_n252), .A3(new_n369), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n202), .A2(G68), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n206), .B(G13), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n385), .A2(new_n386), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n377), .A2(new_n378), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n304), .B1(new_n890), .B2(new_n363), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n891), .B2(new_n379), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n676), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n414), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n411), .B1(new_n892), .B2(new_n399), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT101), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n676), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n388), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n401), .A2(KEYINPUT101), .A3(new_n411), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n411), .C1(new_n892), .C2(new_n676), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n388), .A2(KEYINPUT99), .A3(new_n400), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT99), .B1(new_n388), .B2(new_n400), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n894), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT100), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n406), .A2(new_n408), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n903), .B1(new_n912), .B2(new_n899), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT99), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n401), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT37), .B1(new_n892), .B2(new_n405), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n408), .A2(KEYINPUT99), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n899), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n895), .B2(new_n893), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n909), .B1(new_n414), .B2(new_n893), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT102), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n919), .A2(KEYINPUT100), .A3(new_n920), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT100), .B1(new_n919), .B2(new_n920), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT102), .B(new_n923), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n910), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n337), .A2(new_n678), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n357), .A2(new_n361), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT14), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n353), .A3(new_n349), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n337), .B(new_n678), .C1(new_n934), .C2(new_n360), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n878), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n724), .A2(new_n725), .ZN(new_n939));
  INV_X1    g0739(.A(new_n503), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n628), .A2(new_n552), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n679), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n942), .A3(new_n727), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(KEYINPUT40), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n899), .B1(new_n661), .B2(new_n663), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n914), .B2(new_n921), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n946), .B1(new_n948), .B2(KEYINPUT38), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n937), .B1(new_n726), .B2(new_n727), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n929), .A2(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n953), .A2(new_n443), .A3(new_n943), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n443), .B2(new_n943), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n954), .A2(new_n955), .A3(new_n710), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n931), .A2(new_n935), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n839), .A2(new_n840), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n678), .B1(new_n841), .B2(new_n828), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n957), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n961), .A2(new_n949), .B1(new_n662), .B2(new_n676), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n894), .B1(new_n925), .B2(new_n926), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n909), .B1(new_n922), .B2(new_n923), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT39), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n934), .A2(new_n337), .A3(new_n679), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT102), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n946), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n969), .A2(new_n927), .B1(new_n909), .B2(new_n908), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n965), .B(new_n967), .C1(new_n970), .C2(KEYINPUT39), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n743), .A2(new_n443), .A3(new_n746), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n668), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n956), .A2(new_n975), .B1(new_n206), .B2(new_n749), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT103), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n956), .A2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n976), .A2(KEYINPUT103), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n888), .B1(new_n979), .B2(new_n980), .ZN(G367));
  NAND2_X1  g0781(.A1(new_n761), .A2(new_n237), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n770), .B1(new_n699), .B2(new_n582), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n753), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n734), .B1(new_n648), .B2(new_n679), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n634), .A2(new_n584), .A3(new_n641), .A4(new_n678), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G303), .ZN(new_n988));
  INV_X1    g0788(.A(G283), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n861), .A2(new_n988), .B1(new_n809), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT46), .B1(new_n788), .B2(G116), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT109), .Z(new_n992));
  NAND3_X1  g0792(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n374), .C1(new_n794), .C2(new_n774), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n790), .A2(new_n868), .B1(new_n782), .B2(new_n222), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n990), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n996), .B1(new_n420), .B2(new_n798), .C1(new_n997), .C2(new_n804), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n798), .A2(new_n331), .ZN(new_n999));
  INV_X1    g0799(.A(G150), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n861), .A2(new_n1000), .B1(new_n790), .B2(new_n860), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT110), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n806), .A2(G137), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n780), .A2(G50), .B1(G58), .B2(new_n788), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n859), .B2(new_n774), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n782), .A2(new_n252), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1007), .A2(new_n374), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT110), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1005), .B(new_n1009), .C1(new_n1010), .C2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n998), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n984), .B1(new_n824), .B2(new_n987), .C1(new_n1013), .C2(new_n821), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n643), .B1(new_n550), .B2(new_n679), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n543), .B2(new_n679), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n696), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT45), .Z(new_n1018));
  NOR2_X1   g0818(.A1(new_n696), .A2(new_n1016), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n692), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n690), .A2(new_n694), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT108), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n684), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1025), .B(new_n1027), .Z(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n747), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n747), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n702), .B(KEYINPUT41), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n751), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT105), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n1035));
  NAND3_X1  g0835(.A1(new_n985), .A2(new_n1035), .A3(new_n986), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(KEYINPUT106), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n695), .A2(new_n1016), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT42), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n543), .B1(new_n1015), .B2(new_n621), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n679), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n692), .A2(new_n1016), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1036), .A2(KEYINPUT106), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1044), .B(new_n1045), .Z(new_n1046));
  OAI21_X1  g0846(.A(new_n1014), .B1(new_n1032), .B2(new_n1046), .ZN(G387));
  NAND2_X1  g0847(.A1(new_n1028), .A2(new_n751), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n374), .B1(new_n782), .B2(new_n471), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G322), .A2(new_n791), .B1(new_n775), .B2(G311), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n809), .B2(new_n988), .C1(new_n997), .C2(new_n861), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1051), .A2(new_n1052), .B1(G294), .B2(new_n788), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .C1(new_n989), .C2(new_n798), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT49), .Z(new_n1055));
  AOI211_X1 g0855(.A(new_n1049), .B(new_n1055), .C1(G326), .C2(new_n806), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n812), .A2(new_n582), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n861), .A2(new_n202), .B1(new_n809), .B2(new_n331), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n790), .A2(new_n859), .B1(new_n787), .B2(new_n252), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n383), .A2(new_n775), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n374), .B1(new_n783), .B2(G97), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G150), .B2(new_n806), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n768), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n234), .A2(new_n262), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT111), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT111), .ZN(new_n1069));
  AOI211_X1 g0869(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n283), .A2(new_n202), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT50), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n762), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(KEYINPUT112), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(KEYINPUT112), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1068), .A2(new_n1069), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(G107), .B2(new_n210), .C1(new_n704), .C2(new_n755), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n753), .B1(new_n1078), .B2(new_n769), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1065), .B(new_n1079), .C1(new_n690), .C2(new_n824), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1048), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1029), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n702), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1028), .A2(new_n747), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G393));
  XNOR2_X1  g0886(.A(new_n1021), .B(new_n693), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n1082), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n1089), .A3(new_n703), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n751), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n242), .A2(new_n761), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n769), .B1(new_n222), .B2(new_n210), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n752), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n785), .A2(G159), .B1(new_n791), .B2(G150), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  OAI21_X1  g0896(.A(new_n255), .B1(new_n782), .B2(new_n568), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n202), .A2(new_n774), .B1(new_n787), .B2(new_n331), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n283), .C2(new_n780), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n252), .B2(new_n798), .C1(new_n860), .C2(new_n804), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n806), .A2(G322), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n785), .A2(G311), .B1(new_n791), .B2(G317), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT52), .Z(new_n1104));
  OAI22_X1  g0904(.A1(new_n809), .A2(new_n794), .B1(new_n989), .B2(new_n787), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1105), .A2(new_n255), .A3(new_n814), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n798), .A2(new_n471), .B1(new_n988), .B2(new_n774), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT113), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1101), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT114), .Z(new_n1111));
  AOI21_X1  g0911(.A(new_n1094), .B1(new_n1111), .B2(new_n768), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n824), .B2(new_n1016), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1090), .A2(new_n1091), .A3(new_n1113), .ZN(G390));
  NAND4_X1  g0914(.A1(new_n943), .A2(G330), .A3(new_n878), .A4(new_n936), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n878), .B1(new_n738), .B2(new_n742), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n957), .B1(new_n1117), .B2(new_n960), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n929), .A2(new_n966), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT39), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n929), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n958), .A2(new_n960), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n936), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1122), .A2(new_n965), .B1(new_n1124), .B2(new_n966), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1116), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n965), .B1(new_n970), .B2(KEYINPUT39), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n959), .B1(new_n839), .B2(new_n840), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n966), .B1(new_n1128), .B2(new_n957), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n1115), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n943), .A2(G330), .A3(new_n878), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n957), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1128), .B1(new_n1134), .B2(new_n1115), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n741), .A2(new_n679), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT86), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n741), .A2(new_n739), .A3(new_n679), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n959), .B1(new_n1139), .B2(new_n878), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1134), .A2(new_n1115), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1135), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n728), .A2(new_n443), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n973), .A2(new_n668), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1132), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1126), .A2(new_n1131), .A3(new_n1146), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n703), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1126), .A2(new_n751), .A3(new_n1131), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1127), .A2(new_n765), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n752), .B1(new_n383), .B2(new_n856), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n374), .B1(new_n780), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT53), .B1(new_n787), .B2(new_n1000), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n775), .A2(G137), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n861), .B2(new_n866), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n790), .A2(new_n1161), .B1(new_n782), .B2(new_n202), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n1000), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1158), .A2(new_n1160), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(G125), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n804), .C1(new_n859), .C2(new_n798), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n804), .A2(new_n794), .B1(new_n331), .B2(new_n782), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT117), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n785), .A2(G116), .B1(new_n791), .B2(G283), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n780), .A2(G97), .B1(G107), .B2(new_n775), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1171), .B2(KEYINPUT115), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G77), .B2(new_n812), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n374), .B1(new_n787), .B2(new_n568), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1171), .A2(KEYINPUT115), .B1(new_n1174), .B2(KEYINPUT116), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(KEYINPUT116), .C2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1166), .B1(new_n1168), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1153), .B1(new_n1177), .B2(new_n768), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1152), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1150), .A2(new_n1151), .A3(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1145), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1149), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n962), .A2(new_n971), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n315), .A2(new_n316), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n320), .A2(new_n676), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n660), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n319), .B2(new_n325), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n953), .B2(G330), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n969), .A2(new_n927), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n944), .B1(new_n1198), .B2(new_n910), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT40), .B1(new_n949), .B2(new_n950), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n1195), .A4(new_n710), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1184), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT120), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n953), .A2(G330), .A3(new_n1196), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n938), .A2(new_n943), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n952), .B1(new_n964), .B2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1206), .B(G330), .C1(new_n970), .C2(new_n944), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1195), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n972), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1203), .A3(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n972), .A2(new_n1204), .A3(new_n1208), .A4(KEYINPUT120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1181), .B1(new_n1183), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1149), .A2(new_n1182), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1181), .B1(new_n1202), .B2(new_n1209), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n702), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n752), .B1(G50), .B2(new_n856), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1196), .A2(new_n766), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n374), .A2(new_n261), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n782), .A2(new_n220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G77), .C2(new_n788), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n804), .B2(new_n989), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT118), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n785), .A2(G107), .B1(G97), .B2(new_n775), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n471), .B2(new_n790), .C1(new_n430), .C2(new_n809), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1224), .A2(new_n999), .A3(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT58), .Z(new_n1228));
  OAI211_X1 g1028(.A(new_n1220), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n785), .A2(G128), .B1(new_n788), .B2(new_n1155), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n790), .A2(new_n1165), .B1(new_n774), .B2(new_n866), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G137), .B2(new_n780), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(new_n798), .C2(new_n1000), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT119), .Z(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n463), .B(new_n261), .C1(new_n782), .C2(new_n859), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n806), .B2(G124), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT59), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1228), .B(new_n1229), .C1(new_n1236), .C2(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1218), .B(new_n1219), .C1(new_n768), .C2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n751), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1217), .A2(new_n1244), .ZN(G375));
  INV_X1    g1045(.A(new_n1143), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(KEYINPUT121), .A3(new_n751), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n752), .B1(G68), .B2(new_n856), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT122), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n785), .A2(G137), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n774), .B2(new_n1154), .C1(new_n809), .C2(new_n1000), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n790), .A2(new_n866), .B1(new_n787), .B2(new_n859), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1251), .A2(new_n374), .A3(new_n1252), .A4(new_n1221), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n202), .B2(new_n798), .C1(new_n804), .C2(new_n1161), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G107), .A2(new_n780), .B1(new_n785), .B2(G283), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n794), .B2(new_n790), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n222), .A2(new_n787), .B1(new_n774), .B2(new_n471), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1256), .A2(new_n255), .A3(new_n1257), .A4(new_n1008), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1258), .B(new_n1057), .C1(new_n988), .C2(new_n804), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1249), .B1(new_n821), .B2(new_n1260), .C1(new_n936), .C2(new_n766), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT121), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1143), .B2(new_n750), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1247), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1246), .A2(new_n1182), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1031), .A3(new_n1147), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(G381));
  NOR3_X1   g1069(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G375), .A2(G378), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1085), .A2(new_n826), .A3(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT123), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1271), .A3(new_n1274), .ZN(G407));
  NAND2_X1  g1075(.A1(new_n677), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1271), .A2(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT124), .Z(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(G213), .A3(G407), .ZN(G409));
  NAND4_X1  g1080(.A1(new_n1243), .A2(KEYINPUT125), .A3(new_n1031), .A4(new_n1214), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1210), .A2(new_n1031), .A3(new_n1211), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1183), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1202), .A2(new_n1209), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1242), .B1(new_n1285), .B2(new_n751), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1281), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  INV_X1    g1088(.A(G378), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1217), .A2(G378), .A3(new_n1244), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1288), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1276), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1277), .A2(G2897), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1266), .B1(KEYINPUT60), .B2(new_n1147), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1143), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n703), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1265), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1272), .A2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G384), .B(new_n1265), .C1(new_n1296), .C2(new_n1298), .ZN(new_n1301));
  AOI211_X1 g1101(.A(KEYINPUT127), .B(new_n1295), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G2897), .B(new_n1277), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1293), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n1291), .A3(new_n1290), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1303), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1276), .A4(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1276), .B(new_n1312), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT62), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1308), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(G390), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G387), .A2(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G390), .B(new_n1014), .C1(new_n1032), .C2(new_n1046), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1085), .B(G396), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1320), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1316), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1314), .A2(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1276), .A4(new_n1312), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1308), .A2(new_n1323), .A3(new_n1327), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1325), .A2(new_n1329), .ZN(G405));
  XNOR2_X1  g1130(.A(G375), .B(new_n1289), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1303), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1323), .ZN(G402));
endmodule


