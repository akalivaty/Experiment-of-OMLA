//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  OR3_X1    g0004(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT64), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G50), .B2(G226), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G97), .A2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G77), .A2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n224), .A2(new_n225), .B1(new_n206), .B2(new_n205), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n204), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n217), .A2(new_n212), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n210), .B(new_n227), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(G250), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(KEYINPUT68), .B(G107), .ZN(new_n244));
  INV_X1    g0044(.A(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT13), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI211_X1 g0060(.A(G232), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n268), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1698), .B1(new_n266), .B2(new_n267), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n271), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n258), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n277), .B(new_n203), .C1(G41), .C2(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G238), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n255), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(G1), .B(G13), .C1(new_n265), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n270), .B2(new_n272), .ZN(new_n284));
  INV_X1    g0084(.A(new_n280), .ZN(new_n285));
  NOR4_X1   g0085(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT13), .A4(new_n258), .ZN(new_n286));
  OAI21_X1  g0086(.A(G169), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n273), .A2(new_n274), .ZN(new_n289));
  INV_X1    g0089(.A(new_n258), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(new_n280), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n275), .A2(new_n255), .A3(new_n280), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G179), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(G169), .C1(new_n281), .C2(new_n286), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n288), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT74), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n204), .A2(G68), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n265), .A2(new_n300), .A3(G20), .ZN(new_n301));
  NOR3_X1   g0101(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI211_X1 g0105(.A(new_n299), .B(new_n301), .C1(new_n305), .C2(G50), .ZN(new_n306));
  NAND3_X1  g0106(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n228), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT11), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  INV_X1    g0111(.A(new_n304), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(new_n302), .ZN(new_n313));
  INV_X1    g0113(.A(G50), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n204), .B2(G68), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n311), .B(new_n308), .C1(new_n315), .C2(new_n301), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n203), .A2(G20), .ZN(new_n318));
  INV_X1    g0118(.A(G13), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OR3_X1    g0121(.A1(new_n321), .A2(KEYINPUT12), .A3(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT12), .B1(new_n321), .B2(G68), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n308), .B1(new_n203), .B2(G20), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(new_n323), .B1(G68), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n317), .A2(KEYINPUT73), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT73), .B1(new_n317), .B2(new_n325), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n298), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n317), .A2(new_n325), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n317), .A2(KEYINPUT73), .A3(new_n325), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(KEYINPUT74), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n297), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n292), .A2(new_n293), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n332), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n292), .A2(G190), .A3(new_n293), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT72), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n341), .A3(G200), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(new_n339), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT75), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G222), .ZN(new_n348));
  INV_X1    g0148(.A(G223), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n268), .B(new_n348), .C1(new_n349), .C2(new_n347), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n274), .C1(G77), .C2(new_n268), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n279), .A2(G226), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n290), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT8), .B(G58), .Z(new_n355));
  NOR2_X1   g0155(.A1(new_n265), .A2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n313), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n308), .B1(new_n314), .B2(new_n320), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n324), .A2(G50), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n353), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n354), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT9), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n363), .A2(new_n368), .B1(G200), .B2(new_n353), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n369), .B1(new_n368), .B2(new_n363), .C1(new_n370), .C2(new_n353), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G238), .A2(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n268), .B(new_n375), .C1(new_n218), .C2(G1698), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n274), .C1(G107), .C2(new_n268), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n290), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(G244), .B2(new_n279), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(G169), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT15), .B(G87), .Z(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n356), .B1(G20), .B2(G77), .ZN(new_n382));
  INV_X1    g0182(.A(new_n355), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n313), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n308), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n324), .A2(G77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n320), .A2(new_n300), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n380), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n379), .B2(G190), .ZN(new_n392));
  INV_X1    g0192(.A(G200), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n379), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n355), .A2(new_n318), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT79), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n320), .A2(new_n308), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n397), .A2(new_n398), .B1(new_n320), .B2(new_n383), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n259), .A2(new_n260), .ZN(new_n401));
  AND2_X1   g0201(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n404), .A3(new_n204), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n266), .A2(new_n204), .A3(new_n267), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT76), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n410), .A3(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(G68), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(G58), .B(G68), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n305), .A2(G159), .B1(new_n413), .B2(G20), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(new_n308), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT78), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n267), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n259), .A2(new_n260), .A3(G20), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n418), .C1(new_n419), .C2(new_n404), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(KEYINPUT78), .A3(KEYINPUT7), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G68), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n414), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n400), .B1(new_n416), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n349), .A2(new_n347), .ZN(new_n427));
  INV_X1    g0227(.A(G226), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n429), .C1(new_n259), .C2(new_n260), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n283), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n258), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n279), .A2(G232), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(G190), .A3(new_n434), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n425), .A2(new_n308), .A3(new_n415), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(new_n436), .A3(new_n437), .A4(new_n399), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n415), .A2(new_n308), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT16), .B1(new_n422), .B2(new_n414), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n399), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n433), .A2(G179), .A3(new_n434), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n364), .B1(new_n433), .B2(new_n434), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT18), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  AOI211_X1 g0251(.A(new_n451), .B(new_n448), .C1(new_n439), .C2(new_n399), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n438), .B(new_n442), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n453), .A2(new_n454), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n374), .B(new_n395), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n346), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n204), .A2(G107), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT23), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  AOI21_X1  g0262(.A(G20), .B1(new_n266), .B2(new_n267), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G87), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n204), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT22), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n459), .B(new_n461), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n465), .B(KEYINPUT22), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(KEYINPUT24), .A3(new_n459), .A4(new_n461), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n471), .A3(new_n308), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT87), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(KEYINPUT25), .C1(new_n321), .C2(G107), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n265), .A2(G1), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n320), .A2(new_n308), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G107), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G107), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n473), .A2(KEYINPUT25), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(KEYINPUT25), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n320), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n222), .A2(new_n347), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n268), .B(new_n483), .C1(G257), .C2(new_n347), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G294), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  INV_X1    g0287(.A(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G1), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n274), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n486), .A2(new_n274), .B1(G264), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n203), .A2(G45), .A3(G274), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n496), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n487), .A2(new_n498), .A3(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n393), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G190), .B2(new_n501), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n478), .A2(new_n482), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT88), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n472), .A2(new_n482), .A3(new_n474), .A4(new_n477), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n491), .A2(new_n389), .A3(new_n500), .ZN(new_n507));
  AOI21_X1  g0307(.A(G169), .B1(new_n491), .B2(new_n500), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n505), .B1(new_n504), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n321), .A2(G116), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n476), .B2(G116), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n245), .A2(G20), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n308), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n204), .B1(new_n522), .B2(G33), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT85), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT85), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(new_n265), .B2(G97), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n524), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n521), .B(KEYINPUT20), .C1(new_n526), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT86), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n521), .B1(new_n526), .B2(new_n529), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT85), .B1(new_n523), .B2(new_n525), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n528), .A2(new_n527), .A3(new_n524), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n520), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT86), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT20), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n518), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n347), .A2(G257), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G264), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n259), .C2(new_n260), .ZN(new_n545));
  INV_X1    g0345(.A(G303), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n266), .A2(new_n546), .A3(new_n267), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n274), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n490), .A2(G270), .B1(new_n497), .B2(new_n499), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n364), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n515), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n539), .B1(new_n538), .B2(KEYINPUT20), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n538), .A2(KEYINPUT20), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n517), .B1(new_n559), .B2(new_n540), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT21), .A3(new_n554), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n552), .A2(new_n553), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n389), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n535), .A2(new_n541), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n552), .A2(new_n553), .A3(G190), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n517), .A4(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n556), .A2(new_n561), .A3(new_n564), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n420), .A2(G107), .A3(new_n421), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n305), .A2(G77), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n479), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n522), .A2(new_n479), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n575), .B2(KEYINPUT6), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n570), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n308), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n321), .A2(G97), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n476), .B2(G97), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  INV_X1    g0383(.A(G244), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n401), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n347), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n524), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n268), .A2(G250), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n347), .B1(new_n588), .B2(KEYINPUT4), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n274), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G257), .A3(new_n283), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n495), .A2(new_n492), .A3(new_n496), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT81), .B1(new_n487), .B2(new_n498), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n364), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT82), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n500), .A2(new_n600), .A3(new_n592), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n590), .A2(new_n599), .A3(new_n389), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n582), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n590), .A2(new_n599), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  INV_X1    g0405(.A(new_n581), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n578), .B2(new_n308), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n590), .A2(G190), .A3(new_n596), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n221), .A2(new_n522), .A3(new_n479), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G97), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n204), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT19), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n204), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n612), .A2(G20), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(KEYINPUT19), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n381), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n308), .B1(new_n320), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n476), .A2(new_n381), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT83), .ZN(new_n622));
  NOR2_X1   g0422(.A1(G238), .A2(G1698), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n268), .B(new_n624), .C1(G244), .C2(new_n347), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G116), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n283), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G250), .B1(new_n488), .B2(G1), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n274), .B1(new_n496), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n364), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT83), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n619), .A2(new_n631), .A3(new_n620), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n259), .A2(new_n260), .B1(G244), .B2(new_n347), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n626), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n629), .B1(new_n634), .B2(new_n274), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n389), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n622), .A2(new_n630), .A3(new_n632), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n476), .A2(G87), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n635), .A2(G190), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n639), .B(new_n640), .C1(new_n393), .C2(new_n635), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n569), .A2(new_n610), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n458), .A2(new_n514), .A3(new_n643), .ZN(G372));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n635), .B2(new_n393), .ZN(new_n647));
  OAI211_X1 g0447(.A(KEYINPUT90), .B(G200), .C1(new_n627), .C2(new_n629), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n639), .A2(new_n647), .A3(new_n648), .A4(new_n640), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT89), .B1(new_n635), .B2(G169), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(new_n364), .C1(new_n627), .C2(new_n629), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n650), .A2(new_n621), .A3(new_n652), .A4(new_n636), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n645), .B1(new_n603), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT91), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n637), .A2(new_n641), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n582), .A2(new_n602), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n598), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n660), .B(new_n645), .C1(new_n603), .C2(new_n654), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n656), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n510), .A2(new_n556), .A3(new_n561), .A4(new_n564), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n603), .A2(new_n609), .A3(new_n649), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n504), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n653), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n458), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n452), .A2(new_n450), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n391), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n343), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n335), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n438), .A2(new_n442), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n371), .B(KEYINPUT10), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n367), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n556), .A2(new_n561), .A3(new_n564), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n319), .A2(G20), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n203), .ZN(new_n680));
  XNOR2_X1  g0480(.A(KEYINPUT92), .B(KEYINPUT27), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n542), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT93), .B1(new_n569), .B2(new_n688), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT94), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n691), .B(new_n695), .C1(new_n689), .C2(new_n692), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G330), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n510), .A2(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n506), .A2(new_n686), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n514), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n678), .A2(new_n687), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n513), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n510), .A2(new_n686), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n208), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n611), .A2(G116), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n709), .A2(new_n203), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT95), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT95), .ZN(new_n714));
  INV_X1    g0514(.A(new_n709), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n713), .B(new_n714), .C1(new_n231), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT97), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n666), .A2(new_n719), .A3(new_n687), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(new_n666), .B2(new_n687), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n658), .A2(new_n598), .A3(new_n649), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT26), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n657), .A2(new_n645), .A3(new_n598), .A4(new_n658), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n665), .A2(new_n653), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n687), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n643), .B(new_n687), .C1(new_n511), .C2(new_n512), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n590), .A2(new_n596), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT96), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n491), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n563), .A2(new_n732), .A3(new_n736), .A4(new_n635), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n733), .A2(new_n734), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n501), .B1(new_n627), .B2(new_n629), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n604), .A2(new_n389), .A3(new_n562), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n686), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n745), .A3(new_n686), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(G330), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n730), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n717), .B1(new_n749), .B2(G1), .ZN(G364));
  AOI21_X1  g0550(.A(new_n228), .B1(G20), .B2(new_n364), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT99), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT99), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n204), .A2(new_n370), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n389), .A2(new_n393), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n204), .B1(new_n760), .B2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(G294), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT102), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n204), .A2(G190), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT101), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT101), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n766), .A2(new_n767), .A3(new_n760), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n268), .B1(new_n768), .B2(G329), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(new_n765), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G317), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT33), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(KEYINPUT33), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n389), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n765), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n769), .B(new_n775), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n756), .A2(new_n777), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n764), .B(new_n779), .C1(G322), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n393), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n766), .A2(new_n784), .A3(new_n767), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n756), .A2(new_n784), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n782), .B1(new_n783), .B2(new_n785), .C1(new_n546), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT103), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n768), .A2(G159), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT32), .Z(new_n790));
  OAI22_X1  g0590(.A1(new_n780), .A2(new_n217), .B1(new_n778), .B2(new_n300), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT100), .Z(new_n792));
  INV_X1    g0592(.A(new_n785), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G107), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n758), .A2(new_n314), .B1(new_n770), .B2(new_n212), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n786), .A2(new_n221), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n761), .A2(new_n522), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n401), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n790), .A2(new_n792), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n755), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n754), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n208), .A2(G355), .A3(new_n268), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n253), .A2(G45), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n708), .A2(new_n268), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(G45), .B2(new_n232), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n805), .B1(G116), .B2(new_n208), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n800), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n203), .B1(new_n679), .B2(G45), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n709), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n694), .A2(new_n696), .ZN(new_n815));
  INV_X1    g0615(.A(new_n803), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n811), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n814), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n697), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(G330), .B2(new_n815), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  AND3_X1   g0622(.A1(new_n656), .A2(new_n659), .A3(new_n661), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n665), .A2(new_n653), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n687), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT97), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n388), .A2(new_n686), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n394), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n391), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n670), .A2(new_n687), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n826), .A2(new_n720), .A3(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n687), .B(new_n831), .C1(new_n823), .C2(new_n824), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n748), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n747), .A3(new_n834), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n818), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n786), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n793), .A2(G68), .B1(G50), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(KEYINPUT105), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n758), .A2(new_n842), .B1(new_n770), .B2(new_n359), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT104), .ZN(new_n844));
  INV_X1    g0644(.A(G143), .ZN(new_n845));
  INV_X1    g0645(.A(G159), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(new_n845), .B2(new_n780), .C1(new_n846), .C2(new_n778), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  INV_X1    g0648(.A(new_n761), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n840), .A2(KEYINPUT105), .B1(G58), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n268), .A3(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n841), .B(new_n851), .C1(G132), .C2(new_n768), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n778), .A2(new_n245), .B1(new_n761), .B2(new_n522), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n758), .A2(new_n546), .B1(new_n770), .B2(new_n783), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n768), .C2(G311), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n268), .B1(new_n839), .B2(G107), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(new_n762), .C2(new_n780), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G87), .B2(new_n793), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n754), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n754), .A2(new_n801), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n859), .B1(G77), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n801), .B2(new_n832), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n838), .B1(new_n818), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT106), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n864), .B(new_n865), .ZN(G384));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(new_n684), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n453), .A2(new_n445), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n448), .A2(new_n684), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n445), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n440), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(new_n874), .A3(new_n440), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(KEYINPUT109), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT109), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n867), .B1(new_n869), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT16), .B1(new_n412), .B2(new_n414), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n399), .B1(new_n443), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n868), .B(new_n882), .C1(new_n673), .C2(new_n668), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n870), .ZN(new_n884));
  INV_X1    g0684(.A(new_n440), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n875), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n334), .A2(new_n686), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT108), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n297), .A2(new_n334), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n297), .B2(new_n334), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n343), .B(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n344), .A2(new_n334), .A3(new_n686), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n832), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT110), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n744), .A2(new_n897), .A3(new_n746), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n744), .B2(new_n746), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n889), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n883), .B2(new_n887), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT40), .B1(new_n903), .B2(new_n888), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n458), .B1(new_n898), .B2(new_n899), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(G330), .ZN(new_n909));
  INV_X1    g0709(.A(new_n676), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n730), .B2(new_n458), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n894), .A2(new_n895), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n888), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT107), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n834), .A2(new_n914), .A3(new_n830), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n834), .B2(new_n830), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n912), .B(new_n913), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n876), .A2(new_n878), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n453), .A2(new_n445), .A3(new_n868), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n892), .A2(new_n893), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n686), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n669), .A2(new_n868), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n917), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n911), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n909), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n203), .B2(new_n679), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n245), .B1(new_n576), .B2(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n229), .C1(KEYINPUT35), .C2(new_n576), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  OAI21_X1  g0736(.A(G77), .B1(new_n217), .B2(new_n212), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n231), .A2(new_n937), .B1(G50), .B2(new_n212), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G1), .A3(new_n319), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n936), .A3(new_n939), .ZN(G367));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n603), .B(new_n609), .C1(new_n607), .C2(new_n687), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n658), .A2(new_n598), .A3(new_n686), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n704), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT111), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n609), .A2(new_n506), .A3(new_n509), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n686), .B1(new_n947), .B2(new_n603), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n704), .A2(new_n941), .A3(new_n944), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n639), .A2(new_n687), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n653), .A3(new_n649), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n653), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n952), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n949), .A2(new_n950), .A3(new_n957), .A4(new_n951), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n944), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n702), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n966), .B(new_n960), .C1(new_n962), .C2(new_n963), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n709), .B(KEYINPUT41), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT45), .B1(new_n706), .B2(new_n944), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  NOR4_X1   g0773(.A1(new_n704), .A2(new_n973), .A3(new_n705), .A4(new_n965), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT44), .B1(new_n706), .B2(new_n944), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n977), .B(new_n965), .C1(new_n704), .C2(new_n705), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n975), .A2(new_n702), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n972), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n976), .A2(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n701), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n699), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n703), .B1(new_n510), .B2(new_n687), .C1(new_n513), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n513), .B2(new_n703), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n986), .A2(new_n815), .A3(KEYINPUT113), .A4(G330), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT113), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n697), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n694), .A2(KEYINPUT113), .A3(G330), .A4(new_n696), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n987), .B1(new_n991), .B2(new_n986), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n749), .A2(new_n992), .A3(KEYINPUT114), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT114), .B1(new_n749), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n983), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n971), .B1(new_n995), .B2(new_n749), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n968), .B(new_n969), .C1(new_n996), .C2(new_n813), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n268), .B1(new_n785), .B2(new_n300), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G58), .A2(new_n839), .B1(new_n771), .B2(G159), .ZN(new_n999));
  INV_X1    g0799(.A(new_n768), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n842), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n778), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n998), .B(new_n1001), .C1(G50), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n761), .A2(new_n212), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G150), .B2(new_n781), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT116), .Z(new_n1006));
  OAI211_X1 g0806(.A(new_n1003), .B(new_n1006), .C1(new_n845), .C2(new_n758), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n778), .A2(new_n783), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n786), .A2(new_n245), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n401), .B1(new_n479), .B2(new_n761), .C1(new_n1009), .C2(KEYINPUT46), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT46), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n758), .A2(new_n776), .B1(new_n780), .B2(new_n546), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT115), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1010), .B(new_n1014), .C1(G97), .C2(new_n793), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n768), .A2(G317), .B1(G294), .B2(new_n771), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1007), .B1(new_n1008), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT117), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n754), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n956), .A2(new_n816), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n808), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n804), .B1(new_n208), .B2(new_n618), .C1(new_n1024), .C2(new_n242), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n814), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n997), .A2(new_n1026), .ZN(G387));
  NOR3_X1   g0827(.A1(new_n238), .A2(new_n488), .A3(new_n268), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n383), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT50), .B1(new_n383), .B2(G50), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(G68), .A2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n488), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n711), .B1(new_n1032), .B2(new_n401), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n208), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1034), .B(new_n804), .C1(new_n479), .C2(new_n208), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT118), .B(G150), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n768), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n849), .A2(new_n381), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n522), .C2(new_n785), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n401), .B1(new_n1002), .B2(G68), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n300), .B2(new_n786), .C1(new_n846), .C2(new_n758), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n383), .A2(new_n770), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n780), .A2(new_n314), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n758), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G322), .A2(new_n1045), .B1(new_n771), .B2(G311), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n546), .B2(new_n778), .C1(new_n772), .C2(new_n780), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT48), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n783), .B2(new_n761), .C1(new_n762), .C2(new_n786), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT49), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n401), .B1(new_n1000), .B2(new_n759), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G116), .B2(new_n793), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1044), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n814), .B(new_n1035), .C1(new_n1053), .C2(new_n755), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n700), .B2(new_n803), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n992), .B2(new_n813), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n749), .A2(new_n992), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n709), .B1(new_n749), .B2(new_n992), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n983), .A2(new_n813), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n249), .A2(new_n808), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n803), .B(new_n754), .C1(new_n708), .C2(G97), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n818), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n768), .A2(G322), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n794), .B(new_n1065), .C1(new_n783), .C2(new_n786), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n268), .B(new_n1066), .C1(G303), .C2(new_n771), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G317), .A2(new_n1045), .B1(new_n781), .B2(G311), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1068), .A2(KEYINPUT52), .B1(G116), .B2(new_n849), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(KEYINPUT52), .B2(new_n1068), .C1(new_n762), .C2(new_n778), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n768), .A2(G143), .B1(G68), .B2(new_n839), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT119), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n268), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n383), .A2(new_n778), .B1(new_n300), .B2(new_n761), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1072), .A2(new_n1073), .B1(G87), .B2(new_n793), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n771), .A2(G50), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n758), .A2(new_n359), .B1(new_n780), .B2(new_n846), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1071), .A2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1064), .B1(new_n816), .B2(new_n944), .C1(new_n1082), .C2(new_n755), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1061), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n995), .B1(new_n983), .B2(new_n1058), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n715), .ZN(G390));
  AOI21_X1  g0887(.A(KEYINPUT39), .B1(new_n880), .B2(new_n888), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n922), .A2(new_n902), .A3(new_n918), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1090), .A2(new_n802), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1000), .A2(new_n762), .B1(new_n212), .B2(new_n785), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n761), .A2(new_n300), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n401), .B1(new_n770), .B2(new_n479), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n758), .A2(new_n783), .B1(new_n786), .B2(new_n221), .ZN(new_n1095));
  NOR4_X1   g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n522), .B2(new_n778), .C1(new_n245), .C2(new_n780), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n268), .B1(new_n778), .B2(new_n1099), .C1(new_n785), .C2(new_n314), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G125), .B2(new_n768), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n781), .A2(G132), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n839), .A2(new_n1036), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT53), .Z(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n758), .A2(new_n1105), .B1(new_n770), .B2(new_n842), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G159), .B2(new_n849), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n755), .B1(new_n1097), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n814), .B1(new_n355), .B2(new_n861), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1091), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(G330), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n925), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1113), .A2(new_n1114), .B1(new_n923), .B2(new_n926), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n727), .A2(new_n687), .A3(new_n829), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n830), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT120), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT120), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1119), .A3(new_n830), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n912), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n925), .B1(new_n888), .B2(new_n880), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1112), .B1(new_n1115), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n923), .A2(new_n926), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n894), .A2(new_n895), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n834), .A2(new_n830), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT107), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n834), .A2(new_n914), .A3(new_n830), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1125), .B1(new_n1130), .B2(new_n925), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n744), .A2(G330), .A3(new_n746), .A4(new_n831), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(new_n1126), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1111), .B1(new_n1136), .B2(new_n813), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT29), .B1(new_n826), .B2(new_n720), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n729), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n458), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n458), .B(G330), .C1(new_n898), .C2(new_n899), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n676), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1133), .A2(new_n1126), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1112), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n915), .A2(new_n916), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n831), .C1(new_n898), .C2(new_n899), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1126), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1120), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1119), .B1(new_n1116), .B2(new_n830), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1150), .A2(new_n1151), .B1(new_n1133), .B2(new_n1126), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1142), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n709), .B1(new_n1136), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1152), .B1(new_n1126), .B2(new_n1148), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1145), .B1(new_n1112), .B2(new_n1143), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n911), .B(new_n1141), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1124), .B2(new_n1135), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1137), .B1(new_n1156), .B2(new_n1160), .ZN(G378));
  AND3_X1   g0961(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1112), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1155), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1142), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(G330), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n901), .B2(new_n905), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n374), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n374), .A2(new_n1171), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n363), .A2(new_n868), .ZN(new_n1174));
  OR3_X1    g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n930), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n917), .A2(new_n927), .A3(new_n929), .A4(new_n1177), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1169), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1169), .B1(new_n1180), .B2(new_n1179), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1167), .A2(KEYINPUT57), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1142), .B1(new_n1136), .B2(new_n1155), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n906), .A2(G330), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n928), .B1(new_n1090), .B2(new_n925), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1177), .B1(new_n1188), .B2(new_n917), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1180), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1169), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1185), .B1(new_n1186), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1184), .A2(new_n1194), .A3(new_n709), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G50), .B1(new_n267), .B2(new_n282), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n785), .A2(new_n217), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G41), .B1(new_n768), .B2(G283), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n522), .B2(new_n770), .C1(new_n245), .C2(new_n758), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(G107), .C2(new_n781), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n268), .B(new_n1004), .C1(new_n381), .C2(new_n1002), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n300), .C2(new_n786), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT121), .Z(new_n1205));
  NAND2_X1  g1005(.A1(new_n771), .A2(G132), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G128), .A2(new_n781), .B1(new_n1002), .B2(G137), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1045), .A2(G125), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n839), .A2(new_n1098), .B1(new_n849), .B2(G150), .ZN(new_n1209));
  AND4_X1   g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT59), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(G33), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G41), .B1(new_n768), .B2(G124), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n846), .C2(new_n785), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1202), .A2(new_n1203), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n754), .B1(new_n1205), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT122), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1177), .A2(new_n801), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1218), .A2(new_n814), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(G50), .B2(new_n861), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1193), .B2(new_n812), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1195), .A2(new_n1223), .ZN(G375));
  NOR2_X1   g1024(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT123), .B1(new_n1225), .B2(new_n812), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1126), .A2(new_n801), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n860), .A2(new_n212), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n758), .A2(new_n762), .B1(new_n778), .B2(new_n479), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G116), .B2(new_n771), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT124), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G303), .B2(new_n768), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n793), .A2(G77), .B1(G283), .B2(new_n781), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1038), .A3(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n268), .B(new_n1234), .C1(G97), .C2(new_n839), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1197), .B1(G132), .B2(new_n1045), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n1105), .B2(new_n1000), .C1(new_n846), .C2(new_n786), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n780), .A2(new_n842), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1099), .A2(new_n770), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n268), .B1(new_n761), .B2(new_n314), .C1(new_n359), .C2(new_n778), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n754), .B1(new_n1235), .B2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1227), .A2(new_n814), .A3(new_n1228), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n813), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1226), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1225), .A2(new_n1142), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n970), .A3(new_n1159), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(G381));
  NOR2_X1   g1049(.A1(G375), .A2(G378), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n979), .A2(new_n982), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT114), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1057), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n749), .A2(new_n992), .A3(KEYINPUT114), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n983), .A2(new_n1058), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1084), .B1(new_n1258), .B2(new_n709), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n997), .A2(new_n1026), .A3(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1260), .A2(G384), .A3(G381), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1251), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1263), .B2(new_n1262), .ZN(G407));
  NAND2_X1  g1065(.A1(new_n685), .A2(G213), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT126), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1250), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT127), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1268), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1269), .A4(new_n1270), .ZN(G409));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1195), .B2(new_n1223), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1186), .A2(new_n1193), .A3(new_n971), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1274), .A2(G378), .A3(new_n1222), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1273), .A2(new_n1267), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1247), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1147), .A2(new_n1154), .A3(KEYINPUT60), .A4(new_n1142), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n709), .A3(new_n1159), .A4(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(new_n1246), .A3(G384), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n864), .B(KEYINPUT106), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1159), .A3(new_n709), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT60), .B1(new_n1225), .B2(new_n1142), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1226), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1281), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1276), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1267), .A2(G2897), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1281), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1267), .B1(G375), .B2(G378), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1275), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1290), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(G393), .B(new_n821), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n968), .A2(new_n969), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n749), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n970), .B1(new_n1256), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1302), .B1(new_n1304), .B2(new_n812), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1026), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1305), .A2(G390), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1259), .B1(new_n997), .B2(new_n1026), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1301), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(G390), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1301), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1260), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  NOR4_X1   g1113(.A1(new_n1273), .A2(new_n1267), .A3(new_n1275), .A4(new_n1288), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(KEYINPUT63), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1300), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  OAI22_X1  g1118(.A1(new_n1314), .A2(new_n1318), .B1(new_n1276), .B2(new_n1295), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1296), .A2(new_n1318), .A3(new_n1289), .A4(new_n1297), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1316), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1313), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1322), .ZN(G405));
  NOR2_X1   g1123(.A1(new_n1250), .A2(new_n1273), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1313), .A2(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1309), .B(new_n1312), .C1(new_n1250), .C2(new_n1273), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1325), .A2(new_n1289), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1289), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


