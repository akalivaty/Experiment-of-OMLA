

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XNOR2_X1 U322 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U323 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U324 ( .A(n302), .B(n301), .ZN(n290) );
  XOR2_X1 U325 ( .A(G15GAT), .B(G113GAT), .Z(n291) );
  NOR2_X1 U326 ( .A1(n457), .A2(n462), .ZN(n458) );
  INV_X1 U327 ( .A(KEYINPUT20), .ZN(n296) );
  XNOR2_X1 U328 ( .A(n297), .B(n296), .ZN(n298) );
  INV_X1 U329 ( .A(KEYINPUT55), .ZN(n445) );
  XNOR2_X1 U330 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U331 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U332 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n450) );
  XOR2_X1 U334 ( .A(n290), .B(n320), .Z(n525) );
  XNOR2_X1 U335 ( .A(n472), .B(n471), .ZN(n496) );
  XNOR2_X1 U336 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U337 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(G190GAT), .B(G134GAT), .Z(n383) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(G43GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n291), .B(n292), .ZN(n354) );
  XOR2_X1 U341 ( .A(n383), .B(n354), .Z(n294) );
  NAND2_X1 U342 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U344 ( .A(G99GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n295), .B(G120GAT), .ZN(n363) );
  XNOR2_X1 U346 ( .A(n363), .B(KEYINPUT81), .ZN(n297) );
  XOR2_X1 U347 ( .A(n300), .B(KEYINPUT82), .Z(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT0), .B(G127GAT), .Z(n423) );
  XNOR2_X1 U349 ( .A(n423), .B(KEYINPUT84), .ZN(n301) );
  XOR2_X1 U350 ( .A(G176GAT), .B(KEYINPUT83), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n305) );
  XOR2_X1 U354 ( .A(n306), .B(n305), .Z(n320) );
  XOR2_X1 U355 ( .A(G92GAT), .B(G204GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(G36GAT), .B(G190GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U358 ( .A(KEYINPUT97), .B(n309), .Z(n311) );
  NAND2_X1 U359 ( .A1(G226GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U361 ( .A(G64GAT), .B(KEYINPUT98), .Z(n313) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G8GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(n315), .B(n314), .Z(n322) );
  XNOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n316), .B(KEYINPUT21), .ZN(n317) );
  XOR2_X1 U367 ( .A(n317), .B(KEYINPUT89), .Z(n319) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(G218GAT), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n442) );
  XNOR2_X1 U370 ( .A(n320), .B(n442), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n513) );
  XOR2_X1 U372 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n332) );
  NAND2_X1 U375 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XOR2_X1 U376 ( .A(G78GAT), .B(G155GAT), .Z(n326) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(G71GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U379 ( .A(G22GAT), .B(G211GAT), .Z(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n340) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(G8GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n333), .B(KEYINPUT69), .ZN(n353) );
  XOR2_X1 U385 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n335) );
  XNOR2_X1 U386 ( .A(G183GAT), .B(G127GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n353), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(G57GAT), .B(G64GAT), .Z(n337) );
  XOR2_X1 U390 ( .A(KEYINPUT13), .B(n337), .Z(n371) );
  XOR2_X1 U391 ( .A(n338), .B(n371), .Z(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n560) );
  XOR2_X1 U393 ( .A(KEYINPUT7), .B(G50GAT), .Z(n342) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(n343), .Z(n392) );
  XOR2_X1 U397 ( .A(G141GAT), .B(G22GAT), .Z(n433) );
  XOR2_X1 U398 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n345) );
  XNOR2_X1 U399 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U401 ( .A(n433), .B(n346), .Z(n348) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n350) );
  XNOR2_X1 U405 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n352), .B(n351), .Z(n356) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U410 ( .A(n392), .B(n357), .Z(n566) );
  INV_X1 U411 ( .A(n566), .ZN(n542) );
  XNOR2_X1 U412 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n372) );
  XOR2_X1 U413 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n359) );
  NAND2_X1 U414 ( .A1(G230GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U416 ( .A(n360), .B(KEYINPUT32), .Z(n365) );
  XOR2_X1 U417 ( .A(G78GAT), .B(G148GAT), .Z(n362) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G204GAT), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n436) );
  XNOR2_X1 U420 ( .A(n363), .B(n436), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U422 ( .A(G85GAT), .B(G92GAT), .Z(n384) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(n384), .ZN(n367) );
  INV_X1 U424 ( .A(KEYINPUT73), .ZN(n366) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n571) );
  XNOR2_X1 U426 ( .A(n372), .B(n571), .ZN(n556) );
  AND2_X1 U427 ( .A1(n542), .A2(n556), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n373), .B(KEYINPUT46), .ZN(n374) );
  NOR2_X1 U429 ( .A1(n560), .A2(n374), .ZN(n395) );
  XOR2_X1 U430 ( .A(KEYINPUT76), .B(G106GAT), .Z(n376) );
  XNOR2_X1 U431 ( .A(G99GAT), .B(G162GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n391) );
  XOR2_X1 U433 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n378) );
  XNOR2_X1 U434 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U436 ( .A(KEYINPUT74), .B(KEYINPUT77), .Z(n380) );
  XNOR2_X1 U437 ( .A(KEYINPUT75), .B(KEYINPUT11), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U439 ( .A(n382), .B(n381), .Z(n389) );
  XOR2_X1 U440 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U443 ( .A(G43GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n394) );
  INV_X1 U446 ( .A(n392), .ZN(n393) );
  XOR2_X1 U447 ( .A(n394), .B(n393), .Z(n549) );
  INV_X1 U448 ( .A(n549), .ZN(n397) );
  NAND2_X1 U449 ( .A1(n395), .A2(n397), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n396), .B(KEYINPUT47), .ZN(n402) );
  XNOR2_X1 U451 ( .A(KEYINPUT36), .B(n397), .ZN(n578) );
  INV_X1 U452 ( .A(n560), .ZN(n574) );
  NOR2_X1 U453 ( .A1(n578), .A2(n574), .ZN(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT45), .B(n398), .ZN(n399) );
  NAND2_X1 U455 ( .A1(n399), .A2(n571), .ZN(n400) );
  XNOR2_X1 U456 ( .A(KEYINPUT72), .B(n542), .ZN(n553) );
  NOR2_X1 U457 ( .A1(n400), .A2(n553), .ZN(n401) );
  NOR2_X1 U458 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U459 ( .A(KEYINPUT48), .B(n403), .ZN(n521) );
  NOR2_X1 U460 ( .A1(n513), .A2(n521), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n404), .B(KEYINPUT54), .ZN(n429) );
  XOR2_X1 U462 ( .A(KEYINPUT3), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U463 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U465 ( .A(KEYINPUT90), .B(n407), .Z(n441) );
  XOR2_X1 U466 ( .A(KEYINPUT96), .B(G148GAT), .Z(n409) );
  XNOR2_X1 U467 ( .A(G113GAT), .B(G120GAT), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G134GAT), .Z(n411) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G141GAT), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n427) );
  XOR2_X1 U473 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n415) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(G57GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U479 ( .A(n419), .B(n418), .Z(n425) );
  XOR2_X1 U480 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n421) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n441), .B(n428), .ZN(n522) );
  NAND2_X1 U487 ( .A1(n429), .A2(n522), .ZN(n563) );
  XOR2_X1 U488 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n431) );
  XNOR2_X1 U489 ( .A(KEYINPUT22), .B(KEYINPUT86), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U491 ( .A(n432), .B(KEYINPUT23), .Z(n435) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U494 ( .A(KEYINPUT91), .B(n436), .Z(n438) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U497 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n462) );
  NOR2_X1 U500 ( .A1(n563), .A2(n462), .ZN(n448) );
  XNOR2_X1 U501 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n446) );
  NOR2_X1 U502 ( .A1(n525), .A2(n449), .ZN(n561) );
  NAND2_X1 U503 ( .A1(n561), .A2(n549), .ZN(n453) );
  XOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n451) );
  INV_X1 U505 ( .A(G36GAT), .ZN(n475) );
  NAND2_X1 U506 ( .A1(n462), .A2(n525), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT26), .ZN(n564) );
  XNOR2_X1 U508 ( .A(n513), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT27), .ZN(n524) );
  INV_X1 U510 ( .A(n524), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n564), .A2(n456), .ZN(n461) );
  NOR2_X1 U512 ( .A1(n525), .A2(n513), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT25), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n459), .A2(n522), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n461), .A2(n460), .ZN(n467) );
  XOR2_X1 U516 ( .A(n462), .B(KEYINPUT28), .Z(n527) );
  NAND2_X1 U517 ( .A1(n527), .A2(n524), .ZN(n464) );
  XNOR2_X1 U518 ( .A(KEYINPUT85), .B(n525), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n465), .A2(n522), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n468), .B(KEYINPUT100), .ZN(n477) );
  NOR2_X1 U523 ( .A1(n578), .A2(n560), .ZN(n469) );
  AND2_X1 U524 ( .A1(n477), .A2(n469), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT37), .ZN(n511) );
  NAND2_X1 U526 ( .A1(n553), .A2(n571), .ZN(n479) );
  NOR2_X1 U527 ( .A1(n511), .A2(n479), .ZN(n472) );
  XNOR2_X1 U528 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n513), .A2(n496), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT106), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(G1329GAT) );
  NOR2_X1 U532 ( .A1(n549), .A2(n574), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT16), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n500) );
  OR2_X1 U535 ( .A1(n479), .A2(n500), .ZN(n487) );
  NOR2_X1 U536 ( .A1(n522), .A2(n487), .ZN(n480) );
  XOR2_X1 U537 ( .A(n480), .B(KEYINPUT34), .Z(n481) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U539 ( .A1(n513), .A2(n487), .ZN(n483) );
  XNOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1325GAT) );
  NOR2_X1 U542 ( .A1(n525), .A2(n487), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n527), .A2(n487), .ZN(n489) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  NOR2_X1 U549 ( .A1(n496), .A2(n522), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n525), .A2(n496), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n498) );
  NOR2_X1 U558 ( .A1(n527), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  NAND2_X1 U561 ( .A1(n566), .A2(n556), .ZN(n510) );
  NOR2_X1 U562 ( .A1(n510), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT110), .B(n501), .Z(n506) );
  NOR2_X1 U564 ( .A1(n506), .A2(n522), .ZN(n502) );
  XOR2_X1 U565 ( .A(n502), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n506), .ZN(n504) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n525), .A2(n506), .ZN(n505) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  XNOR2_X1 U571 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n508) );
  NOR2_X1 U572 ( .A1(n527), .A2(n506), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  OR2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U576 ( .A1(n522), .A2(n518), .ZN(n512) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n512), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n518), .ZN(n514) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n518), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G99GAT), .B(n517), .ZN(G1338GAT) );
  NOR2_X1 U584 ( .A1(n527), .A2(n518), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n541) );
  NOR2_X1 U589 ( .A1(n525), .A2(n541), .ZN(n526) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(n526), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(KEYINPUT115), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n553), .A2(n538), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n532) );
  NAND2_X1 U596 ( .A1(n538), .A2(n556), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT116), .Z(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n536) );
  NAND2_X1 U601 ( .A1(n538), .A2(n560), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n549), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n564), .A2(n541), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n550), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n545) );
  NAND2_X1 U611 ( .A1(n550), .A2(n556), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n550), .A2(n560), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT120), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  XOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT123), .Z(n555) );
  NAND2_X1 U621 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  NAND2_X1 U624 ( .A1(n561), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT125), .B(n565), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n566), .A2(n577), .ZN(n570) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT126), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n577), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

