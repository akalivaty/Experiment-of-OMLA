

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741;

  XNOR2_X1 U378 ( .A(n487), .B(n488), .ZN(n724) );
  NOR2_X1 U379 ( .A1(n666), .A2(n665), .ZN(n663) );
  INV_X1 U380 ( .A(G953), .ZN(n718) );
  INV_X2 U381 ( .A(G143), .ZN(n445) );
  AND2_X2 U382 ( .A1(n408), .A2(n362), .ZN(n600) );
  NOR2_X1 U383 ( .A1(n662), .A2(n547), .ZN(n619) );
  NAND2_X1 U384 ( .A1(n586), .A2(n662), .ZN(n641) );
  NOR2_X1 U385 ( .A1(n543), .A2(n418), .ZN(n417) );
  XNOR2_X1 U386 ( .A(n518), .B(n363), .ZN(n418) );
  XNOR2_X1 U387 ( .A(n486), .B(n485), .ZN(n543) );
  XNOR2_X1 U388 ( .A(n539), .B(KEYINPUT108), .ZN(n631) );
  XNOR2_X1 U389 ( .A(n474), .B(n373), .ZN(n487) );
  NOR2_X2 U390 ( .A1(n736), .A2(KEYINPUT44), .ZN(n386) );
  XNOR2_X2 U391 ( .A(n724), .B(G146), .ZN(n515) );
  NOR2_X1 U392 ( .A1(G902), .A2(G237), .ZN(n449) );
  XOR2_X1 U393 ( .A(KEYINPUT4), .B(G131), .Z(n488) );
  XNOR2_X1 U394 ( .A(n372), .B(G140), .ZN(n497) );
  INV_X1 U395 ( .A(G137), .ZN(n372) );
  NOR2_X1 U396 ( .A1(n614), .A2(n460), .ZN(n552) );
  XNOR2_X1 U397 ( .A(n406), .B(n404), .ZN(n498) );
  XNOR2_X1 U398 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n406) );
  NOR2_X1 U399 ( .A1(n405), .A2(G953), .ZN(n404) );
  INV_X1 U400 ( .A(G234), .ZN(n405) );
  XNOR2_X1 U401 ( .A(n421), .B(n419), .ZN(n699) );
  XNOR2_X1 U402 ( .A(n357), .B(n420), .ZN(n419) );
  XNOR2_X1 U403 ( .A(n471), .B(n422), .ZN(n421) );
  XNOR2_X1 U404 ( .A(n465), .B(n467), .ZN(n420) );
  XNOR2_X1 U405 ( .A(n503), .B(KEYINPUT25), .ZN(n432) );
  OR2_X1 U406 ( .A1(n709), .A2(G902), .ZN(n433) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n504) );
  INV_X1 U408 ( .A(KEYINPUT89), .ZN(n395) );
  INV_X1 U409 ( .A(KEYINPUT67), .ZN(n385) );
  XOR2_X1 U410 ( .A(G902), .B(KEYINPUT15), .Z(n460) );
  XNOR2_X1 U411 ( .A(n497), .B(n360), .ZN(n371) );
  NAND2_X1 U412 ( .A1(n596), .A2(n643), .ZN(n602) );
  XNOR2_X1 U413 ( .A(n378), .B(n377), .ZN(n596) );
  INV_X1 U414 ( .A(KEYINPUT48), .ZN(n377) );
  NAND2_X1 U415 ( .A1(n381), .A2(n379), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n413), .B(n412), .ZN(n536) );
  XNOR2_X1 U417 ( .A(G478), .B(KEYINPUT107), .ZN(n412) );
  OR2_X1 U418 ( .A1(n705), .A2(G902), .ZN(n413) );
  OR2_X2 U419 ( .A1(n367), .A2(n364), .ZN(n563) );
  NAND2_X1 U420 ( .A1(n369), .A2(n368), .ZN(n367) );
  NAND2_X1 U421 ( .A1(n495), .A2(n366), .ZN(n365) );
  INV_X1 U422 ( .A(n519), .ZN(n669) );
  XOR2_X1 U423 ( .A(G116), .B(G107), .Z(n478) );
  INV_X1 U424 ( .A(KEYINPUT76), .ZN(n438) );
  XNOR2_X1 U425 ( .A(n358), .B(n441), .ZN(n511) );
  XNOR2_X1 U426 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U427 ( .A(G113), .B(G104), .ZN(n442) );
  XOR2_X1 U428 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n476) );
  XNOR2_X1 U429 ( .A(G122), .B(KEYINPUT106), .ZN(n475) );
  INV_X1 U430 ( .A(G134), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n712), .B(n389), .ZN(n614) );
  XNOR2_X1 U432 ( .A(n390), .B(n444), .ZN(n389) );
  XNOR2_X1 U433 ( .A(n447), .B(n391), .ZN(n390) );
  XNOR2_X1 U434 ( .A(n552), .B(n551), .ZN(n582) );
  NOR2_X1 U435 ( .A1(n585), .A2(n397), .ZN(n591) );
  NAND2_X1 U436 ( .A1(n631), .A2(n650), .ZN(n397) );
  XNOR2_X1 U437 ( .A(n525), .B(KEYINPUT34), .ZN(n431) );
  XNOR2_X1 U438 ( .A(n473), .B(n423), .ZN(n538) );
  XNOR2_X1 U439 ( .A(n472), .B(n424), .ZN(n423) );
  INV_X1 U440 ( .A(G475), .ZN(n424) );
  BUF_X1 U441 ( .A(n521), .Z(n662) );
  XNOR2_X1 U442 ( .A(KEYINPUT22), .B(KEYINPUT75), .ZN(n485) );
  XNOR2_X1 U443 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U444 ( .A(n427), .B(n425), .ZN(n500) );
  INV_X1 U445 ( .A(KEYINPUT64), .ZN(n599) );
  NOR2_X1 U446 ( .A1(G952), .A2(n718), .ZN(n711) );
  INV_X1 U447 ( .A(KEYINPUT90), .ZN(n388) );
  XNOR2_X1 U448 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U449 ( .A(n590), .B(n380), .ZN(n379) );
  INV_X1 U450 ( .A(KEYINPUT69), .ZN(n380) );
  NOR2_X1 U451 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U452 ( .A(n382), .B(KEYINPUT46), .ZN(n381) );
  NOR2_X1 U453 ( .A1(n739), .A2(n741), .ZN(n382) );
  NAND2_X1 U454 ( .A1(n370), .A2(G902), .ZN(n368) );
  XNOR2_X1 U455 ( .A(G137), .B(G116), .ZN(n507) );
  XOR2_X1 U456 ( .A(KEYINPUT98), .B(G113), .Z(n508) );
  XOR2_X1 U457 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n506) );
  XNOR2_X1 U458 ( .A(n466), .B(n468), .ZN(n422) );
  XNOR2_X1 U459 ( .A(G143), .B(G131), .ZN(n464) );
  OR2_X1 U460 ( .A1(n597), .A2(n598), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n392), .B(n448), .ZN(n391) );
  XNOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT79), .ZN(n392) );
  NAND2_X1 U463 ( .A1(n536), .A2(n538), .ZN(n653) );
  NOR2_X1 U464 ( .A1(n653), .A2(n665), .ZN(n483) );
  NOR2_X1 U465 ( .A1(n602), .A2(n597), .ZN(n731) );
  XNOR2_X1 U466 ( .A(n435), .B(n428), .ZN(n427) );
  XNOR2_X1 U467 ( .A(KEYINPUT23), .B(KEYINPUT94), .ZN(n435) );
  XNOR2_X1 U468 ( .A(KEYINPUT24), .B(G110), .ZN(n428) );
  XNOR2_X1 U469 ( .A(n426), .B(G128), .ZN(n425) );
  INV_X1 U470 ( .A(G119), .ZN(n426) );
  XNOR2_X1 U471 ( .A(n491), .B(n371), .ZN(n493) );
  NOR2_X1 U472 ( .A1(n602), .A2(n356), .ZN(n403) );
  AND2_X1 U473 ( .A1(n578), .A2(n651), .ZN(n557) );
  INV_X1 U474 ( .A(KEYINPUT80), .ZN(n363) );
  XNOR2_X1 U475 ( .A(n552), .B(n401), .ZN(n594) );
  INV_X1 U476 ( .A(n551), .ZN(n401) );
  AND2_X1 U477 ( .A1(n376), .A2(n374), .ZN(n578) );
  XNOR2_X1 U478 ( .A(n554), .B(n375), .ZN(n374) );
  NOR2_X1 U479 ( .A1(n555), .A2(n558), .ZN(n376) );
  INV_X1 U480 ( .A(KEYINPUT30), .ZN(n375) );
  NAND2_X1 U481 ( .A1(n582), .A2(n650), .ZN(n402) );
  XNOR2_X1 U482 ( .A(n605), .B(KEYINPUT62), .ZN(n606) );
  XNOR2_X1 U483 ( .A(n440), .B(n478), .ZN(n393) );
  XNOR2_X1 U484 ( .A(n511), .B(n470), .ZN(n394) );
  XNOR2_X1 U485 ( .A(n481), .B(n482), .ZN(n705) );
  XNOR2_X1 U486 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U487 ( .A(n411), .B(n410), .ZN(n586) );
  INV_X1 U488 ( .A(KEYINPUT36), .ZN(n410) );
  NAND2_X1 U489 ( .A1(n591), .A2(n582), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n526), .B(KEYINPUT85), .ZN(n429) );
  NOR2_X1 U491 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U492 ( .A1(n415), .A2(n359), .ZN(n625) );
  XNOR2_X1 U493 ( .A(n708), .B(n398), .ZN(n710) );
  XNOR2_X1 U494 ( .A(n709), .B(KEYINPUT122), .ZN(n398) );
  XOR2_X1 U495 ( .A(KEYINPUT81), .B(n601), .Z(n356) );
  XOR2_X1 U496 ( .A(n464), .B(G140), .Z(n357) );
  XOR2_X1 U497 ( .A(G101), .B(G119), .Z(n358) );
  AND2_X1 U498 ( .A1(n592), .A2(n520), .ZN(n359) );
  AND2_X1 U499 ( .A1(n718), .A2(G227), .ZN(n360) );
  INV_X1 U500 ( .A(G902), .ZN(n366) );
  XOR2_X1 U501 ( .A(n451), .B(KEYINPUT19), .Z(n361) );
  XNOR2_X1 U502 ( .A(n394), .B(n393), .ZN(n712) );
  XOR2_X1 U503 ( .A(n437), .B(KEYINPUT65), .Z(n362) );
  NAND2_X1 U504 ( .A1(n692), .A2(n370), .ZN(n369) );
  XNOR2_X2 U505 ( .A(n515), .B(n494), .ZN(n692) );
  XNOR2_X2 U506 ( .A(n563), .B(KEYINPUT1), .ZN(n521) );
  NOR2_X1 U507 ( .A1(n692), .A2(n365), .ZN(n364) );
  INV_X1 U508 ( .A(n495), .ZN(n370) );
  XNOR2_X2 U509 ( .A(n445), .B(G128), .ZN(n474) );
  XNOR2_X1 U510 ( .A(n383), .B(KEYINPUT74), .ZN(n414) );
  NAND2_X1 U511 ( .A1(n387), .A2(n384), .ZN(n383) );
  XNOR2_X1 U512 ( .A(n386), .B(n385), .ZN(n384) );
  XNOR2_X1 U513 ( .A(n527), .B(n388), .ZN(n387) );
  NAND2_X1 U514 ( .A1(n737), .A2(n625), .ZN(n527) );
  XNOR2_X1 U515 ( .A(n417), .B(n416), .ZN(n737) );
  NOR2_X1 U516 ( .A1(n533), .A2(n484), .ZN(n486) );
  XNOR2_X2 U517 ( .A(n524), .B(n523), .ZN(n661) );
  NAND2_X1 U518 ( .A1(n431), .A2(n577), .ZN(n430) );
  XNOR2_X1 U519 ( .A(n396), .B(n395), .ZN(n529) );
  NAND2_X1 U520 ( .A1(n736), .A2(KEYINPUT44), .ZN(n396) );
  AND2_X4 U521 ( .A1(n604), .A2(n603), .ZN(n707) );
  NAND2_X1 U522 ( .A1(n731), .A2(n719), .ZN(n645) );
  XNOR2_X2 U523 ( .A(n600), .B(n599), .ZN(n604) );
  XNOR2_X1 U524 ( .A(n399), .B(n703), .ZN(G60) );
  NOR2_X2 U525 ( .A1(n702), .A2(n711), .ZN(n399) );
  XNOR2_X1 U526 ( .A(n400), .B(n618), .ZN(G51) );
  NOR2_X2 U527 ( .A1(n617), .A2(n711), .ZN(n400) );
  INV_X1 U528 ( .A(n458), .ZN(n571) );
  XNOR2_X2 U529 ( .A(n402), .B(n361), .ZN(n458) );
  AND2_X1 U530 ( .A1(n719), .A2(n403), .ZN(n649) );
  XNOR2_X2 U531 ( .A(n550), .B(KEYINPUT45), .ZN(n719) );
  NAND2_X1 U532 ( .A1(n719), .A2(n407), .ZN(n408) );
  NOR2_X1 U533 ( .A1(n602), .A2(n409), .ZN(n407) );
  NAND2_X1 U534 ( .A1(n414), .A2(n434), .ZN(n550) );
  INV_X1 U535 ( .A(n543), .ZN(n415) );
  INV_X1 U536 ( .A(KEYINPUT32), .ZN(n416) );
  XNOR2_X2 U537 ( .A(n430), .B(n429), .ZN(n736) );
  XNOR2_X2 U538 ( .A(n433), .B(n432), .ZN(n666) );
  XNOR2_X1 U539 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X2 U540 ( .A1(n608), .A2(n711), .ZN(n610) );
  AND2_X1 U541 ( .A1(n436), .A2(n549), .ZN(n434) );
  AND2_X1 U542 ( .A1(n529), .A2(n528), .ZN(n436) );
  INV_X1 U543 ( .A(n469), .ZN(n443) );
  XNOR2_X1 U544 ( .A(n510), .B(n509), .ZN(n513) );
  XNOR2_X1 U545 ( .A(n474), .B(n446), .ZN(n447) );
  XNOR2_X1 U546 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U547 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U548 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n523) );
  XNOR2_X1 U549 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U550 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n568) );
  INV_X1 U551 ( .A(KEYINPUT63), .ZN(n609) );
  XNOR2_X1 U552 ( .A(n569), .B(n568), .ZN(n739) );
  NAND2_X1 U553 ( .A1(n460), .A2(KEYINPUT2), .ZN(n437) );
  XNOR2_X1 U554 ( .A(G110), .B(KEYINPUT16), .ZN(n439) );
  XNOR2_X1 U555 ( .A(n442), .B(G122), .ZN(n470) );
  XNOR2_X1 U556 ( .A(n443), .B(KEYINPUT17), .ZN(n444) );
  AND2_X1 U557 ( .A1(G224), .A2(n718), .ZN(n446) );
  INV_X1 U558 ( .A(KEYINPUT18), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n449), .B(KEYINPUT77), .ZN(n450) );
  NAND2_X1 U560 ( .A1(G210), .A2(n450), .ZN(n551) );
  NAND2_X1 U561 ( .A1(G214), .A2(n450), .ZN(n650) );
  INV_X1 U562 ( .A(KEYINPUT66), .ZN(n451) );
  NAND2_X1 U563 ( .A1(G898), .A2(G953), .ZN(n456) );
  NAND2_X1 U564 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U565 ( .A(n452), .B(KEYINPUT14), .ZN(n683) );
  OR2_X1 U566 ( .A1(n718), .A2(G902), .ZN(n453) );
  NAND2_X1 U567 ( .A1(n683), .A2(n453), .ZN(n455) );
  NOR2_X1 U568 ( .A1(G953), .A2(G952), .ZN(n454) );
  NOR2_X1 U569 ( .A1(n455), .A2(n454), .ZN(n553) );
  AND2_X1 U570 ( .A1(n456), .A2(n553), .ZN(n457) );
  NAND2_X1 U571 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X2 U572 ( .A(n459), .B(KEYINPUT0), .ZN(n533) );
  XOR2_X1 U573 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n462) );
  INV_X1 U574 ( .A(n460), .ZN(n598) );
  NAND2_X1 U575 ( .A1(G234), .A2(n598), .ZN(n461) );
  XNOR2_X1 U576 ( .A(n462), .B(n461), .ZN(n502) );
  NAND2_X1 U577 ( .A1(n502), .A2(G221), .ZN(n463) );
  XNOR2_X1 U578 ( .A(n463), .B(KEYINPUT21), .ZN(n665) );
  XOR2_X1 U579 ( .A(KEYINPUT103), .B(KEYINPUT101), .Z(n466) );
  NAND2_X1 U580 ( .A1(G214), .A2(n504), .ZN(n465) );
  XOR2_X1 U581 ( .A(KEYINPUT100), .B(KEYINPUT102), .Z(n468) );
  XNOR2_X1 U582 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n467) );
  XNOR2_X1 U583 ( .A(KEYINPUT10), .B(n469), .ZN(n496) );
  XNOR2_X1 U584 ( .A(n470), .B(n496), .ZN(n471) );
  NOR2_X1 U585 ( .A1(G902), .A2(n699), .ZN(n473) );
  XNOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U588 ( .A(n487), .B(n477), .ZN(n482) );
  XOR2_X1 U589 ( .A(n478), .B(KEYINPUT105), .Z(n480) );
  NAND2_X1 U590 ( .A1(G217), .A2(n498), .ZN(n479) );
  XNOR2_X1 U591 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U592 ( .A(KEYINPUT110), .B(n483), .Z(n484) );
  XOR2_X1 U593 ( .A(G107), .B(G110), .Z(n490) );
  XNOR2_X1 U594 ( .A(G101), .B(G104), .ZN(n489) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U596 ( .A(KEYINPUT78), .B(KEYINPUT93), .ZN(n492) );
  XNOR2_X1 U597 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U598 ( .A(KEYINPUT71), .B(G469), .ZN(n495) );
  INV_X1 U599 ( .A(n662), .ZN(n592) );
  XNOR2_X1 U600 ( .A(n497), .B(n496), .ZN(n725) );
  NAND2_X1 U601 ( .A1(G221), .A2(n498), .ZN(n499) );
  XNOR2_X1 U602 ( .A(n725), .B(n501), .ZN(n709) );
  NAND2_X1 U603 ( .A1(G217), .A2(n502), .ZN(n503) );
  INV_X1 U604 ( .A(n666), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n504), .A2(G210), .ZN(n505) );
  XNOR2_X1 U606 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X1 U607 ( .A(n508), .B(n507), .ZN(n509) );
  INV_X1 U608 ( .A(n511), .ZN(n512) );
  XNOR2_X1 U609 ( .A(n515), .B(n514), .ZN(n605) );
  NOR2_X1 U610 ( .A1(G902), .A2(n605), .ZN(n516) );
  XNOR2_X1 U611 ( .A(n516), .B(G472), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n519), .B(KEYINPUT6), .ZN(n522) );
  OR2_X1 U613 ( .A1(n545), .A2(n522), .ZN(n517) );
  NOR2_X1 U614 ( .A1(n592), .A2(n517), .ZN(n518) );
  INV_X1 U615 ( .A(n669), .ZN(n561) );
  AND2_X1 U616 ( .A1(n561), .A2(n666), .ZN(n520) );
  AND2_X2 U617 ( .A1(n521), .A2(n663), .ZN(n532) );
  NAND2_X1 U618 ( .A1(n532), .A2(n522), .ZN(n524) );
  NOR2_X2 U619 ( .A1(n661), .A2(n533), .ZN(n525) );
  NOR2_X1 U620 ( .A1(n538), .A2(n536), .ZN(n577) );
  INV_X1 U621 ( .A(KEYINPUT35), .ZN(n526) );
  NAND2_X1 U622 ( .A1(n527), .A2(KEYINPUT44), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n563), .A2(n663), .ZN(n530) );
  XNOR2_X1 U624 ( .A(KEYINPUT96), .B(n530), .ZN(n555) );
  NOR2_X1 U625 ( .A1(n555), .A2(n533), .ZN(n531) );
  NAND2_X1 U626 ( .A1(n531), .A2(n561), .ZN(n621) );
  NAND2_X1 U627 ( .A1(n669), .A2(n532), .ZN(n673) );
  NOR2_X1 U628 ( .A1(n533), .A2(n673), .ZN(n535) );
  XOR2_X1 U629 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n534) );
  XNOR2_X1 U630 ( .A(n535), .B(n534), .ZN(n637) );
  NAND2_X1 U631 ( .A1(n621), .A2(n637), .ZN(n541) );
  INV_X1 U632 ( .A(n536), .ZN(n537) );
  NAND2_X1 U633 ( .A1(n537), .A2(n538), .ZN(n638) );
  INV_X1 U634 ( .A(n638), .ZN(n626) );
  NOR2_X1 U635 ( .A1(n626), .A2(n631), .ZN(n655) );
  INV_X1 U636 ( .A(n655), .ZN(n540) );
  NAND2_X1 U637 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U638 ( .A(n542), .B(KEYINPUT109), .ZN(n548) );
  NOR2_X1 U639 ( .A1(n522), .A2(n543), .ZN(n544) );
  XNOR2_X1 U640 ( .A(n544), .B(KEYINPUT88), .ZN(n546) );
  NAND2_X1 U641 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U642 ( .A1(n548), .A2(n619), .ZN(n549) );
  XNOR2_X1 U643 ( .A(KEYINPUT38), .B(n594), .ZN(n651) );
  NAND2_X1 U644 ( .A1(G953), .A2(G900), .ZN(n729) );
  NAND2_X1 U645 ( .A1(n553), .A2(n729), .ZN(n558) );
  NAND2_X1 U646 ( .A1(n669), .A2(n650), .ZN(n554) );
  XNOR2_X1 U647 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n556) );
  XNOR2_X1 U648 ( .A(n557), .B(n556), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n567), .A2(n626), .ZN(n642) );
  INV_X1 U650 ( .A(n642), .ZN(n597) );
  NOR2_X1 U651 ( .A1(n665), .A2(n558), .ZN(n559) );
  XNOR2_X1 U652 ( .A(KEYINPUT70), .B(n559), .ZN(n560) );
  NAND2_X1 U653 ( .A1(n560), .A2(n666), .ZN(n583) );
  NOR2_X1 U654 ( .A1(n583), .A2(n561), .ZN(n562) );
  XNOR2_X1 U655 ( .A(KEYINPUT28), .B(n562), .ZN(n564) );
  NAND2_X1 U656 ( .A1(n564), .A2(n563), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n651), .A2(n650), .ZN(n654) );
  NOR2_X1 U658 ( .A1(n653), .A2(n654), .ZN(n565) );
  XNOR2_X1 U659 ( .A(n565), .B(KEYINPUT41), .ZN(n677) );
  NOR2_X1 U660 ( .A1(n570), .A2(n677), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n566), .B(KEYINPUT42), .ZN(n741) );
  NAND2_X1 U662 ( .A1(n567), .A2(n631), .ZN(n569) );
  NAND2_X1 U663 ( .A1(KEYINPUT84), .A2(n655), .ZN(n572) );
  NOR2_X1 U664 ( .A1(n571), .A2(n570), .ZN(n632) );
  NAND2_X1 U665 ( .A1(n572), .A2(n632), .ZN(n573) );
  NAND2_X1 U666 ( .A1(n573), .A2(KEYINPUT47), .ZN(n576) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(n655), .ZN(n574) );
  NAND2_X1 U668 ( .A1(n574), .A2(n632), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n576), .A2(n575), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U671 ( .A1(n594), .A2(n579), .ZN(n630) );
  AND2_X1 U672 ( .A1(n655), .A2(KEYINPUT47), .ZN(n580) );
  NOR2_X1 U673 ( .A1(KEYINPUT84), .A2(n580), .ZN(n581) );
  NOR2_X1 U674 ( .A1(n630), .A2(n581), .ZN(n587) );
  INV_X1 U675 ( .A(n583), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n584), .A2(n522), .ZN(n585) );
  NAND2_X1 U677 ( .A1(n587), .A2(n641), .ZN(n588) );
  NAND2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U679 ( .A(n593), .B(KEYINPUT43), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n595), .A2(n594), .ZN(n643) );
  NAND2_X1 U681 ( .A1(KEYINPUT2), .A2(n642), .ZN(n601) );
  INV_X1 U682 ( .A(n649), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n707), .A2(G472), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n610), .B(n609), .ZN(G57) );
  NAND2_X1 U685 ( .A1(n707), .A2(G210), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n612) );
  XNOR2_X1 U687 ( .A(KEYINPUT91), .B(KEYINPUT83), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT86), .B(KEYINPUT56), .ZN(n618) );
  XOR2_X1 U692 ( .A(G101), .B(n619), .Z(G3) );
  INV_X1 U693 ( .A(n631), .ZN(n635) );
  NOR2_X1 U694 ( .A1(n635), .A2(n621), .ZN(n620) );
  XOR2_X1 U695 ( .A(G104), .B(n620), .Z(G6) );
  NOR2_X1 U696 ( .A1(n638), .A2(n621), .ZN(n623) );
  XNOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U699 ( .A(G107), .B(n624), .ZN(G9) );
  XNOR2_X1 U700 ( .A(G110), .B(n625), .ZN(G12) );
  XOR2_X1 U701 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n628) );
  NAND2_X1 U702 ( .A1(n626), .A2(n632), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U704 ( .A(G128), .B(n629), .ZN(G30) );
  XOR2_X1 U705 ( .A(G143), .B(n630), .Z(G45) );
  XOR2_X1 U706 ( .A(G146), .B(KEYINPUT113), .Z(n634) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(G48) );
  NOR2_X1 U709 ( .A1(n635), .A2(n637), .ZN(n636) );
  XOR2_X1 U710 ( .A(G113), .B(n636), .Z(G15) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U712 ( .A(G116), .B(n639), .Z(G18) );
  XOR2_X1 U713 ( .A(G125), .B(KEYINPUT37), .Z(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G27) );
  XNOR2_X1 U715 ( .A(G134), .B(n642), .ZN(G36) );
  XNOR2_X1 U716 ( .A(G140), .B(n643), .ZN(G42) );
  NOR2_X1 U717 ( .A1(n677), .A2(n661), .ZN(n644) );
  NOR2_X1 U718 ( .A1(G953), .A2(n644), .ZN(n689) );
  INV_X1 U719 ( .A(KEYINPUT2), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U721 ( .A(KEYINPUT82), .B(n647), .Z(n648) );
  NOR2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n687) );
  NOR2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT116), .ZN(n657) );
  NOR2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(n659), .Z(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n680) );
  XOR2_X1 U730 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n676) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U732 ( .A(KEYINPUT50), .B(n664), .Z(n672) );
  NAND2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(KEYINPUT49), .B(n667), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U736 ( .A(KEYINPUT114), .B(n670), .ZN(n671) );
  NAND2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U739 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U742 ( .A(n681), .B(KEYINPUT118), .ZN(n682) );
  XNOR2_X1 U743 ( .A(n682), .B(KEYINPUT52), .ZN(n685) );
  NAND2_X1 U744 ( .A1(n683), .A2(G952), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n690), .B(KEYINPUT119), .ZN(n691) );
  XNOR2_X1 U749 ( .A(KEYINPUT53), .B(n691), .ZN(G75) );
  XNOR2_X1 U750 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n692), .B(KEYINPUT57), .ZN(n693) );
  XNOR2_X1 U752 ( .A(n694), .B(n693), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n707), .A2(G469), .ZN(n695) );
  XOR2_X1 U754 ( .A(n696), .B(n695), .Z(n697) );
  NOR2_X1 U755 ( .A1(n711), .A2(n697), .ZN(G54) );
  NAND2_X1 U756 ( .A1(n707), .A2(G475), .ZN(n701) );
  XOR2_X1 U757 ( .A(KEYINPUT59), .B(KEYINPUT92), .Z(n698) );
  XOR2_X1 U758 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n703) );
  NAND2_X1 U759 ( .A1(G478), .A2(n707), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U761 ( .A1(n711), .A2(n706), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n707), .A2(G217), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(G66) );
  OR2_X1 U764 ( .A1(G898), .A2(n718), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n714), .B(KEYINPUT124), .ZN(n723) );
  XOR2_X1 U767 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n716) );
  NAND2_X1 U768 ( .A1(G224), .A2(G953), .ZN(n715) );
  XNOR2_X1 U769 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n717), .A2(G898), .ZN(n721) );
  NAND2_X1 U771 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U772 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U773 ( .A(n723), .B(n722), .Z(G69) );
  BUF_X1 U774 ( .A(n724), .Z(n726) );
  XOR2_X1 U775 ( .A(n726), .B(n725), .Z(n730) );
  XNOR2_X1 U776 ( .A(n730), .B(G227), .ZN(n727) );
  XNOR2_X1 U777 ( .A(KEYINPUT125), .B(n727), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n734) );
  XOR2_X1 U779 ( .A(n731), .B(n730), .Z(n732) );
  NOR2_X1 U780 ( .A1(G953), .A2(n732), .ZN(n733) );
  NOR2_X1 U781 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U783 ( .A(n736), .B(G122), .Z(G24) );
  BUF_X1 U784 ( .A(n737), .Z(n738) );
  XNOR2_X1 U785 ( .A(G119), .B(n738), .ZN(G21) );
  XNOR2_X1 U786 ( .A(G131), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n740), .B(n739), .ZN(G33) );
  XOR2_X1 U788 ( .A(G137), .B(n741), .Z(G39) );
endmodule

