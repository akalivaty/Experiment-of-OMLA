//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n213), .B(new_n219), .C1(G116), .C2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G58), .B2(G232), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n205), .B(new_n224), .C1(KEYINPUT65), .C2(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n204), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n210), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n218), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n217), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT25), .B1(new_n251), .B2(new_n217), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n217), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n203), .A2(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n250), .A2(new_n255), .A3(new_n228), .A4(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n253), .A2(new_n254), .B1(G107), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n203), .B(G45), .C1(new_n260), .C2(KEYINPUT5), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT5), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G41), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT77), .A3(new_n203), .A4(G45), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n267), .A2(G274), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G250), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n274), .B1(G257), .B2(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G294), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n269), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n263), .A2(new_n270), .A3(new_n266), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G264), .A3(new_n269), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n271), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G200), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n271), .A2(new_n287), .A3(new_n281), .A4(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT81), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n204), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT22), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(KEYINPUT22), .A3(new_n204), .A4(G87), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT23), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n217), .A3(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n217), .A2(KEYINPUT68), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G107), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n204), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n302), .B(new_n303), .C1(new_n307), .C2(new_n301), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT24), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n300), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n293), .A2(new_n299), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT24), .B1(new_n312), .B2(new_n308), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n256), .A2(new_n228), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n290), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n315), .ZN(new_n317));
  AOI211_X1 g0117(.A(KEYINPUT81), .B(new_n317), .C1(new_n311), .C2(new_n313), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n259), .B(new_n289), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n259), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n310), .B1(new_n300), .B2(new_n309), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n312), .A2(new_n308), .A3(KEYINPUT24), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT81), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n314), .A2(new_n290), .A3(new_n315), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n284), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G179), .B2(new_n284), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n319), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n273), .A2(G222), .ZN(new_n332));
  INV_X1    g0132(.A(G223), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n298), .B(new_n332), .C1(new_n333), .C2(new_n273), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(new_n280), .C1(G77), .C2(new_n298), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n336));
  INV_X1    g0136(.A(G274), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n269), .A2(new_n336), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n335), .B(new_n339), .C1(new_n222), .C2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n287), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT70), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT10), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n251), .A2(new_n221), .ZN(new_n349));
  INV_X1    g0149(.A(G150), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G20), .A2(G33), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR3_X1   g0152(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n350), .A2(new_n352), .B1(new_n353), .B2(new_n204), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT8), .B(G58), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n204), .A2(G33), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n315), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n251), .A2(new_n315), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(KEYINPUT66), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n204), .A2(G1), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT67), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(KEYINPUT66), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n349), .B(new_n358), .C1(new_n365), .C2(new_n221), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT9), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n347), .A2(new_n348), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n343), .A2(new_n344), .A3(new_n367), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n348), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n341), .A2(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n341), .A2(new_n327), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G238), .A2(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n298), .B(new_n375), .C1(new_n234), .C2(G1698), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT68), .B(G107), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n280), .C1(new_n377), .C2(new_n298), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n339), .C1(new_n212), .C2(new_n340), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(G200), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n287), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n362), .A2(new_n315), .A3(new_n251), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G77), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT15), .B(G87), .Z(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n356), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n355), .A2(new_n352), .B1(new_n204), .B2(new_n211), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n315), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n383), .B(new_n388), .C1(G77), .C2(new_n250), .ZN(new_n389));
  OR3_X1    g0189(.A1(new_n380), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n371), .A2(new_n374), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT73), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G58), .B2(G68), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n351), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n296), .A2(new_n204), .A3(new_n297), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n297), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT72), .B1(new_n400), .B2(G68), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT72), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n402), .B(new_n215), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT16), .B(new_n395), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n392), .B(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G58), .A2(G68), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n409), .A2(new_n204), .B1(new_n410), .B2(new_n352), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n215), .B1(new_n398), .B2(new_n399), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n315), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n355), .ZN(new_n415));
  MUX2_X1   g0215(.A(new_n250), .B(new_n365), .S(new_n415), .Z(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT74), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G33), .A3(G87), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n333), .A2(new_n273), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n222), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(new_n275), .C2(new_n276), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n269), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G179), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n269), .A2(G232), .A3(new_n336), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n426), .A2(new_n427), .A3(new_n338), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n428), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(new_n421), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n296), .A2(new_n297), .B1(new_n222), .B2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n423), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n339), .B(new_n430), .C1(new_n433), .C2(new_n269), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n429), .B1(G169), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n417), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n417), .A2(KEYINPUT18), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n285), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n422), .A2(new_n425), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n428), .B1(new_n442), .B2(new_n280), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n287), .A3(new_n339), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(KEYINPUT75), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  AOI21_X1  g0246(.A(G200), .B1(new_n443), .B2(new_n339), .ZN(new_n447));
  NOR4_X1   g0247(.A1(new_n426), .A2(G190), .A3(new_n338), .A4(new_n428), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n414), .A2(new_n416), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT17), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n447), .A2(new_n448), .A3(new_n446), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT75), .B1(new_n441), .B2(new_n444), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g0254(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n455));
  NAND4_X1  g0255(.A1(new_n454), .A2(new_n414), .A3(new_n416), .A4(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n439), .A2(new_n440), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT13), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n222), .A2(new_n273), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n298), .B(new_n459), .C1(G232), .C2(new_n273), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n338), .B1(new_n462), .B2(new_n280), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n340), .A2(new_n216), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n458), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n269), .B1(new_n460), .B2(new_n461), .ZN(new_n467));
  NOR4_X1   g0267(.A1(new_n467), .A2(KEYINPUT13), .A3(new_n338), .A4(new_n464), .ZN(new_n468));
  OAI21_X1  g0268(.A(G169), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n470));
  INV_X1    g0270(.A(new_n466), .ZN(new_n471));
  INV_X1    g0271(.A(new_n468), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(G179), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT14), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(G169), .C1(new_n466), .C2(new_n468), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n382), .A2(G68), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT71), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n352), .A2(new_n221), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n356), .A2(new_n211), .B1(new_n204), .B2(G68), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n315), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g0281(.A(new_n481), .B(KEYINPUT11), .Z(new_n482));
  NOR2_X1   g0282(.A1(new_n250), .A2(G68), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT12), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n379), .A2(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n379), .A2(new_n327), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n389), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n457), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(G200), .B1(new_n466), .B2(new_n468), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n471), .A2(G190), .A3(new_n472), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n391), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n273), .A2(G257), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n298), .B(new_n498), .C1(new_n218), .C2(new_n273), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(new_n280), .C1(G303), .C2(new_n298), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n282), .A2(G270), .A3(new_n269), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n271), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  INV_X1    g0304(.A(G97), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n504), .B(new_n204), .C1(G33), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n244), .A2(G20), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n315), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n506), .A2(KEYINPUT20), .A3(new_n315), .A4(new_n507), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(G116), .B2(new_n258), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n251), .A2(new_n244), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n503), .B(new_n515), .C1(new_n287), .C2(new_n502), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n271), .A2(new_n500), .A3(new_n501), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G179), .A3(new_n514), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n327), .B1(new_n512), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n502), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(KEYINPUT21), .A3(new_n502), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n516), .A2(new_n518), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n251), .A2(new_n505), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n258), .A2(G97), .ZN(new_n527));
  INV_X1    g0327(.A(new_n377), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n398), .B2(new_n399), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n505), .A2(new_n217), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n204), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n352), .A2(new_n211), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n526), .B(new_n527), .C1(new_n537), .C2(new_n317), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G1698), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(G244), .C1(new_n276), .C2(new_n275), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n212), .B1(new_n296), .B2(new_n297), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n504), .C1(new_n543), .C2(KEYINPUT4), .ZN(new_n544));
  OAI21_X1  g0344(.A(G250), .B1(new_n275), .B2(new_n276), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n273), .B1(new_n545), .B2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n280), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n282), .A2(G257), .A3(new_n269), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n271), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n282), .A2(G257), .A3(new_n269), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n282), .A2(new_n337), .A3(new_n280), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(G190), .A3(new_n547), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n539), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(KEYINPUT78), .A3(new_n427), .A4(new_n547), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n547), .A2(new_n271), .A3(new_n427), .A4(new_n548), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT78), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n549), .A2(new_n327), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n538), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n204), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT79), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n298), .A2(new_n564), .A3(new_n204), .A4(G68), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n204), .B1(new_n461), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n505), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n377), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n566), .B1(new_n356), .B2(new_n505), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n563), .A2(new_n565), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n315), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n385), .A2(new_n251), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n216), .A2(new_n273), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n212), .A2(G1698), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n275), .C2(new_n276), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n269), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G45), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n272), .B1(new_n580), .B2(G1), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n203), .A2(new_n337), .A3(G45), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n269), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(G200), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n258), .A2(G87), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n573), .A2(new_n574), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n579), .A2(new_n584), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G190), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n572), .A2(new_n315), .B1(new_n251), .B2(new_n385), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(KEYINPUT80), .A3(new_n585), .A4(new_n586), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n258), .A2(new_n384), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n592), .A2(new_n595), .B1(new_n427), .B2(new_n590), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G169), .B2(new_n590), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n555), .A2(new_n561), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n331), .A2(new_n497), .A3(new_n525), .A4(new_n599), .ZN(G372));
  AND3_X1   g0400(.A1(new_n522), .A2(new_n518), .A3(new_n523), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n326), .B2(new_n329), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n573), .A2(new_n574), .A3(new_n586), .ZN(new_n603));
  INV_X1    g0403(.A(new_n579), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n269), .A2(new_n581), .A3(new_n582), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(G200), .B1(new_n590), .B2(G190), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n555), .A2(new_n561), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n602), .A2(new_n319), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n579), .B1(new_n605), .B2(new_n607), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT83), .B1(new_n614), .B2(G169), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n609), .A2(new_n616), .A3(new_n327), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n596), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n561), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n596), .A2(new_n618), .B1(new_n603), .B2(new_n610), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n594), .A2(new_n597), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT26), .B1(new_n624), .B2(new_n561), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n613), .A2(new_n619), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n497), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n374), .ZN(new_n628));
  INV_X1    g0428(.A(new_n491), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n495), .A2(new_n629), .B1(new_n476), .B2(new_n487), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n451), .A2(new_n456), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT18), .B1(new_n417), .B2(new_n436), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n438), .B(new_n435), .C1(new_n414), .C2(new_n416), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n371), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(new_n635), .ZN(G369));
  INV_X1    g0436(.A(G13), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(G20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n203), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT27), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(G213), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n326), .A2(new_n329), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n326), .A2(new_n647), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n330), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(KEYINPUT85), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n648), .A2(KEYINPUT85), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT86), .ZN(new_n654));
  INV_X1    g0454(.A(new_n601), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n647), .A2(new_n515), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n524), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G330), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n601), .A2(new_n646), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n326), .A2(new_n329), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n647), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n207), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G1), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n377), .A2(G116), .A3(new_n569), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(new_n230), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n556), .A2(new_n559), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n560), .A2(new_n538), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n622), .A2(new_n674), .A3(KEYINPUT26), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n621), .B1(new_n624), .B2(new_n561), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n620), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n622), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n613), .A3(new_n619), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n647), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n626), .A2(new_n647), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(KEYINPUT29), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n549), .A2(new_n284), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT88), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n517), .A2(G179), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n549), .A2(KEYINPUT88), .A3(new_n284), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n689), .A2(new_n609), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n590), .A2(new_n281), .A3(new_n283), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n517), .A3(G179), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n553), .B(new_n547), .C1(KEYINPUT87), .C2(new_n694), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n549), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n271), .A2(G179), .A3(new_n500), .A4(new_n501), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(KEYINPUT87), .B2(new_n694), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n702), .A3(KEYINPUT30), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n692), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(new_n705), .A3(new_n646), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n704), .B2(new_n646), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n330), .A2(new_n598), .A3(new_n524), .A4(new_n646), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n686), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n673), .B1(new_n713), .B2(G1), .ZN(G364));
  AOI21_X1  g0514(.A(new_n670), .B1(G45), .B2(new_n638), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n660), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(G330), .B2(new_n658), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n228), .B1(G20), .B2(new_n327), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n427), .A2(new_n285), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n287), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n204), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G97), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n204), .A2(new_n287), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n427), .A2(new_n285), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G50), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n720), .A2(new_n204), .A3(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G159), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT32), .Z(new_n734));
  NOR2_X1   g0534(.A1(new_n204), .A2(G190), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G68), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n726), .A2(new_n731), .A3(new_n734), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n427), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n735), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n211), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n727), .A2(new_n740), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G58), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n285), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n727), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G87), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n751), .A2(new_n735), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n298), .C1(new_n217), .C2(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n739), .A2(new_n742), .A3(new_n750), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n275), .A2(new_n276), .ZN(new_n761));
  INV_X1    g0561(.A(G303), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n755), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  INV_X1    g0564(.A(new_n741), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n732), .A2(G329), .B1(G311), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n758), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n730), .A2(G326), .B1(new_n767), .B2(G283), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n737), .A2(new_n769), .ZN(new_n770));
  AND3_X1   g0570(.A1(new_n766), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n764), .B(new_n771), .C1(new_n772), .C2(new_n722), .ZN(new_n773));
  INV_X1    g0573(.A(new_n748), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(G322), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n718), .B1(new_n760), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n667), .A2(new_n761), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G355), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n248), .A2(G45), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT90), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n667), .A2(new_n298), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G45), .B2(new_n230), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n778), .B1(G116), .B2(new_n207), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n718), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n776), .A2(new_n715), .A3(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT96), .Z(new_n790));
  INV_X1    g0590(.A(new_n786), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n658), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n717), .B1(new_n790), .B2(new_n792), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n646), .A2(new_n389), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n390), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n491), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n629), .A2(new_n647), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n685), .B(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(new_n712), .ZN(new_n800));
  INV_X1    g0600(.A(new_n715), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n755), .A2(new_n221), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G137), .A2(new_n730), .B1(new_n737), .B2(G150), .ZN(new_n804));
  INV_X1    g0604(.A(G143), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n410), .B2(new_n741), .C1(new_n748), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT34), .ZN(new_n807));
  INV_X1    g0607(.A(new_n722), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n761), .B1(new_n808), .B2(G58), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n215), .C2(new_n758), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n803), .B(new_n810), .C1(G132), .C2(new_n732), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n761), .B1(new_n748), .B2(new_n772), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n730), .A2(G303), .B1(new_n765), .B2(G116), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n736), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT97), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n756), .A2(G107), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n816), .A2(KEYINPUT97), .B1(G311), .B2(new_n732), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n726), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n812), .B(new_n820), .C1(G87), .C2(new_n767), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n718), .B1(new_n811), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n718), .A2(new_n784), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n211), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n798), .A2(new_n784), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n822), .A2(new_n715), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n802), .A2(new_n826), .ZN(G384));
  NAND2_X1  g0627(.A1(new_n404), .A2(new_n315), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT7), .B1(new_n761), .B2(new_n204), .ZN(new_n829));
  INV_X1    g0629(.A(new_n399), .ZN(new_n830));
  OAI21_X1  g0630(.A(G68), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n402), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n412), .A2(KEYINPUT72), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT16), .B1(new_n834), .B2(new_n395), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n416), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n644), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT102), .B1(new_n457), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT102), .ZN(new_n840));
  INV_X1    g0640(.A(new_n838), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n632), .A2(new_n633), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(new_n841), .C1(new_n631), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  AND4_X1   g0644(.A1(new_n414), .A2(new_n416), .A3(new_n449), .A4(new_n445), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n414), .A2(new_n416), .B1(new_n435), .B2(new_n644), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n836), .A2(new_n436), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n838), .A2(new_n848), .A3(new_n450), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(KEYINPUT37), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n853), .B(new_n850), .C1(new_n839), .C2(new_n843), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT99), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n476), .A2(new_n487), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n476), .B2(new_n487), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n646), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(new_n846), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n845), .A2(new_n846), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n417), .A2(new_n837), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n457), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n853), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT39), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  OR3_X1    g0673(.A1(new_n856), .A2(new_n862), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n797), .B1(new_n685), .B2(new_n798), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n486), .A2(new_n647), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n495), .B(new_n877), .C1(new_n858), .C2(new_n859), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n476), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT100), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(new_n476), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n875), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n886), .B(new_n888), .C1(new_n854), .C2(new_n852), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n842), .A2(new_n644), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n874), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n686), .A2(new_n497), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n635), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n891), .B(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n865), .A2(new_n450), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n867), .B(new_n897), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n457), .A2(new_n870), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT105), .B1(new_n854), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT104), .B1(new_n708), .B2(new_n709), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n798), .B1(new_n878), .B2(new_n883), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n331), .A2(new_n525), .A3(new_n599), .A4(new_n647), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n904), .B(new_n905), .C1(new_n707), .C2(new_n706), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n863), .A2(new_n909), .A3(new_n872), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n901), .A2(new_n908), .A3(new_n910), .A4(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n852), .A2(new_n854), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(new_n907), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n497), .A2(new_n902), .A3(new_n906), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n915), .B(new_n916), .Z(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n711), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n896), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n894), .B(KEYINPUT106), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n919), .B1(new_n203), .B2(new_n638), .C1(new_n920), .C2(new_n918), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n533), .A2(new_n534), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n244), .B1(new_n922), .B2(KEYINPUT35), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n229), .C1(KEYINPUT35), .C2(new_n922), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n393), .A2(G77), .A3(new_n231), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT98), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(G50), .B2(new_n215), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n637), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n925), .A3(new_n929), .ZN(G367));
  OAI211_X1 g0730(.A(new_n555), .B(new_n561), .C1(new_n539), .C2(new_n647), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n620), .A2(new_n646), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n663), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n933), .B(KEYINPUT108), .Z(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n664), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n647), .B1(new_n938), .B2(new_n620), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT43), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n647), .A2(new_n603), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n619), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n622), .B2(new_n942), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT107), .Z(new_n945));
  OAI21_X1  g0745(.A(new_n940), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n654), .A2(new_n660), .A3(new_n937), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  INV_X1    g0749(.A(new_n945), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n948), .B2(new_n949), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n668), .B(KEYINPUT41), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n663), .A2(new_n665), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT109), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(new_n934), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n957), .B2(new_n934), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n957), .A2(new_n934), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n660), .A3(new_n654), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n963), .A2(new_n661), .A3(new_n965), .A4(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n654), .B(new_n662), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n660), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(new_n713), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n956), .B1(new_n973), .B2(new_n713), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n638), .A2(G45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(G1), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n953), .B(new_n954), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n781), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n787), .B1(new_n207), .B2(new_n385), .C1(new_n240), .C2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT110), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n725), .A2(G68), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n761), .B1(new_n765), .B2(G50), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n410), .B2(new_n736), .C1(new_n755), .C2(new_n749), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G150), .B2(new_n774), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n211), .B2(new_n758), .C1(new_n805), .C2(new_n729), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n982), .B(new_n986), .C1(G137), .C2(new_n732), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n755), .A2(new_n244), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT46), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n298), .B1(new_n774), .B2(G303), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT111), .B(G311), .Z(new_n991));
  AOI22_X1  g0791(.A1(new_n730), .A2(new_n991), .B1(new_n765), .B2(G283), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n732), .A2(G317), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G294), .A2(new_n737), .B1(new_n767), .B2(G97), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n990), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n989), .B(new_n995), .C1(new_n377), .C2(new_n808), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n987), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  AOI21_X1  g0798(.A(new_n980), .B1(new_n998), .B2(new_n718), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n715), .C1(new_n791), .C2(new_n950), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n977), .A2(new_n1000), .ZN(G387));
  NOR2_X1   g0801(.A1(new_n972), .A2(new_n669), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n713), .B2(new_n971), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n971), .A2(new_n976), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n978), .B1(new_n237), .B2(G45), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n671), .B2(new_n777), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n415), .A2(new_n221), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n215), .A2(new_n211), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1008), .A2(G45), .A3(new_n1009), .A4(new_n671), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1006), .A2(new_n1010), .B1(G107), .B2(new_n207), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n801), .B1(new_n1011), .B2(new_n787), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n725), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n385), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n732), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1016), .A2(new_n350), .B1(new_n755), .B2(new_n211), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n767), .A2(G97), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n774), .A2(G50), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n298), .B1(new_n736), .B2(new_n355), .C1(new_n410), .C2(new_n729), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G68), .B2(new_n765), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n774), .A2(G317), .B1(G303), .B2(new_n765), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n730), .A2(G322), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n737), .A2(new_n991), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n814), .B2(new_n722), .C1(new_n772), .C2(new_n755), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT49), .Z(new_n1030));
  NAND2_X1  g0830(.A1(new_n732), .A2(G326), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n761), .C1(new_n244), .C2(new_n758), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1023), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT113), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n718), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1013), .B1(new_n654), .B2(new_n791), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1003), .A2(new_n1004), .A3(new_n1036), .ZN(G393));
  NAND3_X1  g0837(.A1(new_n968), .A2(new_n976), .A3(new_n969), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n774), .A2(G311), .B1(G317), .B2(new_n730), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G303), .B2(new_n737), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n732), .A2(G322), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n808), .A2(G116), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n217), .A2(new_n758), .B1(new_n741), .B2(new_n772), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n298), .B(new_n1044), .C1(new_n756), .C2(G283), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1014), .A2(new_n211), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n732), .A2(G143), .B1(G87), .B2(new_n767), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n298), .C1(new_n215), .C2(new_n755), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT115), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n748), .A2(new_n410), .B1(new_n350), .B2(new_n729), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT51), .Z(new_n1052));
  NOR2_X1   g0852(.A1(new_n736), .A2(new_n221), .ZN(new_n1053));
  OR4_X1    g0853(.A1(new_n1047), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n741), .A2(new_n355), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1046), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n718), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n245), .A2(new_n781), .B1(G97), .B2(new_n667), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n787), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n715), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT114), .Z(new_n1061));
  OAI211_X1 g0861(.A(new_n1057), .B(new_n1061), .C1(new_n937), .C2(new_n791), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n973), .A2(new_n668), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n972), .B1(new_n968), .B2(new_n969), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1038), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(G390));
  NAND3_X1  g0865(.A1(new_n682), .A2(new_n647), .A3(new_n796), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n797), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n861), .B1(new_n1067), .B2(new_n884), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1068), .A2(new_n901), .A3(new_n910), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT116), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n885), .A2(new_n862), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n856), .B2(new_n873), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n901), .A3(new_n910), .A4(KEYINPUT116), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n908), .A2(G330), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n798), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n712), .A2(new_n1078), .A3(new_n884), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n710), .A2(new_n711), .A3(new_n798), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n884), .A2(new_n1083), .B1(new_n907), .B2(new_n711), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n875), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n902), .A2(new_n1086), .A3(G330), .A4(new_n906), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1087), .A2(new_n1078), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n902), .A2(G330), .A3(new_n906), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT117), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n884), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1079), .A2(new_n797), .A3(new_n1066), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1091), .A2(KEYINPUT118), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT118), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n884), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1090), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1087), .A2(new_n1078), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1092), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1085), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n916), .A2(G330), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n893), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1082), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1085), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT118), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1098), .A2(new_n1099), .A3(new_n1094), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1103), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1077), .B(new_n1081), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1110), .A3(new_n668), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n784), .B1(new_n856), .B2(new_n873), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n528), .A2(new_n736), .B1(new_n741), .B2(new_n505), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT119), .Z(new_n1114));
  NOR2_X1   g0914(.A1(new_n1016), .A2(new_n772), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1115), .B(new_n1047), .C1(G116), .C2(new_n774), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n730), .A2(G283), .B1(new_n767), .B2(G68), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n757), .A2(new_n761), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT120), .Z(new_n1119));
  AND4_X1   g0919(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n725), .A2(G159), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n737), .A2(G137), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n755), .A2(new_n350), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT54), .B(G143), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n765), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(G128), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n729), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G132), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n748), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n761), .B1(new_n732), .B2(G125), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n221), .B2(new_n758), .ZN(new_n1133));
  NOR4_X1   g0933(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n718), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1112), .A2(new_n715), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n355), .B2(new_n823), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1082), .B2(new_n976), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1111), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT121), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1111), .A2(new_n1141), .A3(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(G378));
  NAND3_X1  g0943(.A1(new_n911), .A2(new_n914), .A3(G330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n371), .A2(new_n374), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1146));
  OR2_X1    g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n837), .A2(new_n366), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1147), .A2(new_n366), .A3(new_n837), .A4(new_n1148), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1144), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1155), .A2(new_n914), .A3(new_n911), .A4(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n891), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n874), .A2(new_n890), .A3(new_n889), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n976), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1153), .A2(new_n785), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n981), .B1(new_n244), .B2(new_n729), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT122), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n761), .B1(new_n748), .B2(new_n217), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n260), .B1(new_n755), .B2(new_n211), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n385), .A2(new_n741), .B1(new_n505), .B2(new_n736), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n749), .B2(new_n758), .C1(new_n814), .C2(new_n1016), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT58), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n221), .B1(new_n275), .B2(G41), .ZN(new_n1173));
  INV_X1    g0973(.A(G124), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n260), .B1(new_n1016), .B2(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n725), .A2(G150), .B1(G128), .B2(new_n774), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n756), .A2(new_n1125), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G125), .A2(new_n730), .B1(new_n737), .B2(G132), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G137), .B2(new_n765), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT59), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(new_n1175), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .C1(new_n410), .C2(new_n758), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1172), .A2(new_n1173), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n718), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n823), .A2(new_n221), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1164), .A2(new_n1185), .A3(new_n715), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1162), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1109), .B1(new_n1082), .B2(new_n1101), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n669), .B1(new_n1191), .B2(KEYINPUT57), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1188), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G375));
  NOR2_X1   g0996(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n955), .A3(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n528), .A2(new_n741), .B1(new_n758), .B2(new_n211), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n736), .A2(new_n244), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1015), .A2(new_n298), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n774), .A2(G283), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1016), .A2(new_n762), .B1(new_n755), .B2(new_n505), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT123), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n730), .A2(G294), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n774), .A2(G137), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n761), .B1(new_n737), .B2(new_n1125), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n1130), .B2(new_n729), .C1(new_n1016), .C2(new_n1128), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n725), .B2(G50), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G58), .A2(new_n767), .B1(new_n765), .B2(G150), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n410), .C2(new_n755), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1208), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT124), .Z(new_n1216));
  OAI221_X1 g1016(.A(new_n715), .B1(new_n785), .B2(new_n884), .C1(new_n1216), .C2(new_n1035), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n215), .B2(new_n823), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1101), .B2(new_n976), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1200), .A2(new_n1219), .ZN(G381));
  INV_X1    g1020(.A(G390), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n977), .A3(new_n1000), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1222), .A2(G396), .A3(G393), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G375), .A2(new_n1139), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G384), .A3(G381), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(G407));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G343), .C2(new_n1225), .ZN(G409));
  INV_X1    g1028(.A(new_n1188), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1191), .A2(new_n955), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1139), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1103), .B1(new_n1234), .B2(new_n1108), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(KEYINPUT57), .A3(new_n1161), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n668), .A3(new_n1194), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1111), .A2(new_n1141), .A3(new_n1138), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1141), .B1(new_n1111), .B2(new_n1138), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1237), .B(new_n1229), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1195), .B2(G378), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1233), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n669), .B1(new_n1197), .B2(KEYINPUT60), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n1199), .C1(KEYINPUT60), .C2(new_n1197), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1246), .A2(G384), .A3(new_n1219), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G384), .B1(new_n1246), .B2(new_n1219), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(G213), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(G343), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1244), .A2(new_n1249), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1195), .A2(G378), .A3(new_n1242), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1251), .B1(new_n1256), .B2(new_n1233), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1249), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(G2897), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1249), .A2(G2897), .A3(new_n1251), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1257), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1253), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1254), .A2(new_n1255), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1251), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1266), .A2(new_n1265), .A3(new_n1251), .ZN(new_n1269));
  OAI211_X1 g1069(.A(KEYINPUT63), .B(new_n1249), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(G390), .ZN(new_n1272));
  XOR2_X1   g1072(.A(G393), .B(G396), .Z(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1272), .A2(new_n1222), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1272), .B2(new_n1222), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1264), .A2(new_n1270), .A3(new_n1271), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1267), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1271), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1283), .B(KEYINPUT62), .C1(new_n1257), .C2(new_n1249), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(KEYINPUT62), .B(new_n1249), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1282), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1278), .B1(new_n1289), .B2(new_n1277), .ZN(G405));
  AOI22_X1  g1090(.A1(new_n1254), .A2(new_n1255), .B1(new_n1232), .B2(G375), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1277), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1258), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1249), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


