//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206));
  INV_X1    g005(.A(G85gat), .ZN(new_n207));
  INV_X1    g006(.A(G92gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(KEYINPUT8), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT93), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n212), .A3(new_n209), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G99gat), .B(G106gat), .Z(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n215), .A3(new_n213), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G71gat), .B(G78gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT88), .ZN(new_n222));
  AND2_X1   g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT9), .ZN(new_n224));
  INV_X1    g023(.A(G57gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G64gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n225), .A2(G64gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(KEYINPUT89), .B2(new_n226), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(KEYINPUT89), .B2(new_n226), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n224), .A3(new_n221), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT90), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n233), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n202), .B1(new_n220), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n234), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n219), .A2(KEYINPUT94), .A3(new_n238), .A4(new_n235), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G230gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT95), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT95), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n248), .A3(new_n245), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(KEYINPUT96), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT10), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n240), .A2(new_n251), .A3(new_n241), .A4(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n239), .A3(KEYINPUT10), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n245), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G176gat), .B(G204gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT96), .B1(new_n247), .B2(new_n249), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT97), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n249), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT96), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT97), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n250), .A4(new_n259), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n258), .B1(new_n263), .B2(new_n254), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n239), .A2(KEYINPUT21), .ZN(new_n271));
  XOR2_X1   g070(.A(G127gat), .B(G155gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G8gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n275), .A2(G1gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n276), .B2(KEYINPUT84), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT16), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(G1gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n277), .B(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(new_n239), .B2(KEYINPUT21), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n273), .B(new_n282), .Z(new_n283));
  NAND2_X1  g082(.A1(G231gat), .A2(G233gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT91), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G183gat), .B(G211gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n283), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G29gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n297), .B2(G36gat), .ZN(new_n298));
  INV_X1    g097(.A(G50gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G43gat), .ZN(new_n300));
  INV_X1    g099(.A(G43gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G50gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT15), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT83), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT15), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n306), .B(new_n307), .C1(new_n305), .C2(new_n302), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n308), .A2(new_n298), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n304), .B1(new_n309), .B2(new_n303), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n310), .A2(KEYINPUT17), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(KEYINPUT17), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n219), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n313), .B(new_n314), .C1(new_n310), .C2(new_n219), .ZN(new_n315));
  XOR2_X1   g114(.A(G190gat), .B(G218gat), .Z(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  XNOR2_X1  g116(.A(G134gat), .B(G162gat), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n317), .A2(new_n320), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n292), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n270), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT98), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n270), .A2(new_n325), .A3(KEYINPUT98), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n281), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n311), .A2(new_n332), .A3(new_n312), .ZN(new_n333));
  INV_X1    g132(.A(new_n310), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n281), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(KEYINPUT85), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n334), .B2(new_n281), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n331), .B(new_n333), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n331), .B(KEYINPUT13), .Z(new_n341));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n334), .B2(new_n281), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n332), .A2(KEYINPUT86), .A3(new_n310), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(new_n344), .C1(new_n336), .C2(new_n338), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n340), .A2(KEYINPUT18), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G141gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(G197gat), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT11), .B(G169gat), .Z(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n350), .B(KEYINPUT12), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT18), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n354), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT87), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n346), .A2(new_n352), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n336), .A2(new_n338), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n359), .A2(KEYINPUT18), .A3(new_n331), .A4(new_n333), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n341), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n351), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366));
  AND2_X1   g165(.A1(G113gat), .A2(G120gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(G113gat), .A2(G120gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(G127gat), .A2(G134gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(G127gat), .A2(G134gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT69), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n366), .B(new_n369), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G113gat), .ZN(new_n375));
  INV_X1    g174(.A(G120gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G113gat), .A2(G120gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n366), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n373), .A3(new_n378), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G141gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G148gat), .ZN(new_n385));
  INV_X1    g184(.A(G148gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G141gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT2), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n392), .A2(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G155gat), .B(G162gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n395), .A3(new_n390), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n383), .A2(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n388), .A2(new_n395), .A3(new_n390), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n395), .B1(new_n390), .B2(new_n388), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n374), .A2(new_n382), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT4), .B1(new_n401), .B2(new_n402), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n374), .A2(new_n382), .A3(KEYINPUT70), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT70), .B1(new_n374), .B2(new_n382), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n410), .A2(new_n411), .A3(new_n397), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n406), .B(new_n409), .C1(new_n412), .C2(KEYINPUT4), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT74), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n415), .B(KEYINPUT3), .C1(new_n399), .C2(new_n400), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n394), .A2(new_n417), .A3(new_n396), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n383), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT74), .B1(new_n401), .B2(new_n417), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n402), .B1(new_n401), .B2(new_n417), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT75), .A4(new_n416), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n408), .B1(new_n413), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n411), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n374), .A2(new_n382), .A3(KEYINPUT70), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n401), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n406), .A2(KEYINPUT5), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT76), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n425), .A2(KEYINPUT76), .A3(new_n433), .A4(new_n434), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n426), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G1gat), .B(G29gat), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(G57gat), .B(G85gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT6), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n426), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n427), .B1(new_n412), .B2(KEYINPUT4), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n421), .B2(new_n424), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT76), .B1(new_n447), .B2(new_n434), .ZN(new_n448));
  INV_X1    g247(.A(new_n438), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n443), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n454), .B2(new_n445), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G197gat), .B(G204gat), .ZN(new_n458));
  INV_X1    g257(.A(G211gat), .ZN(new_n459));
  INV_X1    g258(.A(G218gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n458), .B1(KEYINPUT22), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G211gat), .B(G218gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT65), .B(G183gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT66), .B(G190gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(G183gat), .A2(G190gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT24), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT24), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(G183gat), .A3(G190gat), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n467), .A2(new_n468), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G169gat), .ZN(new_n474));
  INV_X1    g273(.A(G176gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT23), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT23), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(G169gat), .B2(G176gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(G169gat), .A2(G176gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT25), .A4(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n466), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n470), .A2(new_n472), .ZN(new_n482));
  INV_X1    g281(.A(G183gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT65), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G183gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G190gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT66), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G190gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n482), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n480), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT67), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n470), .A2(new_n472), .B1(new_n483), .B2(new_n488), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT26), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT26), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(G169gat), .B2(G176gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n479), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n501), .B(new_n469), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(G169gat), .A2(G176gat), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n508), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(KEYINPUT68), .C1(new_n504), .C2(new_n503), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT27), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n467), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT28), .B1(new_n515), .B2(new_n468), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G183gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n468), .A2(new_n517), .A3(KEYINPUT28), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n511), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n500), .A2(new_n520), .A3(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n481), .A2(new_n495), .A3(new_n499), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n512), .B1(new_n487), .B2(KEYINPUT27), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(new_n492), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n532), .A2(new_n518), .B1(new_n507), .B2(new_n510), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n528), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n500), .A2(new_n520), .A3(KEYINPUT73), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT29), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n465), .B(new_n527), .C1(new_n536), .C2(new_n526), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n526), .A3(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n524), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n538), .B(new_n464), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G8gat), .B(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G64gat), .B(G92gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n537), .A2(new_n542), .ZN(new_n549));
  INV_X1    g348(.A(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n537), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n545), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n457), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n417), .B1(new_n464), .B2(KEYINPUT29), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n418), .A2(new_n540), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n556), .A2(new_n397), .B1(new_n464), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G78gat), .B(G106gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G228gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G22gat), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G50gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n560), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI22_X1  g365(.A1(new_n529), .A2(new_n533), .B1(new_n410), .B2(new_n411), .ZN(new_n567));
  INV_X1    g366(.A(G227gat), .ZN(new_n568));
  INV_X1    g367(.A(G233gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n500), .A2(new_n520), .A3(new_n430), .A4(new_n429), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT34), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G15gat), .B(G43gat), .Z(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G99gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n570), .B(KEYINPUT64), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n567), .B2(new_n572), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n582), .B2(KEYINPUT33), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n580), .A2(KEYINPUT34), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n572), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n585), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n576), .A2(new_n586), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT71), .B1(new_n573), .B2(KEYINPUT34), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n589), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n583), .A2(new_n585), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n596), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n555), .A2(new_n566), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n537), .A2(new_n603), .A3(new_n542), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n550), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n537), .B2(new_n542), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT38), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n443), .B(KEYINPUT77), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n450), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n444), .A2(new_n611), .B1(KEYINPUT6), .B2(new_n455), .ZN(new_n612));
  INV_X1    g411(.A(new_n546), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n604), .A2(new_n614), .A3(new_n550), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT79), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n534), .A2(new_n535), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n526), .B1(new_n617), .B2(new_n540), .ZN(new_n618));
  INV_X1    g417(.A(new_n527), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n616), .B(new_n464), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n524), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT72), .B1(new_n500), .B2(new_n520), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n621), .A2(new_n622), .A3(new_n541), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n500), .A2(new_n520), .A3(KEYINPUT73), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT73), .B1(new_n500), .B2(new_n520), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n624), .A2(new_n625), .A3(new_n525), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n465), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT79), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n540), .B1(new_n624), .B2(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n525), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n465), .B1(new_n630), .B2(new_n527), .ZN(new_n631));
  OAI211_X1 g430(.A(KEYINPUT37), .B(new_n620), .C1(new_n628), .C2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n613), .B1(new_n615), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(KEYINPUT80), .B(KEYINPUT38), .C1(new_n605), .C2(new_n606), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n609), .A2(new_n612), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n405), .B1(new_n425), .B2(new_n433), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n610), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT78), .ZN(new_n640));
  INV_X1    g439(.A(new_n404), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n637), .B1(new_n641), .B2(new_n405), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n447), .B2(new_n405), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n638), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n610), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n454), .B2(new_n445), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n638), .B2(new_n643), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n566), .B1(new_n648), .B2(new_n553), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n635), .A2(KEYINPUT81), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT81), .B1(new_n635), .B2(new_n649), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n602), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n590), .A2(new_n596), .A3(new_n565), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n443), .B(new_n445), .C1(new_n448), .C2(new_n449), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT6), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n654), .B(new_n655), .C1(new_n439), .C2(new_n645), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n456), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT35), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .A4(new_n554), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT82), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n599), .A2(new_n566), .A3(new_n553), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n662), .A2(KEYINPUT82), .A3(new_n658), .A4(new_n657), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n457), .A3(new_n554), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT35), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n365), .B1(new_n652), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n330), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n457), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT100), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT99), .B(G1gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1324gat));
  NAND3_X1  g471(.A1(new_n330), .A2(new_n553), .A3(new_n667), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT16), .B(G8gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n675), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n673), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n675), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(G1325gat));
  NAND2_X1  g481(.A1(new_n598), .A2(new_n601), .ZN(new_n683));
  OAI21_X1  g482(.A(G15gat), .B1(new_n668), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n599), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n668), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n668), .A2(new_n565), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n555), .A2(new_n566), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n683), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n609), .A2(new_n634), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n615), .A2(new_n632), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n693), .A2(new_n456), .A3(new_n656), .A4(new_n546), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n649), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT81), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n635), .A2(KEYINPUT81), .A3(new_n649), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n323), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n652), .A2(new_n666), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(KEYINPUT44), .A3(new_n323), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n358), .A2(new_n363), .A3(KEYINPUT103), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT103), .B1(new_n358), .B2(new_n363), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n292), .ZN(new_n711));
  INV_X1    g510(.A(new_n269), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n262), .B2(new_n267), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n706), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n457), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n324), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n667), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(G29gat), .A3(new_n457), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(new_n722), .ZN(G1328gat));
  OAI21_X1  g522(.A(G36gat), .B1(new_n716), .B2(new_n554), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n719), .A2(G36gat), .A3(new_n554), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1329gat));
  NAND4_X1  g526(.A1(new_n667), .A2(new_n301), .A3(new_n597), .A4(new_n718), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(KEYINPUT47), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n716), .B2(new_n683), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G43gat), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n716), .A2(KEYINPUT104), .A3(new_n683), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n683), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n715), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n728), .B1(new_n735), .B2(new_n301), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n738), .ZN(G1330gat));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n565), .A2(G50gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n719), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n667), .B2(new_n718), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n714), .A2(new_n710), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n703), .A2(new_n566), .A3(new_n705), .A4(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G50gat), .B1(new_n747), .B2(new_n748), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT48), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n747), .A2(new_n754), .A3(G50gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n747), .B2(G50gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n743), .B2(new_n744), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n740), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT44), .B1(new_n704), .B2(new_n323), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n702), .B(new_n324), .C1(new_n652), .C2(new_n666), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(KEYINPUT107), .A3(new_n566), .A4(new_n746), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n749), .A3(G50gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n757), .B1(new_n765), .B2(new_n745), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT108), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n760), .A2(new_n768), .ZN(G1331gat));
  NOR3_X1   g568(.A1(new_n325), .A2(new_n713), .A3(new_n709), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n704), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n457), .B(KEYINPUT109), .Z(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n553), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT49), .B(G64gat), .Z(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n771), .A2(G71gat), .A3(new_n734), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n599), .B(KEYINPUT110), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(G71gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n566), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT112), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT111), .B(G78gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  NOR3_X1   g586(.A1(new_n713), .A2(new_n709), .A3(new_n292), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n763), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n457), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n292), .A2(new_n709), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n704), .A2(new_n323), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT51), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n270), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n457), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n207), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n791), .B1(new_n797), .B2(new_n799), .ZN(G1336gat));
  NAND2_X1  g599(.A1(new_n789), .A2(new_n553), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n793), .B(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n713), .A2(G92gat), .A3(new_n554), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n805), .B(KEYINPUT114), .Z(new_n808));
  AOI22_X1  g607(.A1(new_n801), .A2(G92gat), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n790), .B2(new_n683), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n599), .A2(G99gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n797), .B2(new_n813), .ZN(G1338gat));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n703), .A2(new_n566), .A3(new_n705), .A4(new_n788), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n713), .A2(G106gat), .A3(new_n565), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n818), .A2(KEYINPUT115), .B1(new_n804), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n821), .A3(G106gat), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  INV_X1    g623(.A(new_n819), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n794), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n804), .A2(KEYINPUT116), .A3(new_n819), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT53), .B1(new_n817), .B2(G106gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n815), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n804), .A2(new_n819), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n832), .A2(new_n833), .A3(new_n822), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT117), .B(new_n829), .C1(new_n834), .C2(new_n816), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(G1339gat));
  NAND2_X1  g635(.A1(new_n326), .A2(new_n710), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n252), .A2(new_n253), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n244), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n252), .A2(new_n245), .A3(new_n253), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n257), .B1(new_n254), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT55), .B1(new_n841), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n268), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n331), .B1(new_n359), .B2(new_n333), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n345), .A2(new_n341), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n350), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n358), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(KEYINPUT118), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n323), .B1(new_n854), .B2(new_n851), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n847), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n847), .A2(new_n710), .B1(new_n713), .B2(new_n851), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n324), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n837), .B1(new_n858), .B2(new_n292), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n798), .A2(new_n554), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n599), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n565), .A3(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n375), .A3(new_n365), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n859), .A2(new_n772), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n662), .A3(new_n709), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n375), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n862), .B2(new_n713), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n662), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n713), .A2(G120gat), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT119), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n868), .B2(new_n870), .ZN(G1341gat));
  OR3_X1    g670(.A1(new_n868), .A2(G127gat), .A3(new_n711), .ZN(new_n872));
  OAI21_X1  g671(.A(G127gat), .B1(new_n862), .B2(new_n711), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(KEYINPUT120), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1342gat));
  OR2_X1    g677(.A1(new_n324), .A2(G134gat), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n868), .A2(KEYINPUT56), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n862), .B2(new_n324), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT56), .B1(new_n868), .B2(new_n879), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n268), .A2(new_n709), .A3(new_n846), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n713), .A2(new_n851), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n324), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n847), .A2(new_n853), .A3(new_n855), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n292), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n837), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n885), .B(new_n566), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n734), .A2(new_n860), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n270), .A2(new_n852), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n268), .A2(new_n364), .A3(new_n846), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n323), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n711), .B1(new_n896), .B2(new_n856), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n565), .B1(new_n897), .B2(new_n837), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n892), .B(new_n893), .C1(new_n898), .C2(new_n885), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n884), .B1(new_n899), .B2(new_n365), .ZN(new_n900));
  INV_X1    g699(.A(new_n893), .ZN(new_n901));
  INV_X1    g700(.A(new_n895), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n324), .B1(new_n902), .B2(new_n887), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n292), .B1(new_n903), .B2(new_n889), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n566), .B1(new_n904), .B2(new_n891), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(KEYINPUT123), .A3(new_n364), .A4(new_n892), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n900), .A2(new_n907), .A3(G141gat), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n734), .A2(new_n565), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n772), .B(new_n909), .C1(new_n890), .C2(new_n891), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n859), .A2(KEYINPUT122), .A3(new_n772), .A4(new_n909), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n365), .A2(G141gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n912), .A2(new_n913), .A3(new_n554), .A4(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NOR4_X1   g717(.A1(new_n910), .A2(G141gat), .A3(new_n365), .A4(new_n553), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT57), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n892), .A4(new_n893), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n923), .A3(new_n709), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n924), .B2(G141gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n918), .B1(new_n925), .B2(new_n916), .ZN(G1344gat));
  NAND3_X1  g725(.A1(new_n912), .A2(new_n913), .A3(new_n554), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n927), .A2(G148gat), .A3(new_n713), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n920), .A2(new_n923), .A3(new_n270), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n386), .A2(KEYINPUT59), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n890), .A2(new_n891), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT57), .B1(new_n932), .B2(new_n565), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n328), .A2(new_n364), .A3(new_n329), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n885), .B(new_n566), .C1(new_n934), .C2(new_n904), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n893), .A2(new_n270), .ZN(new_n937));
  OAI21_X1  g736(.A(G148gat), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(KEYINPUT59), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n928), .B1(new_n931), .B2(new_n939), .ZN(G1345gat));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n923), .ZN(new_n941));
  OAI21_X1  g740(.A(G155gat), .B1(new_n941), .B2(new_n711), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n711), .A2(G155gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n927), .B2(new_n943), .ZN(G1346gat));
  NOR2_X1   g743(.A1(new_n324), .A2(G162gat), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n912), .A2(new_n913), .A3(new_n554), .A4(new_n945), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT124), .Z(new_n947));
  OAI21_X1  g746(.A(G162gat), .B1(new_n941), .B2(new_n324), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n798), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n599), .A2(new_n554), .A3(new_n566), .ZN(new_n951));
  AND4_X1   g750(.A1(new_n474), .A2(new_n950), .A3(new_n709), .A4(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n772), .A2(new_n554), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(new_n780), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n859), .A2(new_n565), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n859), .A2(new_n959), .A3(new_n565), .A4(new_n956), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n958), .A2(new_n364), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n954), .B1(new_n474), .B2(new_n961), .ZN(G1348gat));
  NAND2_X1  g761(.A1(new_n950), .A2(new_n951), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n475), .A3(new_n270), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n958), .A2(new_n270), .A3(new_n960), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n475), .ZN(G1349gat));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n292), .A3(new_n960), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n487), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n517), .A3(new_n292), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n964), .A2(new_n468), .A3(new_n323), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n323), .A3(new_n960), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n977), .A2(new_n978), .A3(G190gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n977), .B2(G190gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  NOR3_X1   g780(.A1(new_n772), .A2(new_n554), .A3(new_n734), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n933), .A2(new_n935), .A3(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(G197gat), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n983), .A2(new_n984), .A3(new_n365), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n950), .A2(new_n553), .A3(new_n909), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n986), .A2(new_n710), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n985), .B1(new_n984), .B2(new_n987), .ZN(G1352gat));
  NOR3_X1   g787(.A1(new_n986), .A2(G204gat), .A3(new_n713), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(KEYINPUT127), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(G204gat), .B1(new_n983), .B2(new_n713), .ZN(new_n992));
  XNOR2_X1  g791(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n991), .B(new_n992), .C1(new_n989), .C2(new_n993), .ZN(G1353gat));
  NAND4_X1  g793(.A1(new_n933), .A2(new_n935), .A3(new_n292), .A4(new_n982), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n292), .A2(new_n459), .ZN(new_n998));
  OAI22_X1  g797(.A1(new_n996), .A2(new_n997), .B1(new_n986), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n983), .B2(new_n324), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n323), .A2(new_n460), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n986), .B2(new_n1001), .ZN(G1355gat));
endmodule


