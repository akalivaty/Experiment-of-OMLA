

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U549 ( .A(n547), .Z(n876) );
  NOR2_X2 U550 ( .A1(n977), .A2(n694), .ZN(n678) );
  NOR2_X1 U551 ( .A1(n745), .A2(n801), .ZN(n746) );
  NOR2_X1 U552 ( .A1(n682), .A2(n681), .ZN(n691) );
  INV_X1 U553 ( .A(KEYINPUT94), .ZN(n673) );
  XNOR2_X1 U554 ( .A(n709), .B(KEYINPUT30), .ZN(n711) );
  NOR2_X1 U555 ( .A1(n708), .A2(n733), .ZN(n709) );
  XNOR2_X1 U556 ( .A(n744), .B(n743), .ZN(n745) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n743) );
  NOR2_X1 U558 ( .A1(G651), .A2(n628), .ZN(n634) );
  XOR2_X1 U559 ( .A(KEYINPUT6), .B(n524), .Z(n513) );
  NOR2_X1 U560 ( .A1(n965), .A2(n806), .ZN(n514) );
  XNOR2_X1 U561 ( .A(n679), .B(KEYINPUT99), .ZN(n682) );
  INV_X1 U562 ( .A(G168), .ZN(n710) );
  AND2_X1 U563 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U564 ( .A1(n714), .A2(n713), .ZN(n715) );
  BUF_X1 U565 ( .A(n707), .Z(n722) );
  INV_X1 U566 ( .A(KEYINPUT101), .ZN(n720) );
  NOR2_X1 U567 ( .A1(G2084), .A2(n707), .ZN(n706) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  INV_X1 U569 ( .A(KEYINPUT105), .ZN(n752) );
  NOR2_X1 U570 ( .A1(n751), .A2(n750), .ZN(n753) );
  INV_X1 U571 ( .A(G651), .ZN(n519) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n643) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(n521), .ZN(n636) );
  XNOR2_X1 U574 ( .A(n526), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U575 ( .A1(n643), .A2(G89), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n515), .B(KEYINPUT4), .ZN(n517) );
  XOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NOR2_X1 U578 ( .A1(n628), .A2(n519), .ZN(n639) );
  NAND2_X1 U579 ( .A1(G76), .A2(n639), .ZN(n516) );
  NAND2_X1 U580 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(KEYINPUT5), .ZN(n525) );
  NAND2_X1 U582 ( .A1(G51), .A2(n634), .ZN(n523) );
  NOR2_X1 U583 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n520), .Z(n521) );
  NAND2_X1 U585 ( .A1(G63), .A2(n636), .ZN(n522) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n525), .A2(n513), .ZN(n526) );
  XNOR2_X2 U588 ( .A(G2104), .B(KEYINPUT65), .ZN(n534) );
  NOR2_X2 U589 ( .A1(G2105), .A2(n534), .ZN(n546) );
  NAND2_X1 U590 ( .A1(G101), .A2(n546), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT66), .B(n527), .ZN(n529) );
  INV_X1 U592 ( .A(KEYINPUT23), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT17), .B(n530), .Z(n547) );
  NAND2_X1 U595 ( .A1(G137), .A2(n876), .ZN(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n538) );
  NAND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT67), .ZN(n551) );
  BUF_X1 U599 ( .A(n551), .Z(n878) );
  NAND2_X1 U600 ( .A1(G113), .A2(n878), .ZN(n536) );
  AND2_X1 U601 ( .A1(n534), .A2(G2105), .ZN(n879) );
  NAND2_X1 U602 ( .A1(G125), .A2(n879), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X4 U604 ( .A1(n538), .A2(n537), .ZN(G160) );
  NAND2_X1 U605 ( .A1(G53), .A2(n634), .ZN(n540) );
  NAND2_X1 U606 ( .A1(G65), .A2(n636), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT72), .B(n541), .Z(n545) );
  NAND2_X1 U609 ( .A1(n639), .A2(G78), .ZN(n543) );
  NAND2_X1 U610 ( .A1(G91), .A2(n643), .ZN(n542) );
  AND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(G299) );
  BUF_X2 U613 ( .A(n546), .Z(n884) );
  NAND2_X1 U614 ( .A1(G102), .A2(n884), .ZN(n549) );
  NAND2_X1 U615 ( .A1(G138), .A2(n547), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT81), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G126), .A2(n879), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n551), .A2(G114), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT80), .B(n552), .ZN(n553) );
  AND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U623 ( .A1(n636), .A2(G64), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT69), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n643), .A2(G90), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT70), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G77), .A2(n639), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n634), .A2(G52), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(G301) );
  INV_X1 U633 ( .A(G301), .ZN(G171) );
  NAND2_X1 U634 ( .A1(G47), .A2(n634), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G60), .A2(n636), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G72), .A2(n639), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G85), .A2(n643), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n570) );
  OR2_X1 U640 ( .A1(n571), .A2(n570), .ZN(G290) );
  INV_X1 U641 ( .A(G57), .ZN(G237) );
  INV_X1 U642 ( .A(G82), .ZN(G220) );
  NAND2_X1 U643 ( .A1(G94), .A2(G452), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U646 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n823) );
  NAND2_X1 U648 ( .A1(n823), .A2(G567), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U650 ( .A1(n636), .A2(G56), .ZN(n575) );
  XNOR2_X1 U651 ( .A(n575), .B(KEYINPUT14), .ZN(n578) );
  NAND2_X1 U652 ( .A1(G43), .A2(n634), .ZN(n576) );
  XNOR2_X1 U653 ( .A(n576), .B(KEYINPUT74), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n643), .A2(G81), .ZN(n579) );
  XNOR2_X1 U656 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U657 ( .A1(G68), .A2(n639), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n967) );
  NAND2_X1 U661 ( .A1(n967), .A2(G860), .ZN(G153) );
  NAND2_X1 U662 ( .A1(G54), .A2(n634), .ZN(n586) );
  NAND2_X1 U663 ( .A1(G66), .A2(n636), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G79), .A2(n639), .ZN(n588) );
  NAND2_X1 U666 ( .A1(G92), .A2(n643), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U669 ( .A(KEYINPUT15), .B(n591), .Z(n968) );
  NOR2_X1 U670 ( .A1(n968), .A2(G868), .ZN(n592) );
  XNOR2_X1 U671 ( .A(n592), .B(KEYINPUT75), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(G284) );
  XOR2_X1 U674 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U675 ( .A(G868), .ZN(n655) );
  NOR2_X1 U676 ( .A1(G286), .A2(n655), .ZN(n596) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U678 ( .A1(n596), .A2(n595), .ZN(G297) );
  INV_X1 U679 ( .A(G860), .ZN(n619) );
  NAND2_X1 U680 ( .A1(n619), .A2(G559), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n597), .A2(n968), .ZN(n598) );
  XNOR2_X1 U682 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U683 ( .A1(n968), .A2(G868), .ZN(n599) );
  NOR2_X1 U684 ( .A1(G559), .A2(n599), .ZN(n601) );
  AND2_X1 U685 ( .A1(n655), .A2(n967), .ZN(n600) );
  NOR2_X1 U686 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n879), .ZN(n602) );
  XNOR2_X1 U688 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n884), .A2(G99), .ZN(n603) );
  NAND2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U691 ( .A1(G135), .A2(n876), .ZN(n606) );
  NAND2_X1 U692 ( .A1(G111), .A2(n878), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n916) );
  XNOR2_X1 U695 ( .A(G2096), .B(n916), .ZN(n610) );
  INV_X1 U696 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U697 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G80), .A2(n639), .ZN(n612) );
  NAND2_X1 U699 ( .A1(G93), .A2(n643), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n634), .A2(G55), .ZN(n613) );
  XNOR2_X1 U702 ( .A(n613), .B(KEYINPUT76), .ZN(n615) );
  NAND2_X1 U703 ( .A1(G67), .A2(n636), .ZN(n614) );
  NAND2_X1 U704 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U705 ( .A1(n617), .A2(n616), .ZN(n654) );
  NAND2_X1 U706 ( .A1(G559), .A2(n968), .ZN(n618) );
  XNOR2_X1 U707 ( .A(n618), .B(n967), .ZN(n652) );
  NAND2_X1 U708 ( .A1(n619), .A2(n652), .ZN(n620) );
  XNOR2_X1 U709 ( .A(n620), .B(KEYINPUT77), .ZN(n621) );
  XOR2_X1 U710 ( .A(n654), .B(n621), .Z(G145) );
  NAND2_X1 U711 ( .A1(G75), .A2(n639), .ZN(n623) );
  NAND2_X1 U712 ( .A1(G88), .A2(n643), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U714 ( .A1(G50), .A2(n634), .ZN(n625) );
  NAND2_X1 U715 ( .A1(G62), .A2(n636), .ZN(n624) );
  NAND2_X1 U716 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U717 ( .A1(n627), .A2(n626), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G87), .A2(n628), .ZN(n630) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U720 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U721 ( .A1(n636), .A2(n631), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(G49), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G48), .A2(n634), .ZN(n635) );
  XNOR2_X1 U725 ( .A(n635), .B(KEYINPUT78), .ZN(n638) );
  NAND2_X1 U726 ( .A1(G61), .A2(n636), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G73), .A2(n639), .ZN(n640) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n643), .A2(G86), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(G305) );
  XNOR2_X1 U733 ( .A(G166), .B(G290), .ZN(n651) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n647) );
  INV_X1 U735 ( .A(G299), .ZN(n977) );
  XNOR2_X1 U736 ( .A(G288), .B(n977), .ZN(n646) );
  XNOR2_X1 U737 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U738 ( .A(n654), .B(n648), .Z(n649) );
  XNOR2_X1 U739 ( .A(n649), .B(G305), .ZN(n650) );
  XNOR2_X1 U740 ( .A(n651), .B(n650), .ZN(n892) );
  XNOR2_X1 U741 ( .A(n652), .B(n892), .ZN(n653) );
  NAND2_X1 U742 ( .A1(n653), .A2(G868), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U751 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n662) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U754 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U755 ( .A1(G96), .A2(n664), .ZN(n828) );
  NAND2_X1 U756 ( .A1(n828), .A2(G2106), .ZN(n668) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n665) );
  NOR2_X1 U758 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U759 ( .A1(G108), .A2(n666), .ZN(n829) );
  NAND2_X1 U760 ( .A1(n829), .A2(G567), .ZN(n667) );
  NAND2_X1 U761 ( .A1(n668), .A2(n667), .ZN(n830) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n669) );
  NOR2_X1 U763 ( .A1(n830), .A2(n669), .ZN(n827) );
  NAND2_X1 U764 ( .A1(n827), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  AND2_X2 U766 ( .A1(G160), .A2(G40), .ZN(n670) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n754) );
  NAND2_X2 U768 ( .A1(n670), .A2(n754), .ZN(n707) );
  XNOR2_X2 U769 ( .A(KEYINPUT93), .B(n707), .ZN(n700) );
  NAND2_X1 U770 ( .A1(n700), .A2(G2072), .ZN(n671) );
  XNOR2_X1 U771 ( .A(KEYINPUT27), .B(n671), .ZN(n676) );
  INV_X1 U772 ( .A(n700), .ZN(n672) );
  NAND2_X1 U773 ( .A1(G1956), .A2(n672), .ZN(n674) );
  XNOR2_X1 U774 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U775 ( .A1(n676), .A2(n675), .ZN(n694) );
  XNOR2_X1 U776 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n677) );
  XNOR2_X1 U777 ( .A(n678), .B(n677), .ZN(n698) );
  NAND2_X1 U778 ( .A1(n700), .A2(G2067), .ZN(n679) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n707), .ZN(n680) );
  XOR2_X1 U780 ( .A(KEYINPUT98), .B(n680), .Z(n681) );
  NAND2_X1 U781 ( .A1(n691), .A2(n968), .ZN(n690) );
  XOR2_X1 U782 ( .A(KEYINPUT96), .B(G1996), .Z(n943) );
  NOR2_X1 U783 ( .A1(n707), .A2(n943), .ZN(n684) );
  XOR2_X1 U784 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n683) );
  XNOR2_X1 U785 ( .A(n684), .B(n683), .ZN(n686) );
  NAND2_X1 U786 ( .A1(n722), .A2(G1341), .ZN(n685) );
  NAND2_X1 U787 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U788 ( .A(KEYINPUT97), .B(n687), .ZN(n688) );
  NAND2_X1 U789 ( .A1(n688), .A2(n967), .ZN(n689) );
  NAND2_X1 U790 ( .A1(n690), .A2(n689), .ZN(n693) );
  OR2_X1 U791 ( .A1(n968), .A2(n691), .ZN(n692) );
  NAND2_X1 U792 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U793 ( .A1(n977), .A2(n694), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U796 ( .A(KEYINPUT29), .B(n699), .Z(n704) );
  INV_X1 U797 ( .A(G1961), .ZN(n971) );
  NAND2_X1 U798 ( .A1(n971), .A2(n722), .ZN(n702) );
  XNOR2_X1 U799 ( .A(KEYINPUT25), .B(G2078), .ZN(n944) );
  NAND2_X1 U800 ( .A1(n700), .A2(n944), .ZN(n701) );
  NAND2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n712), .A2(G171), .ZN(n703) );
  NAND2_X1 U803 ( .A1(n704), .A2(n703), .ZN(n719) );
  INV_X1 U804 ( .A(KEYINPUT92), .ZN(n705) );
  XNOR2_X1 U805 ( .A(n706), .B(n705), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n730), .A2(G8), .ZN(n708) );
  NAND2_X1 U807 ( .A1(G8), .A2(n707), .ZN(n801) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n801), .ZN(n733) );
  NOR2_X1 U809 ( .A1(G171), .A2(n712), .ZN(n713) );
  XNOR2_X1 U810 ( .A(n715), .B(KEYINPUT100), .ZN(n716) );
  INV_X1 U811 ( .A(n716), .ZN(n717) );
  XNOR2_X1 U812 ( .A(n717), .B(KEYINPUT31), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n732) );
  NAND2_X1 U814 ( .A1(G286), .A2(n732), .ZN(n721) );
  XNOR2_X1 U815 ( .A(n721), .B(n720), .ZN(n727) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n801), .ZN(n724) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n722), .ZN(n723) );
  NOR2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U819 ( .A1(G303), .A2(n725), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n728), .A2(G8), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(KEYINPUT32), .ZN(n796) );
  INV_X1 U823 ( .A(n730), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n731), .A2(G8), .ZN(n736) );
  INV_X1 U825 ( .A(n732), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n797) );
  NAND2_X1 U828 ( .A1(G288), .A2(G1976), .ZN(n737) );
  XNOR2_X1 U829 ( .A(n737), .B(KEYINPUT102), .ZN(n976) );
  AND2_X1 U830 ( .A1(n797), .A2(n976), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n796), .A2(n738), .ZN(n742) );
  INV_X1 U832 ( .A(n976), .ZN(n740) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n747) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U835 ( .A1(n747), .A2(n739), .ZN(n975) );
  OR2_X1 U836 ( .A1(n740), .A2(n975), .ZN(n741) );
  AND2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U838 ( .A1(KEYINPUT33), .A2(n746), .ZN(n751) );
  NAND2_X1 U839 ( .A1(KEYINPUT33), .A2(n747), .ZN(n748) );
  NOR2_X1 U840 ( .A1(n801), .A2(n748), .ZN(n749) );
  XNOR2_X1 U841 ( .A(n749), .B(KEYINPUT104), .ZN(n750) );
  XNOR2_X1 U842 ( .A(n753), .B(n752), .ZN(n791) );
  XNOR2_X1 U843 ( .A(G1981), .B(G305), .ZN(n965) );
  XNOR2_X1 U844 ( .A(G1986), .B(G290), .ZN(n974) );
  NAND2_X1 U845 ( .A1(G160), .A2(G40), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n756), .B(KEYINPUT82), .ZN(n816) );
  NAND2_X1 U848 ( .A1(n974), .A2(n816), .ZN(n790) );
  XNOR2_X1 U849 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  NAND2_X1 U850 ( .A1(n879), .A2(G128), .ZN(n757) );
  XNOR2_X1 U851 ( .A(KEYINPUT85), .B(n757), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n878), .A2(G116), .ZN(n758) );
  XOR2_X1 U853 ( .A(KEYINPUT86), .B(n758), .Z(n759) );
  NOR2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U855 ( .A(KEYINPUT35), .B(n761), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n876), .A2(G140), .ZN(n762) );
  XOR2_X1 U857 ( .A(KEYINPUT83), .B(n762), .Z(n764) );
  NAND2_X1 U858 ( .A1(n884), .A2(G104), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U860 ( .A(KEYINPUT84), .B(n765), .ZN(n766) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n766), .ZN(n767) );
  NOR2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U863 ( .A(KEYINPUT36), .B(n769), .ZN(n873) );
  NOR2_X1 U864 ( .A1(n814), .A2(n873), .ZN(n935) );
  NAND2_X1 U865 ( .A1(n935), .A2(n816), .ZN(n812) );
  NAND2_X1 U866 ( .A1(G141), .A2(n876), .ZN(n771) );
  NAND2_X1 U867 ( .A1(G129), .A2(n879), .ZN(n770) );
  NAND2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U869 ( .A1(n884), .A2(G105), .ZN(n772) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n772), .Z(n773) );
  NOR2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n878), .A2(G117), .ZN(n775) );
  NAND2_X1 U873 ( .A1(n776), .A2(n775), .ZN(n869) );
  NAND2_X1 U874 ( .A1(n869), .A2(G1996), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G95), .A2(n884), .ZN(n777) );
  XNOR2_X1 U876 ( .A(n777), .B(KEYINPUT88), .ZN(n784) );
  NAND2_X1 U877 ( .A1(G131), .A2(n876), .ZN(n779) );
  NAND2_X1 U878 ( .A1(G119), .A2(n879), .ZN(n778) );
  NAND2_X1 U879 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U880 ( .A1(G107), .A2(n878), .ZN(n780) );
  XNOR2_X1 U881 ( .A(KEYINPUT87), .B(n780), .ZN(n781) );
  NOR2_X1 U882 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U883 ( .A1(n784), .A2(n783), .ZN(n868) );
  NAND2_X1 U884 ( .A1(n868), .A2(G1991), .ZN(n785) );
  AND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n923) );
  XNOR2_X1 U886 ( .A(KEYINPUT89), .B(n816), .ZN(n787) );
  NOR2_X1 U887 ( .A1(n923), .A2(n787), .ZN(n809) );
  INV_X1 U888 ( .A(n809), .ZN(n788) );
  AND2_X1 U889 ( .A1(n812), .A2(n788), .ZN(n789) );
  NAND2_X1 U890 ( .A1(n790), .A2(n789), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n791), .A2(n514), .ZN(n821) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U893 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  XNOR2_X1 U894 ( .A(KEYINPUT90), .B(n793), .ZN(n794) );
  NOR2_X1 U895 ( .A1(n801), .A2(n794), .ZN(n795) );
  XOR2_X1 U896 ( .A(KEYINPUT91), .B(n795), .Z(n804) );
  NAND2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n800) );
  NOR2_X1 U898 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U899 ( .A1(G8), .A2(n798), .ZN(n799) );
  NAND2_X1 U900 ( .A1(n800), .A2(n799), .ZN(n802) );
  AND2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n819) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n869), .ZN(n913) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n868), .ZN(n917) );
  NOR2_X1 U907 ( .A1(n807), .A2(n917), .ZN(n808) );
  NOR2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U909 ( .A1(n913), .A2(n810), .ZN(n811) );
  XNOR2_X1 U910 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n814), .A2(n873), .ZN(n932) );
  NAND2_X1 U913 ( .A1(n815), .A2(n932), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(n823), .A2(G2106), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U921 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  INV_X1 U930 ( .A(n830), .ZN(G319) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n832) );
  XNOR2_X1 U932 ( .A(G2067), .B(KEYINPUT108), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U934 ( .A(n833), .B(G2678), .Z(n835) );
  XNOR2_X1 U935 ( .A(G2072), .B(G2090), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2100), .Z(n837) );
  XNOR2_X1 U938 ( .A(G2084), .B(G2078), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1986), .B(G1996), .Z(n841) );
  XNOR2_X1 U942 ( .A(G1981), .B(G1966), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U944 ( .A(G1956), .B(G1961), .Z(n843) );
  XNOR2_X1 U945 ( .A(G1976), .B(G1971), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(G2474), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U950 ( .A(G1991), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G124), .A2(n879), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n884), .A2(G100), .ZN(n851) );
  NAND2_X1 U955 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G136), .A2(n876), .ZN(n854) );
  NAND2_X1 U957 ( .A1(G112), .A2(n878), .ZN(n853) );
  NAND2_X1 U958 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U959 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G106), .A2(n884), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G142), .A2(n876), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT45), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G118), .A2(n878), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n879), .A2(G130), .ZN(n862) );
  XOR2_X1 U967 ( .A(KEYINPUT110), .B(n862), .Z(n863) );
  NOR2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U969 ( .A(n865), .B(KEYINPUT46), .Z(n867) );
  XNOR2_X1 U970 ( .A(n916), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(n872) );
  XNOR2_X1 U972 ( .A(G160), .B(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n873), .B(G162), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n890) );
  NAND2_X1 U977 ( .A1(n876), .A2(G139), .ZN(n877) );
  XNOR2_X1 U978 ( .A(KEYINPUT111), .B(n877), .ZN(n888) );
  NAND2_X1 U979 ( .A1(G115), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G127), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n882), .B(KEYINPUT112), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n883), .B(KEYINPUT47), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n884), .A2(G103), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n924) );
  XOR2_X1 U987 ( .A(n924), .B(G164), .Z(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U989 ( .A1(G37), .A2(n891), .ZN(G395) );
  XOR2_X1 U990 ( .A(n892), .B(G286), .Z(n894) );
  XNOR2_X1 U991 ( .A(G171), .B(n968), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(n967), .ZN(n896) );
  NOR2_X1 U994 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2451), .B(G2430), .Z(n898) );
  XNOR2_X1 U996 ( .A(G2438), .B(G2443), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n904) );
  XOR2_X1 U998 ( .A(G2435), .B(G2454), .Z(n900) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U1001 ( .A(G2446), .B(G2427), .Z(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1004 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(n911), .ZN(G401) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n912) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(KEYINPUT113), .B(n914), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n915), .B(KEYINPUT51), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G160), .B(G2084), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n931) );
  XNOR2_X1 U1023 ( .A(G164), .B(G2078), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(G2072), .B(n924), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n925), .B(KEYINPUT114), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(n928), .B(KEYINPUT50), .ZN(n929) );
  XOR2_X1 U1028 ( .A(KEYINPUT115), .B(n929), .Z(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT52), .B(n936), .Z(n937) );
  NOR2_X1 U1033 ( .A1(KEYINPUT55), .A2(n937), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT116), .B(n938), .Z(n939) );
  NAND2_X1 U1035 ( .A1(G29), .A2(n939), .ZN(n1022) );
  XOR2_X1 U1036 ( .A(G34), .B(KEYINPUT121), .Z(n941) );
  XNOR2_X1 U1037 ( .A(G2084), .B(KEYINPUT54), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(n941), .B(n940), .ZN(n961) );
  XOR2_X1 U1039 ( .A(G2090), .B(G35), .Z(n942) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n942), .ZN(n958) );
  XOR2_X1 U1041 ( .A(n943), .B(G32), .Z(n946) );
  XOR2_X1 U1042 ( .A(n944), .B(G27), .Z(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(n947), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(KEYINPUT119), .B(n952), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n953), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(G25), .B(G1991), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n956), .B(KEYINPUT53), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT120), .B(n959), .Z(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT55), .B(n962), .Z(n963) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n963), .ZN(n1018) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XOR2_X1 U1060 ( .A(G1966), .B(G168), .Z(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n966), .Z(n988) );
  XNOR2_X1 U1063 ( .A(n967), .B(G1341), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n968), .B(G1348), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n986) );
  XNOR2_X1 U1066 ( .A(G171), .B(KEYINPUT122), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n984) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1956), .B(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT123), .B(n982), .Z(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n1016) );
  INV_X1 U1079 ( .A(G16), .ZN(n1014) );
  XNOR2_X1 U1080 ( .A(KEYINPUT125), .B(G1966), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(G21), .ZN(n1004) );
  XNOR2_X1 U1082 ( .A(G1961), .B(G5), .ZN(n1002) );
  XOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .Z(n992) );
  XNOR2_X1 U1084 ( .A(G4), .B(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G6), .B(G1981), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G20), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n999), .B(KEYINPUT124), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(KEYINPUT126), .B(n1020), .Z(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

