

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U550 ( .A(n813), .Z(n519) );
  NAND2_X1 U551 ( .A1(G8), .A2(n727), .ZN(n813) );
  XNOR2_X1 U552 ( .A(KEYINPUT98), .B(n531), .ZN(G164) );
  NOR2_X1 U553 ( .A1(n524), .A2(G2104), .ZN(n893) );
  NOR2_X1 U554 ( .A1(n525), .A2(G2105), .ZN(n889) );
  AND2_X2 U555 ( .A1(n696), .A2(n788), .ZN(n728) );
  NAND2_X1 U556 ( .A1(n809), .A2(n989), .ZN(n765) );
  NAND2_X1 U557 ( .A1(n763), .A2(n762), .ZN(n809) );
  XNOR2_X1 U558 ( .A(n698), .B(KEYINPUT30), .ZN(n699) );
  XNOR2_X2 U559 ( .A(n539), .B(KEYINPUT65), .ZN(G160) );
  INV_X1 U560 ( .A(KEYINPUT111), .ZN(n764) );
  XOR2_X1 U561 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  NAND2_X1 U562 ( .A1(n819), .A2(KEYINPUT33), .ZN(n520) );
  INV_X1 U563 ( .A(KEYINPUT27), .ZN(n729) );
  XNOR2_X1 U564 ( .A(n730), .B(n729), .ZN(n731) );
  INV_X1 U565 ( .A(KEYINPUT107), .ZN(n733) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n743) );
  NOR2_X1 U567 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U568 ( .A(n744), .B(n743), .ZN(n748) );
  OR2_X1 U569 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U570 ( .A1(G651), .A2(n638), .ZN(n653) );
  XNOR2_X1 U571 ( .A(n587), .B(n586), .ZN(n906) );
  INV_X1 U572 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G102), .A2(n889), .ZN(n523) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n521), .Z(n890) );
  NAND2_X1 U576 ( .A1(G138), .A2(n890), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n530) );
  INV_X1 U578 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U579 ( .A1(G126), .A2(n893), .ZN(n527) );
  NOR2_X2 U580 ( .A1(n525), .A2(n524), .ZN(n894) );
  NAND2_X1 U581 ( .A1(G114), .A2(n894), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT97), .B(n528), .Z(n529) );
  NOR2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G137), .A2(n890), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G125), .A2(n893), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G113), .A2(n894), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G101), .A2(n889), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n534), .B(KEYINPUT23), .ZN(n535) );
  NOR2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  INV_X1 U593 ( .A(G651), .ZN(n543) );
  NOR2_X1 U594 ( .A1(G543), .A2(n543), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n540), .Z(n661) );
  NAND2_X1 U596 ( .A1(G64), .A2(n661), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G52), .A2(n653), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n551) );
  INV_X1 U599 ( .A(KEYINPUT67), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n543), .A2(n638), .ZN(n544) );
  XNOR2_X2 U601 ( .A(n545), .B(n544), .ZN(n657) );
  NAND2_X1 U602 ( .A1(n657), .A2(G77), .ZN(n548) );
  NOR2_X1 U603 ( .A1(G543), .A2(G651), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT64), .ZN(n654) );
  NAND2_X1 U605 ( .A1(G90), .A2(n654), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U608 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G120), .ZN(G236) );
  INV_X1 U611 ( .A(G69), .ZN(G235) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(G63), .A2(n661), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G51), .A2(n653), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n554), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G89), .A2(n654), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G76), .A2(n657), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U622 ( .A(KEYINPUT5), .B(n558), .ZN(n559) );
  XNOR2_X1 U623 ( .A(KEYINPUT81), .B(n559), .ZN(n560) );
  NOR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(n562), .Z(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U629 ( .A(G223), .B(KEYINPUT73), .ZN(n840) );
  NAND2_X1 U630 ( .A1(n840), .A2(G567), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U632 ( .A1(n661), .A2(G56), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT14), .B(n565), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT12), .B(KEYINPUT75), .Z(n567) );
  NAND2_X1 U635 ( .A1(G81), .A2(n654), .ZN(n566) );
  XNOR2_X1 U636 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(KEYINPUT74), .B(n568), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n657), .A2(G68), .ZN(n569) );
  XNOR2_X1 U639 ( .A(KEYINPUT76), .B(n569), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(n572), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT77), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G43), .A2(n653), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n995) );
  INV_X1 U646 ( .A(G860), .ZN(n626) );
  OR2_X1 U647 ( .A1(n995), .A2(n626), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  INV_X1 U649 ( .A(G868), .ZN(n597) );
  NOR2_X1 U650 ( .A1(G301), .A2(n597), .ZN(n589) );
  XNOR2_X1 U651 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n654), .A2(G92), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G66), .A2(n661), .ZN(n579) );
  NAND2_X1 U654 ( .A1(G54), .A2(n653), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n657), .A2(G79), .ZN(n580) );
  XOR2_X1 U657 ( .A(n580), .B(KEYINPUT78), .Z(n581) );
  NOR2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U660 ( .A(n585), .B(KEYINPUT79), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n906), .A2(G868), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G53), .A2(n653), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G91), .A2(n654), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G78), .A2(n657), .ZN(n592) );
  XNOR2_X1 U667 ( .A(KEYINPUT71), .B(n592), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n661), .A2(G65), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U671 ( .A1(G286), .A2(n597), .ZN(n599) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n626), .A2(G559), .ZN(n600) );
  INV_X1 U675 ( .A(n906), .ZN(n980) );
  NAND2_X1 U676 ( .A1(n600), .A2(n980), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n995), .ZN(n602) );
  XOR2_X1 U679 ( .A(KEYINPUT82), .B(n602), .Z(n605) );
  NOR2_X1 U680 ( .A1(n906), .A2(G559), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G868), .A2(n603), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(KEYINPUT83), .B(n606), .ZN(G282) );
  XOR2_X1 U684 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n608) );
  NAND2_X1 U685 ( .A1(G123), .A2(n893), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n608), .B(n607), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G111), .A2(n894), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G99), .A2(n889), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT85), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G135), .A2(n890), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n933) );
  XNOR2_X1 U694 ( .A(n933), .B(G2096), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT86), .ZN(n618) );
  INV_X1 U696 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G67), .A2(n661), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G55), .A2(n653), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n657), .A2(G80), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G93), .A2(n654), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n674) );
  NAND2_X1 U705 ( .A1(n980), .A2(G559), .ZN(n625) );
  XOR2_X1 U706 ( .A(n995), .B(n625), .Z(n670) );
  NAND2_X1 U707 ( .A1(n626), .A2(n670), .ZN(n627) );
  XOR2_X1 U708 ( .A(n674), .B(n627), .Z(G145) );
  NAND2_X1 U709 ( .A1(n654), .A2(G85), .ZN(n628) );
  XNOR2_X1 U710 ( .A(n628), .B(KEYINPUT66), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G60), .A2(n661), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G47), .A2(n653), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U714 ( .A(KEYINPUT69), .B(n631), .Z(n634) );
  NAND2_X1 U715 ( .A1(G72), .A2(n657), .ZN(n632) );
  XOR2_X1 U716 ( .A(KEYINPUT68), .B(n632), .Z(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(KEYINPUT70), .B(n637), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G87), .A2(n638), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U723 ( .A1(n661), .A2(n641), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G49), .A2(n653), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT87), .B(n642), .Z(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U727 ( .A(KEYINPUT88), .B(n645), .ZN(G288) );
  NAND2_X1 U728 ( .A1(n657), .A2(G75), .ZN(n647) );
  NAND2_X1 U729 ( .A1(G88), .A2(n654), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U731 ( .A(KEYINPUT89), .B(n648), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G62), .A2(n661), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G50), .A2(n653), .ZN(n649) );
  AND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(G303) );
  NAND2_X1 U736 ( .A1(G48), .A2(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G86), .A2(n654), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n657), .A2(G73), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n658), .Z(n659) );
  NOR2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n661), .A2(G61), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(G305) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n664), .B(KEYINPUT90), .ZN(n667) );
  XNOR2_X1 U746 ( .A(G288), .B(G303), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(G299), .ZN(n669) );
  XNOR2_X1 U750 ( .A(G290), .B(n669), .ZN(n909) );
  XNOR2_X1 U751 ( .A(n909), .B(n670), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n671), .B(KEYINPUT91), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n672), .A2(G868), .ZN(n673) );
  XOR2_X1 U754 ( .A(KEYINPUT92), .B(n673), .Z(n676) );
  NOR2_X1 U755 ( .A1(n674), .A2(G868), .ZN(n675) );
  NOR2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U757 ( .A(KEYINPUT93), .B(n677), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U764 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U767 ( .A1(G218), .A2(n683), .ZN(n684) );
  XNOR2_X1 U768 ( .A(KEYINPUT94), .B(n684), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n685), .A2(G96), .ZN(n845) );
  AND2_X1 U770 ( .A1(G2106), .A2(n845), .ZN(n691) );
  NOR2_X1 U771 ( .A1(G235), .A2(G236), .ZN(n686) );
  XNOR2_X1 U772 ( .A(n686), .B(KEYINPUT95), .ZN(n687) );
  NOR2_X1 U773 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G108), .A2(n688), .ZN(n844) );
  NAND2_X1 U775 ( .A1(G567), .A2(n844), .ZN(n689) );
  XOR2_X1 U776 ( .A(KEYINPUT96), .B(n689), .Z(n690) );
  NOR2_X1 U777 ( .A1(n691), .A2(n690), .ZN(G319) );
  INV_X1 U778 ( .A(G319), .ZN(n693) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n843) );
  NAND2_X1 U781 ( .A1(n843), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(G303), .ZN(G166) );
  NOR2_X1 U783 ( .A1(G1976), .A2(G288), .ZN(n694) );
  XNOR2_X1 U784 ( .A(n694), .B(KEYINPUT110), .ZN(n767) );
  NOR2_X1 U785 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U786 ( .A1(n767), .A2(n695), .ZN(n989) );
  NAND2_X1 U787 ( .A1(G160), .A2(G40), .ZN(n787) );
  XNOR2_X1 U788 ( .A(n787), .B(KEYINPUT105), .ZN(n696) );
  NOR2_X1 U789 ( .A1(G1384), .A2(G164), .ZN(n788) );
  INV_X2 U790 ( .A(n728), .ZN(n727) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n813), .ZN(n758) );
  NOR2_X1 U792 ( .A1(G2084), .A2(n727), .ZN(n757) );
  NOR2_X1 U793 ( .A1(n758), .A2(n757), .ZN(n697) );
  NAND2_X1 U794 ( .A1(G8), .A2(n697), .ZN(n698) );
  NOR2_X1 U795 ( .A1(G168), .A2(n699), .ZN(n703) );
  INV_X1 U796 ( .A(G1961), .ZN(n1002) );
  NAND2_X1 U797 ( .A1(n727), .A2(n1002), .ZN(n701) );
  XNOR2_X1 U798 ( .A(G2078), .B(KEYINPUT25), .ZN(n960) );
  NAND2_X1 U799 ( .A1(n728), .A2(n960), .ZN(n700) );
  NAND2_X1 U800 ( .A1(n701), .A2(n700), .ZN(n745) );
  NOR2_X1 U801 ( .A1(G171), .A2(n745), .ZN(n702) );
  XOR2_X1 U802 ( .A(KEYINPUT31), .B(n704), .Z(n755) );
  INV_X1 U803 ( .A(G8), .ZN(n710) );
  NOR2_X1 U804 ( .A1(G2090), .A2(n727), .ZN(n705) );
  XNOR2_X1 U805 ( .A(KEYINPUT109), .B(n705), .ZN(n708) );
  NOR2_X1 U806 ( .A1(G1971), .A2(n519), .ZN(n706) );
  NOR2_X1 U807 ( .A1(G166), .A2(n706), .ZN(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U809 ( .A1(n710), .A2(n709), .ZN(n750) );
  AND2_X1 U810 ( .A1(n755), .A2(n750), .ZN(n749) );
  NAND2_X1 U811 ( .A1(n906), .A2(G1348), .ZN(n711) );
  NAND2_X1 U812 ( .A1(n711), .A2(KEYINPUT26), .ZN(n712) );
  NOR2_X1 U813 ( .A1(G1341), .A2(n712), .ZN(n713) );
  NOR2_X1 U814 ( .A1(n728), .A2(n713), .ZN(n721) );
  NOR2_X1 U815 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n714) );
  NOR2_X1 U816 ( .A1(n995), .A2(n714), .ZN(n719) );
  NAND2_X1 U817 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n716) );
  NAND2_X1 U818 ( .A1(G2067), .A2(n906), .ZN(n715) );
  NAND2_X1 U819 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U820 ( .A1(n717), .A2(n728), .ZN(n718) );
  NAND2_X1 U821 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U822 ( .A1(n721), .A2(n720), .ZN(n726) );
  NAND2_X1 U823 ( .A1(G1348), .A2(n727), .ZN(n723) );
  NAND2_X1 U824 ( .A1(G2067), .A2(n728), .ZN(n722) );
  NAND2_X1 U825 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U826 ( .A1(n906), .A2(n724), .ZN(n725) );
  NOR2_X1 U827 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U828 ( .A1(G1956), .A2(n727), .ZN(n732) );
  NAND2_X1 U829 ( .A1(n728), .A2(G2072), .ZN(n730) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n734) );
  XNOR2_X1 U831 ( .A(n734), .B(n733), .ZN(n739) );
  NOR2_X1 U832 ( .A1(G299), .A2(n739), .ZN(n736) );
  INV_X1 U833 ( .A(KEYINPUT108), .ZN(n735) );
  XNOR2_X1 U834 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U835 ( .A1(n738), .A2(n737), .ZN(n742) );
  NAND2_X1 U836 ( .A1(G299), .A2(n739), .ZN(n740) );
  XNOR2_X1 U837 ( .A(n740), .B(KEYINPUT28), .ZN(n741) );
  NAND2_X1 U838 ( .A1(n742), .A2(n741), .ZN(n744) );
  AND2_X1 U839 ( .A1(n745), .A2(G171), .ZN(n746) );
  XOR2_X1 U840 ( .A(KEYINPUT106), .B(n746), .Z(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n749), .A2(n756), .ZN(n753) );
  INV_X1 U843 ( .A(n750), .ZN(n751) );
  OR2_X1 U844 ( .A1(n751), .A2(G286), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U846 ( .A(n754), .B(KEYINPUT32), .ZN(n763) );
  AND2_X1 U847 ( .A1(n755), .A2(n756), .ZN(n761) );
  AND2_X1 U848 ( .A1(G8), .A2(n757), .ZN(n759) );
  OR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n765), .B(n764), .ZN(n766) );
  NAND2_X1 U851 ( .A1(G288), .A2(G1976), .ZN(n979) );
  NAND2_X1 U852 ( .A1(n766), .A2(n979), .ZN(n806) );
  INV_X1 U853 ( .A(n767), .ZN(n768) );
  NOR2_X1 U854 ( .A1(n519), .A2(n768), .ZN(n769) );
  NAND2_X1 U855 ( .A1(KEYINPUT33), .A2(n769), .ZN(n803) );
  NAND2_X1 U856 ( .A1(G105), .A2(n889), .ZN(n770) );
  XNOR2_X1 U857 ( .A(n770), .B(KEYINPUT38), .ZN(n777) );
  NAND2_X1 U858 ( .A1(G129), .A2(n893), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G141), .A2(n890), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n894), .A2(G117), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT102), .B(n773), .Z(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n885) );
  NAND2_X1 U865 ( .A1(G1996), .A2(n885), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT103), .ZN(n786) );
  INV_X1 U867 ( .A(G1991), .ZN(n961) );
  NAND2_X1 U868 ( .A1(G95), .A2(n889), .ZN(n780) );
  NAND2_X1 U869 ( .A1(G131), .A2(n890), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G119), .A2(n893), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G107), .A2(n894), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n884) );
  NOR2_X1 U875 ( .A1(n961), .A2(n884), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n940) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n835) );
  INV_X1 U878 ( .A(n835), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n940), .A2(n789), .ZN(n828) );
  XOR2_X1 U880 ( .A(KEYINPUT104), .B(n828), .Z(n802) );
  NAND2_X1 U881 ( .A1(n894), .A2(G116), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT101), .B(n790), .Z(n792) );
  NAND2_X1 U883 ( .A1(n893), .A2(G128), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U885 ( .A(KEYINPUT35), .B(n793), .Z(n800) );
  NAND2_X1 U886 ( .A1(n889), .A2(G104), .ZN(n794) );
  XNOR2_X1 U887 ( .A(KEYINPUT99), .B(n794), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n890), .A2(G140), .ZN(n795) );
  XOR2_X1 U889 ( .A(KEYINPUT100), .B(n795), .Z(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT34), .B(n798), .Z(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n801), .ZN(n903) );
  XNOR2_X1 U894 ( .A(KEYINPUT37), .B(G2067), .ZN(n833) );
  NOR2_X1 U895 ( .A1(n903), .A2(n833), .ZN(n942) );
  NAND2_X1 U896 ( .A1(n835), .A2(n942), .ZN(n831) );
  AND2_X1 U897 ( .A1(n802), .A2(n831), .ZN(n817) );
  NAND2_X1 U898 ( .A1(n803), .A2(n817), .ZN(n804) );
  XNOR2_X1 U899 ( .A(G1981), .B(G305), .ZN(n986) );
  OR2_X1 U900 ( .A1(n804), .A2(n986), .ZN(n818) );
  OR2_X1 U901 ( .A1(n519), .A2(n818), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n822) );
  NOR2_X1 U903 ( .A1(G2090), .A2(G303), .ZN(n807) );
  NAND2_X1 U904 ( .A1(G8), .A2(n807), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n810), .A2(n519), .ZN(n815) );
  NOR2_X1 U907 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XOR2_X1 U908 ( .A(n811), .B(KEYINPUT24), .Z(n812) );
  OR2_X1 U909 ( .A1(n519), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n820) );
  INV_X1 U912 ( .A(n818), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n520), .ZN(n821) );
  OR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U915 ( .A(n823), .B(KEYINPUT112), .ZN(n825) );
  XNOR2_X1 U916 ( .A(G290), .B(G1986), .ZN(n992) );
  NAND2_X1 U917 ( .A1(n992), .A2(n835), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n838) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n885), .ZN(n931) );
  AND2_X1 U920 ( .A1(n961), .A2(n884), .ZN(n934) );
  NOR2_X1 U921 ( .A1(G290), .A2(G1986), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n934), .A2(n826), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  NOR2_X1 U924 ( .A1(n931), .A2(n829), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n830), .B(KEYINPUT39), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n903), .A2(n833), .ZN(n943) );
  NAND2_X1 U928 ( .A1(n834), .A2(n943), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U931 ( .A(n839), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U934 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(G188) );
  XOR2_X1 U937 ( .A(G108), .B(KEYINPUT120), .Z(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1976), .B(G1981), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1971), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U954 ( .A(n856), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U957 ( .A(G2474), .B(G1961), .Z(n860) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1956), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n893), .A2(G124), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G112), .A2(n894), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G100), .A2(n889), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n890), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n871) );
  XNOR2_X1 U970 ( .A(G160), .B(KEYINPUT116), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n883) );
  NAND2_X1 U972 ( .A1(G130), .A2(n893), .ZN(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT115), .B(KEYINPUT45), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G106), .A2(n889), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G142), .A2(n890), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n894), .A2(G118), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT114), .B(n876), .Z(n877) );
  NOR2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n881), .B(G162), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n933), .B(n888), .ZN(n901) );
  NAND2_X1 U987 ( .A1(G103), .A2(n889), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G139), .A2(n890), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U990 ( .A1(G127), .A2(n893), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n945) );
  XNOR2_X1 U995 ( .A(G164), .B(n945), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U997 ( .A(n903), .B(n902), .Z(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(n905) );
  XOR2_X1 U999 ( .A(KEYINPUT117), .B(n905), .Z(G395) );
  XNOR2_X1 U1000 ( .A(G171), .B(KEYINPUT118), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n995), .B(n906), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(n909), .B(G286), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n912), .ZN(G397) );
  XOR2_X1 U1006 ( .A(G2454), .B(G2430), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G2451), .B(G2446), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n921) );
  XOR2_X1 U1009 ( .A(G2443), .B(G2427), .Z(n916) );
  XNOR2_X1 U1010 ( .A(G2438), .B(KEYINPUT113), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1012 ( .A(n917), .B(G2435), .Z(n919) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n922) );
  NAND2_X1 U1016 ( .A1(n922), .A2(G14), .ZN(n929) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n929), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n923) );
  XOR2_X1 U1019 ( .A(KEYINPUT49), .B(n923), .Z(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(KEYINPUT119), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n929), .ZN(G401) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n932), .Z(n936) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n938) );
  XOR2_X1 U1031 ( .A(G160), .B(G2084), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n950) );
  XOR2_X1 U1036 ( .A(G2072), .B(n945), .Z(n947) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n948), .Z(n949) );
  NOR2_X1 U1040 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n951), .ZN(n953) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1044 ( .A1(n954), .A2(G29), .ZN(n1033) );
  XNOR2_X1 U1045 ( .A(G2084), .B(G34), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(n955), .B(KEYINPUT54), .ZN(n973) );
  XOR2_X1 U1047 ( .A(G2090), .B(G35), .Z(n956) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(n956), .ZN(n970) );
  XOR2_X1 U1049 ( .A(G1996), .B(G32), .Z(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n965) );
  XOR2_X1 U1054 ( .A(n960), .B(G27), .Z(n963) );
  XOR2_X1 U1055 ( .A(n961), .B(G25), .Z(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(n968), .B(KEYINPUT53), .ZN(n969) );
  NOR2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1061 ( .A(KEYINPUT122), .B(n971), .Z(n972) );
  NOR2_X1 U1062 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1063 ( .A(KEYINPUT55), .B(n974), .Z(n975) );
  NOR2_X1 U1064 ( .A1(G29), .A2(n975), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(KEYINPUT123), .B(n976), .ZN(n977) );
  NAND2_X1 U1066 ( .A1(n977), .A2(G11), .ZN(n1031) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n1001) );
  XOR2_X1 U1068 ( .A(G1956), .B(G299), .Z(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n984) );
  XNOR2_X1 U1070 ( .A(n980), .B(G1348), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n999) );
  XOR2_X1 U1074 ( .A(G168), .B(G1966), .Z(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n988), .ZN(n994) );
  XNOR2_X1 U1078 ( .A(G171), .B(G1961), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n995), .ZN(n996) );
  NOR2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1085 ( .A1(n1001), .A2(n1000), .ZN(n1029) );
  INV_X1 U1086 ( .A(G16), .ZN(n1027) );
  XNOR2_X1 U1087 ( .A(n1002), .B(G5), .ZN(n1023) );
  XOR2_X1 U1088 ( .A(G1966), .B(G21), .Z(n1014) );
  XNOR2_X1 U1089 ( .A(KEYINPUT59), .B(G4), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(KEYINPUT125), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1348), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1011), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(n1012), .B(KEYINPUT126), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT61), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1114 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

