//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n227), .B(new_n231), .ZN(G358));
  INV_X1    g0032(.A(G50), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(G68), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  XNOR2_X1  g0043(.A(KEYINPUT3), .B(G33), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT67), .B(G1698), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n244), .A2(new_n245), .A3(G222), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(new_n214), .B2(new_n244), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n244), .A2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n247), .B1(new_n250), .B2(G223), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(new_n253), .A3(G274), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  INV_X1    g0061(.A(new_n209), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n252), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT66), .A3(new_n257), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G226), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n253), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n254), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G190), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n265), .B1(new_n266), .B2(new_n269), .C1(new_n251), .C2(new_n253), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G200), .ZN(new_n274));
  INV_X1    g0074(.A(G13), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G1), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n203), .B2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n277), .A2(new_n209), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n267), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G50), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n280), .A2(new_n209), .A3(new_n281), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n210), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G58), .A2(G68), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n210), .B1(new_n293), .B2(new_n233), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n285), .B(new_n295), .C1(G50), .C2(new_n277), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT9), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n272), .A2(new_n274), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n271), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n273), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n305), .A3(new_n296), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT72), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n245), .A2(G226), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G232), .A2(G1698), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n244), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT70), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n253), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n258), .A2(new_n259), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT66), .B1(new_n263), .B2(new_n257), .ZN(new_n318));
  OAI21_X1  g0118(.A(G238), .B1(new_n269), .B2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n253), .B2(new_n268), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT13), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(new_n321), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(new_n260), .B2(new_n264), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n309), .B2(new_n310), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n328), .B1(new_n333), .B2(new_n314), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n326), .A2(new_n327), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n323), .A2(G190), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n283), .A2(G68), .A3(new_n284), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n291), .A2(new_n233), .B1(new_n210), .B2(G68), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n288), .A2(new_n214), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n286), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n277), .A2(G68), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G200), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n323), .B2(new_n335), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n308), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n349), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n346), .A4(new_n336), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n307), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n287), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n284), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n282), .B1(new_n277), .B2(new_n354), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G58), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n235), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n293), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n290), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n368), .A3(G33), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n329), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n329), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(KEYINPUT75), .A3(new_n329), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n365), .B1(new_n379), .B2(G68), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n244), .B2(G20), .ZN(new_n382));
  INV_X1    g0182(.A(new_n331), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n366), .A2(new_n368), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n279), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n382), .B1(new_n385), .B2(new_n371), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n362), .B1(new_n386), .B2(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n286), .B1(new_n387), .B2(KEYINPUT16), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n357), .B1(new_n380), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n245), .A2(G223), .ZN(new_n390));
  INV_X1    g0190(.A(G87), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n374), .A2(new_n390), .B1(new_n279), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G1698), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n266), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n369), .A2(new_n329), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n369), .A2(new_n398), .A3(new_n329), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n253), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n269), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n260), .A2(new_n264), .B1(G232), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G169), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n392), .B1(new_n399), .B2(new_n397), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n403), .B(G179), .C1(new_n406), .C2(new_n253), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n389), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT18), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n389), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  OAI21_X1  g0213(.A(G200), .B1(new_n401), .B2(new_n404), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n403), .B(G190), .C1(new_n406), .C2(new_n253), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n389), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n369), .A2(KEYINPUT75), .A3(new_n329), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT75), .B1(new_n369), .B2(new_n329), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n210), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n372), .B1(new_n421), .B2(new_n381), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n364), .B1(new_n422), .B2(new_n235), .ZN(new_n423));
  INV_X1    g0223(.A(new_n286), .ZN(new_n424));
  INV_X1    g0224(.A(new_n362), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT7), .B1(new_n332), .B2(new_n210), .ZN(new_n426));
  INV_X1    g0226(.A(new_n371), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n331), .B1(new_n428), .B2(G33), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n425), .B1(new_n430), .B2(new_n235), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n431), .B2(new_n363), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n356), .B1(new_n423), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n418), .A2(new_n433), .A3(KEYINPUT17), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n410), .A2(new_n412), .A3(new_n417), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT73), .A2(G169), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n316), .A2(new_n322), .A3(KEYINPUT13), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n327), .B1(new_n326), .B2(new_n334), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n323), .A2(new_n335), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(new_n438), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n323), .A2(G179), .A3(new_n335), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n346), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n244), .A2(new_n245), .A3(G232), .ZN(new_n450));
  INV_X1    g0250(.A(G107), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n244), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n250), .B2(G238), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n253), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n265), .B1(new_n213), .B2(new_n269), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n283), .A2(G77), .A3(new_n284), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n354), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT15), .B(G87), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n288), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n275), .A2(new_n210), .A3(G1), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n461), .A2(new_n286), .B1(new_n214), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n457), .A2(new_n304), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n456), .A2(new_n302), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n458), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n456), .B2(G190), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n348), .B2(new_n456), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n353), .A2(new_n436), .A3(new_n449), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n245), .A2(G244), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n374), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n394), .A2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G244), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(KEYINPUT78), .A3(new_n329), .A4(new_n369), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n474), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT79), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n474), .A2(new_n481), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  INV_X1    g0286(.A(G283), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n279), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G250), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n473), .A2(new_n482), .B1(new_n489), .B2(new_n394), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(new_n244), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n328), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n256), .A2(G1), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n263), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n328), .B1(new_n495), .B2(new_n494), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G257), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n493), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n304), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n282), .B1(new_n267), .B2(G33), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n462), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n451), .A3(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(KEYINPUT6), .B2(new_n508), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT77), .B(G107), .Z(new_n513));
  XNOR2_X1  g0313(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n386), .A2(G107), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(new_n286), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n502), .B1(new_n492), .B2(new_n328), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n302), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n505), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n493), .A2(G190), .A3(new_n503), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n522), .B(new_n518), .C1(new_n348), .C2(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n283), .B1(G1), .B2(new_n279), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n526), .A2(new_n527), .B1(new_n277), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n530), .A3(G20), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n286), .A2(KEYINPUT83), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT83), .B1(new_n286), .B2(new_n534), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n210), .B1(new_n508), .B2(G33), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n488), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n286), .A2(new_n534), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n540), .B1(new_n544), .B2(new_n535), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n532), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n499), .A2(G270), .B1(new_n497), .B2(new_n263), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G264), .A2(G1698), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n478), .B2(new_n501), .ZN(new_n550));
  XOR2_X1   g0350(.A(KEYINPUT82), .B(G303), .Z(new_n551));
  AOI22_X1  g0351(.A1(new_n370), .A2(new_n550), .B1(new_n332), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n548), .B1(new_n552), .B2(new_n253), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G169), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n525), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT81), .B(G116), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n506), .A2(G116), .B1(new_n462), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n533), .B(new_n540), .C1(new_n544), .C2(new_n535), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT21), .A3(G169), .A4(new_n553), .ZN(new_n561));
  INV_X1    g0361(.A(new_n553), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(G179), .A3(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n555), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n553), .A2(G200), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n548), .B(G190), .C1(new_n552), .C2(new_n253), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT84), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n547), .A2(new_n569), .A3(new_n566), .A4(new_n565), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n495), .A2(KEYINPUT80), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT80), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n256), .B2(G1), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n572), .A2(new_n574), .A3(G250), .A4(new_n253), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n263), .A2(new_n495), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n556), .A2(new_n279), .ZN(new_n579));
  INV_X1    g0379(.A(G238), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n478), .A2(new_n580), .B1(new_n479), .B2(new_n394), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n579), .B1(new_n370), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n578), .B1(new_n582), .B2(new_n253), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n369), .A2(new_n210), .A3(G68), .A4(new_n329), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n288), .B2(new_n508), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(new_n314), .B2(KEYINPUT19), .ZN(new_n588));
  NOR3_X1   g0388(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n585), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n286), .B1(new_n462), .B2(new_n460), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n245), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n592), .A2(new_n374), .B1(new_n279), .B2(new_n556), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n577), .B1(new_n593), .B2(new_n328), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n506), .A2(G87), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n584), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n210), .A2(G87), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n332), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n451), .A2(G20), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n531), .A2(new_n210), .A3(G33), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n598), .A2(new_n391), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n370), .A2(new_n210), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n210), .A2(new_n369), .A3(new_n329), .A4(new_n607), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT24), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n286), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n478), .A2(new_n489), .B1(new_n501), .B2(new_n394), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n370), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G294), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n279), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n328), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n499), .A2(G264), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(G190), .A3(new_n498), .A4(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n370), .A2(new_n615), .B1(G33), .B2(G294), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n498), .B(new_n620), .C1(new_n622), .C2(new_n253), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n506), .A2(G107), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n277), .A2(G107), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT25), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n614), .A2(new_n621), .A3(new_n624), .A4(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n619), .A2(new_n302), .A3(new_n498), .A4(new_n620), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n304), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n424), .B1(new_n609), .B2(new_n612), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n628), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n590), .A2(new_n286), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n460), .A2(new_n462), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n636), .C1(new_n460), .C2(new_n526), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n583), .A2(new_n304), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n594), .A2(new_n302), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n597), .A2(new_n630), .A3(new_n634), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n564), .A2(new_n571), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n471), .A2(new_n524), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n306), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n410), .A2(new_n412), .ZN(new_n645));
  INV_X1    g0445(.A(new_n466), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n351), .A2(new_n346), .A3(new_n336), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n646), .A2(new_n647), .B1(new_n448), .B2(new_n447), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n417), .A2(new_n434), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n644), .B1(new_n650), .B2(new_n301), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n584), .A2(new_n595), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT85), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n591), .A2(new_n654), .A3(new_n596), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n591), .B2(new_n596), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n657), .A2(new_n640), .A3(new_n630), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n555), .A2(new_n561), .A3(new_n563), .A4(new_n634), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n521), .A3(new_n659), .A4(new_n523), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT86), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n518), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n504), .B2(G200), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n664), .A2(new_n522), .B1(new_n505), .B2(new_n520), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(KEYINPUT86), .A3(new_n659), .A4(new_n658), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n657), .A2(new_n640), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n505), .A4(new_n520), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n640), .A2(new_n597), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n521), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n671), .A2(new_n673), .A3(new_n640), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n651), .B1(new_n471), .B2(new_n675), .ZN(G369));
  AND2_X1   g0476(.A1(new_n568), .A2(new_n570), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n555), .A2(new_n561), .A3(new_n563), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n276), .A2(new_n210), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(G213), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n547), .A2(new_n686), .ZN(new_n687));
  MUX2_X1   g0487(.A(new_n679), .B(new_n678), .S(new_n687), .Z(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT87), .Z(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n630), .A2(new_n634), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n685), .B1(new_n633), .B2(new_n628), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n634), .B2(new_n686), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n564), .A2(new_n685), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(new_n692), .ZN(new_n698));
  INV_X1    g0498(.A(new_n634), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n686), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT88), .Z(G399));
  INV_X1    g0502(.A(new_n204), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n589), .A2(new_n527), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n704), .A2(new_n267), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n208), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  NOR3_X1   g0508(.A1(new_n675), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n521), .A2(KEYINPUT26), .A3(new_n672), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT26), .B1(new_n521), .B2(new_n668), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n640), .A4(new_n660), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(new_n713), .B2(new_n686), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n548), .B(G179), .C1(new_n552), .C2(new_n253), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n620), .B1(new_n622), .B2(new_n253), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n716), .A2(new_n717), .A3(new_n583), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT90), .B(KEYINPUT30), .C1(new_n519), .C2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT90), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n493), .A2(new_n503), .A3(new_n718), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n493), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n503), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n553), .A2(new_n583), .A3(new_n302), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT89), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT89), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n553), .A2(new_n583), .A3(new_n728), .A4(new_n302), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n623), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n725), .B1(new_n730), .B2(new_n519), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n685), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n730), .A2(new_n519), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n721), .A2(new_n722), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n725), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n686), .A2(new_n733), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n732), .A2(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n679), .A2(new_n665), .A3(new_n641), .A4(new_n686), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n715), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n708), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n275), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n267), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n704), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n209), .B1(G20), .B2(new_n304), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n210), .A2(new_n302), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G190), .A3(new_n348), .ZN(new_n753));
  INV_X1    g0553(.A(G322), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n332), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n210), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n756), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n755), .B(new_n760), .C1(G329), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n752), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(G317), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT33), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n767), .A2(KEYINPUT33), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n210), .A2(new_n348), .A3(G179), .A4(G190), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n772), .A2(G303), .B1(new_n773), .B2(G283), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n302), .A2(new_n348), .A3(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(G326), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n777), .A2(new_n617), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n764), .A2(new_n770), .A3(new_n774), .A4(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n766), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n783), .A2(new_n235), .B1(new_n771), .B2(new_n391), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n763), .A2(G159), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n785), .A2(KEYINPUT32), .B1(new_n233), .B2(new_n778), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT91), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n753), .B(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G58), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n244), .B1(new_n758), .B2(new_n214), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(KEYINPUT32), .B2(new_n785), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n777), .A2(new_n508), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G107), .B2(new_n773), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n787), .A2(new_n791), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n751), .B1(new_n782), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n750), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n703), .A2(new_n332), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G355), .B1(new_n527), .B2(new_n703), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n376), .A2(new_n377), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n703), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n208), .A2(new_n256), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n239), .B2(new_n256), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n803), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n749), .B(new_n797), .C1(new_n801), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n800), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n688), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n690), .A2(new_n749), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n689), .A2(G330), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(G396));
  NOR2_X1   g0617(.A1(new_n675), .A2(new_n685), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n467), .A2(new_n685), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n469), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n466), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n466), .B2(new_n685), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT96), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n470), .A2(new_n686), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n667), .B2(new_n674), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n748), .B1(new_n829), .B2(new_n741), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n742), .A3(new_n828), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n822), .A2(new_n798), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n750), .A2(G77), .A3(new_n798), .ZN(new_n834));
  INV_X1    g0634(.A(new_n773), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n391), .B1(new_n762), .B2(new_n759), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT94), .Z(new_n837));
  OAI21_X1  g0637(.A(new_n332), .B1(new_n758), .B2(new_n556), .ZN(new_n838));
  INV_X1    g0638(.A(new_n753), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(G294), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n794), .B1(G107), .B2(new_n772), .ZN(new_n841));
  INV_X1    g0641(.A(new_n778), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n766), .A2(G283), .B1(new_n842), .B2(G303), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n837), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n835), .A2(new_n235), .B1(new_n777), .B2(new_n358), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n771), .A2(new_n233), .B1(new_n762), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n804), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n842), .A2(G137), .B1(new_n757), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G143), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n289), .B2(new_n783), .C1(new_n789), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n853), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n749), .B(new_n834), .C1(new_n857), .C2(new_n750), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n833), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n832), .A2(new_n859), .ZN(G384));
  OR2_X1    g0660(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n861), .A2(G116), .A3(new_n211), .A4(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT36), .Z(new_n864));
  OAI211_X1 g0664(.A(new_n208), .B(G77), .C1(new_n358), .C2(new_n235), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n267), .B(G13), .C1(new_n865), .C2(new_n234), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n447), .A2(new_n448), .A3(new_n686), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n418), .A2(new_n433), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n379), .A2(G68), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n424), .B1(new_n870), .B2(new_n364), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n421), .A2(new_n381), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n235), .B1(new_n872), .B2(new_n373), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n363), .B1(new_n873), .B2(new_n362), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n356), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n408), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n683), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n389), .A2(new_n416), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n423), .A2(new_n432), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n881), .A2(new_n357), .B1(new_n405), .B2(new_n407), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT99), .B1(new_n433), .B2(new_n683), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT99), .ZN(new_n885));
  INV_X1    g0685(.A(new_n683), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n388), .B1(new_n870), .B2(new_n364), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n356), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n879), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n435), .A2(new_n878), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n892), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n884), .A2(new_n888), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n869), .A2(new_n409), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n901), .A2(new_n891), .B1(new_n435), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n902), .B2(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n435), .A2(new_n899), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n890), .B1(new_n883), .B2(new_n889), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(KEYINPUT100), .A3(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n879), .A2(new_n891), .B1(new_n435), .B2(new_n878), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n910), .A2(KEYINPUT101), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT101), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n903), .B(new_n909), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n868), .B(new_n897), .C1(new_n913), .C2(new_n896), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n448), .A2(new_n685), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n449), .A2(new_n647), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT98), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n350), .A2(new_n352), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n915), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g0722(.A(KEYINPUT98), .B(new_n915), .C1(new_n918), .C2(new_n919), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n466), .A2(new_n685), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT97), .Z(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n827), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n894), .A2(new_n895), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n927), .A2(new_n928), .B1(new_n645), .B2(new_n886), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT102), .B1(new_n914), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n897), .B1(new_n913), .B2(new_n896), .ZN(new_n931));
  INV_X1    g0731(.A(new_n868), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT102), .ZN(new_n934));
  INV_X1    g0734(.A(new_n929), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n651), .ZN(new_n938));
  INV_X1    g0738(.A(new_n471), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n715), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n937), .B(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n725), .B(new_n734), .C1(new_n719), .C2(new_n723), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n737), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n739), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT31), .B1(new_n732), .B2(KEYINPUT103), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT103), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n946), .A3(new_n685), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n924), .A2(new_n823), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  INV_X1    g0751(.A(new_n928), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n735), .A2(KEYINPUT90), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n721), .A2(new_n720), .A3(new_n722), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n731), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT103), .B1(new_n956), .B2(new_n686), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(new_n733), .A3(new_n947), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n642), .A2(new_n524), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n959), .A2(new_n686), .B1(new_n737), .B2(new_n942), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n447), .B1(new_n350), .B2(new_n352), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT98), .B1(new_n962), .B2(new_n915), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n920), .A2(new_n917), .A3(new_n921), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n822), .B1(new_n965), .B2(new_n916), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n907), .A2(KEYINPUT100), .A3(new_n908), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT100), .B1(new_n907), .B2(new_n908), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n910), .A2(KEYINPUT38), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT101), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n910), .A2(KEYINPUT101), .A3(KEYINPUT38), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n967), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n953), .B1(new_n976), .B2(new_n951), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n939), .A3(new_n961), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n951), .B1(new_n894), .B2(new_n895), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n913), .A2(new_n950), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(KEYINPUT40), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n471), .B2(new_n948), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(new_n983), .A3(G330), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n941), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n267), .B2(new_n745), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n941), .A2(new_n984), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n867), .B1(new_n986), .B2(new_n987), .ZN(G367));
  OAI221_X1 g0788(.A(new_n801), .B1(new_n204), .B2(new_n460), .C1(new_n807), .C2(new_n231), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(new_n748), .ZN(new_n990));
  INV_X1    g0790(.A(G159), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n783), .A2(new_n991), .B1(new_n850), .B2(new_n778), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n835), .A2(new_n214), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n332), .B1(new_n839), .B2(G150), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G50), .A2(new_n757), .B1(new_n763), .B2(G137), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n772), .A2(G58), .B1(new_n776), .B2(G68), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n771), .B2(new_n556), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n771), .B2(new_n1001), .C1(new_n783), .C2(new_n617), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n758), .A2(new_n487), .B1(new_n762), .B2(new_n767), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G107), .B2(new_n776), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n790), .A2(new_n551), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n835), .A2(new_n508), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G311), .B2(new_n842), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n804), .A4(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n998), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  OR3_X1    g0811(.A1(new_n655), .A2(new_n656), .A3(new_n686), .ZN(new_n1012));
  MUX2_X1   g0812(.A(new_n640), .B(new_n668), .S(new_n1012), .Z(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT104), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n990), .B1(new_n751), .B2(new_n1011), .C1(new_n1015), .C2(new_n812), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n696), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n521), .B(new_n523), .C1(new_n518), .C2(new_n686), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT105), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n521), .B2(new_n686), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT107), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1019), .A2(new_n634), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n521), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n1025), .A2(KEYINPUT106), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT106), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1027), .A2(new_n686), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1020), .A2(new_n698), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT42), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1024), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1023), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1020), .A2(new_n700), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT44), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n1020), .A2(new_n700), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n696), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n698), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n695), .B2(new_n697), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n690), .B(new_n1046), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1017), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n743), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n743), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n704), .B(KEYINPUT41), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n747), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1016), .B1(new_n1037), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT110), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n1016), .C1(new_n1037), .C2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(G387));
  AOI22_X1  g0858(.A1(new_n802), .A2(new_n705), .B1(new_n451), .B2(new_n703), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n227), .A2(new_n256), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT50), .B1(new_n354), .B2(new_n233), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n354), .A2(KEYINPUT50), .A3(new_n233), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n806), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1059), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n749), .B1(new_n1066), .B2(new_n801), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G68), .A2(new_n757), .B1(new_n763), .B2(G150), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n233), .B2(new_n753), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1007), .B(new_n1069), .C1(new_n354), .C2(new_n766), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n771), .A2(new_n214), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n777), .A2(new_n460), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G159), .C2(new_n842), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n805), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n766), .A2(G311), .B1(new_n551), .B2(new_n757), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n754), .B2(new_n778), .C1(new_n789), .C2(new_n767), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n772), .A2(G294), .B1(new_n776), .B2(G283), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT111), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n835), .A2(new_n556), .B1(new_n762), .B2(new_n779), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n804), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1074), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT112), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1067), .B1(new_n695), .B2(new_n812), .C1(new_n1090), .C2(new_n751), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT113), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n747), .B2(new_n1047), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1047), .A2(new_n743), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1047), .A2(new_n743), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n704), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(G393));
  NAND2_X1  g0897(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1095), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n704), .A3(new_n1049), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1044), .A2(new_n747), .A3(new_n1048), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n777), .A2(new_n556), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n332), .B1(new_n835), .B2(new_n451), .C1(new_n758), .C2(new_n617), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n551), .C2(new_n766), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n759), .A2(new_n753), .B1(new_n778), .B2(new_n767), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT52), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n771), .A2(new_n487), .B1(new_n762), .B2(new_n754), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT115), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1104), .A2(new_n1106), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n783), .A2(new_n233), .B1(new_n771), .B2(new_n235), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n777), .A2(new_n214), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n289), .A2(new_n778), .B1(new_n753), .B2(new_n991), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n758), .A2(new_n287), .B1(new_n762), .B2(new_n850), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G87), .B2(new_n773), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .A4(new_n805), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n751), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n801), .B1(new_n508), .B2(new_n204), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n806), .B2(new_n242), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT114), .Z(new_n1123));
  NOR3_X1   g0923(.A1(new_n1120), .A2(new_n1123), .A3(new_n749), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1020), .B2(new_n812), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1101), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1100), .A2(new_n1126), .ZN(G390));
  NAND2_X1  g0927(.A1(new_n961), .A2(G330), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1128), .A2(new_n471), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n714), .B1(new_n818), .B2(new_n710), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n651), .C1(new_n1130), .C2(new_n471), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n924), .B1(new_n742), .B2(new_n823), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n961), .A2(G330), .A3(new_n966), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1132), .A2(new_n1134), .B1(new_n827), .B2(new_n926), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n742), .A2(new_n823), .A3(new_n924), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n924), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1128), .B2(new_n822), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n926), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n823), .A2(new_n713), .A3(new_n686), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1131), .B1(new_n1135), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n913), .B(new_n868), .C1(new_n1141), .C2(new_n1137), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n927), .A2(new_n868), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n931), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1134), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1145), .B(new_n1136), .C1(new_n931), .C2(new_n1146), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1143), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n704), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1148), .A2(new_n747), .A3(new_n1149), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n750), .A2(new_n798), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n749), .B1(new_n287), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n758), .A2(new_n1157), .B1(new_n846), .B2(new_n753), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n332), .B(new_n1158), .C1(G125), .C2(new_n763), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n771), .A2(KEYINPUT53), .A3(new_n289), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT53), .B1(new_n771), .B2(new_n289), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G137), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n783), .A2(new_n1163), .B1(new_n1164), .B2(new_n778), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n835), .A2(new_n233), .B1(new_n777), .B2(new_n991), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n842), .A2(G283), .B1(new_n757), .B2(G97), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n451), .B2(new_n783), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT116), .Z(new_n1170));
  OAI221_X1 g0970(.A(new_n332), .B1(new_n762), .B2(new_n617), .C1(new_n753), .C2(new_n527), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n835), .A2(new_n235), .B1(new_n391), .B2(new_n771), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n1113), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1162), .A2(new_n1167), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1156), .B1(new_n751), .B2(new_n1174), .C1(new_n931), .C2(new_n799), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1154), .A2(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT117), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(KEYINPUT117), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1153), .B1(new_n1177), .B2(new_n1178), .ZN(G378));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n930), .A2(new_n936), .A3(KEYINPUT121), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n296), .A2(new_n886), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n307), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT120), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n301), .A2(new_n306), .A3(new_n1182), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1182), .B1(new_n301), .B2(new_n306), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n644), .B(new_n1183), .C1(new_n299), .C2(new_n300), .ZN(new_n1189));
  OAI21_X1  g0989(.A(KEYINPUT120), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  AND3_X1   g0991(.A1(new_n1187), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(G330), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n982), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n951), .B1(new_n913), .B2(new_n950), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G330), .B(new_n1194), .C1(new_n1198), .C2(new_n980), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1181), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1131), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1152), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1180), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1194), .B1(new_n977), .B2(G330), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1199), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT122), .B1(new_n1207), .B2(new_n937), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n930), .A2(new_n936), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT122), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1200), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n937), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1180), .B1(new_n1152), .B2(new_n1202), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1204), .A2(new_n1215), .A3(new_n704), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1195), .A2(new_n798), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n766), .A2(G97), .B1(new_n842), .B2(G116), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1071), .B1(G68), .B2(new_n776), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G41), .B1(new_n839), .B2(G107), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n460), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1221), .A2(new_n757), .B1(new_n763), .B2(G283), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n773), .A2(G58), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT118), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n805), .A3(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT58), .Z(new_n1227));
  AOI21_X1  g1027(.A(G41), .B1(new_n805), .B2(G33), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n758), .A2(new_n1163), .B1(new_n1164), .B2(new_n753), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n842), .A2(G125), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n771), .B2(new_n1157), .C1(new_n783), .C2(new_n846), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(G150), .C2(new_n776), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n773), .A2(G159), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1227), .B1(G50), .B2(new_n1228), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT119), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n751), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1240), .B2(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n749), .B1(new_n233), .B2(new_n1155), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1217), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1201), .B2(new_n746), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1216), .A2(new_n1246), .ZN(G375));
  AOI21_X1  g1047(.A(new_n749), .B1(new_n235), .B2(new_n1155), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n839), .A2(G283), .B1(new_n763), .B2(G303), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n332), .C1(new_n451), .C2(new_n758), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G294), .A2(new_n842), .B1(new_n772), .B2(G97), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n556), .B2(new_n783), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1250), .A2(new_n1252), .A3(new_n993), .A4(new_n1072), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n783), .A2(new_n1157), .B1(new_n771), .B2(new_n991), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G150), .A2(new_n757), .B1(new_n763), .B2(G128), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n233), .B2(new_n777), .C1(new_n789), .C2(new_n1163), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G132), .C2(new_n842), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1225), .A2(new_n804), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1248), .B1(new_n1259), .B2(new_n751), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1137), .B2(new_n798), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1135), .A2(new_n1142), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n747), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1144), .A2(new_n1051), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1262), .A2(new_n1202), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(G381));
  OR2_X1    g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1267), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1057), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n704), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1245), .B1(new_n1273), .B2(new_n1204), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1153), .A2(new_n1176), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1271), .A2(new_n1276), .ZN(G407));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n684), .A3(new_n1275), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G213), .B(new_n1278), .C1(new_n1271), .C2(new_n1276), .ZN(G409));
  OAI211_X1 g1079(.A(new_n1016), .B(G390), .C1(new_n1037), .C2(new_n1052), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G393), .B(G396), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1057), .B2(G390), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1281), .B(KEYINPUT125), .ZN(new_n1284));
  INV_X1    g1084(.A(G390), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1053), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1280), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1265), .B1(KEYINPUT60), .B2(new_n1144), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1135), .A2(new_n1131), .A3(new_n1142), .A4(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n704), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1263), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n832), .A3(new_n859), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1263), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1295));
  INV_X1    g1095(.A(G213), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(G343), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G2897), .ZN(new_n1298));
  XOR2_X1   g1098(.A(new_n1298), .B(KEYINPUT124), .Z(new_n1299));
  AND3_X1   g1099(.A1(new_n1294), .A2(new_n1295), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1213), .A2(new_n747), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1152), .A2(new_n1202), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1200), .B1(new_n1209), .B2(KEYINPUT121), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1207), .A2(new_n1181), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1051), .B(new_n1304), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1244), .A3(new_n1307), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1274), .A2(G378), .B1(new_n1275), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1302), .B1(new_n1309), .B2(new_n1297), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1216), .A2(G378), .A3(new_n1246), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1275), .ZN(new_n1314));
  AOI211_X1 g1114(.A(new_n1312), .B(new_n1297), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1310), .B(new_n1311), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1312), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1297), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1289), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1302), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1315), .A2(KEYINPUT63), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1321), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1323), .A2(new_n1330), .ZN(G405));
  AND2_X1   g1131(.A1(G375), .A2(new_n1275), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1313), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT126), .ZN(new_n1335));
  OAI21_X1  g1135(.A(KEYINPUT127), .B1(new_n1312), .B2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(KEYINPUT127), .B2(new_n1312), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1334), .A2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1336), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1289), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1324), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(G402));
endmodule


