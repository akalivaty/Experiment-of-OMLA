//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n463), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n468), .A2(new_n476), .A3(new_n479), .A4(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n475), .B1(new_n482), .B2(new_n486), .ZN(G160));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n485), .C2(G112), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n486), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT69), .B1(new_n489), .B2(new_n471), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n469), .A2(new_n494), .A3(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n497), .B2(G136), .ZN(G162));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n472), .A2(G138), .A3(new_n473), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n468), .A2(new_n476), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT4), .A2(G138), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n485), .A2(new_n508), .B1(G126), .B2(G2105), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n502), .B(new_n506), .C1(new_n509), .C2(new_n469), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(G50), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n519), .B1(new_n524), .B2(G651), .ZN(new_n525));
  AOI211_X1 g100(.A(KEYINPUT71), .B(new_n514), .C1(new_n521), .C2(new_n523), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n516), .B(new_n518), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n512), .A2(new_n516), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(G88), .B(new_n529), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n527), .A2(new_n530), .A3(KEYINPUT72), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT72), .B1(new_n527), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n515), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n536), .B(new_n515), .C1(new_n531), .C2(new_n532), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  XNOR2_X1  g115(.A(KEYINPUT70), .B(KEYINPUT6), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT71), .B1(new_n541), .B2(new_n514), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n524), .A2(new_n519), .A3(G651), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n528), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT74), .B(G89), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n512), .ZN(new_n548));
  INV_X1    g123(.A(G63), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT7), .ZN(new_n551));
  NAND3_X1  g126(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n550), .A2(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n542), .A2(new_n543), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n555), .A2(G543), .A3(new_n516), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G51), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G286));
  INV_X1    g133(.A(G286), .ZN(G168));
  NAND2_X1  g134(.A1(new_n556), .A2(G52), .ZN(new_n560));
  NAND2_X1  g135(.A1(G77), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G64), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n548), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n544), .A2(G90), .B1(G651), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G301));
  INV_X1    g140(.A(G301), .ZN(G171));
  XOR2_X1   g141(.A(KEYINPUT75), .B(G81), .Z(new_n567));
  NAND2_X1  g142(.A1(new_n544), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n514), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n555), .A2(G543), .A3(new_n516), .ZN(new_n571));
  INV_X1    g146(.A(G43), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n568), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  NAND4_X1  g150(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  NAND4_X1  g155(.A1(new_n555), .A2(G53), .A3(G543), .A4(new_n516), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT9), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(KEYINPUT77), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n514), .B1(new_n583), .B2(KEYINPUT77), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(new_n585), .B1(new_n544), .B2(G91), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G299));
  OAI21_X1  g162(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n544), .B2(G87), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n555), .A2(G49), .A3(G543), .A4(new_n516), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  OAI211_X1 g167(.A(G86), .B(new_n529), .C1(new_n525), .C2(new_n526), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT78), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n544), .A2(new_n595), .A3(G86), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n514), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n555), .A2(G48), .A3(G543), .A4(new_n516), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n594), .A2(new_n596), .A3(new_n598), .A4(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n544), .A2(G85), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI221_X1 g178(.A(new_n601), .B1(new_n514), .B2(new_n602), .C1(new_n571), .C2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  OR3_X1    g180(.A1(G171), .A2(KEYINPUT79), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT79), .B1(G171), .B2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n544), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n548), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n556), .A2(G54), .B1(G651), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n616), .ZN(G284));
  OAI211_X1 g192(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n616), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n582), .A2(new_n586), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  XNOR2_X1  g196(.A(G297), .B(KEYINPUT80), .ZN(G280));
  XOR2_X1   g197(.A(KEYINPUT81), .B(G559), .Z(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(G860), .B2(new_n623), .ZN(G148));
  NAND2_X1  g199(.A1(new_n573), .A2(new_n605), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n610), .A2(new_n614), .A3(new_n623), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g204(.A1(new_n497), .A2(G135), .ZN(new_n630));
  OAI221_X1 g205(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n485), .C2(G111), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n490), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(G14), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n656), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n662), .A2(new_n663), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n667), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n675), .A2(new_n680), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n683));
  AOI211_X1 g258(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n686), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g268(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n689), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G29), .A2(G35), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G162), .B2(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G2090), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NOR2_X1   g277(.A1(G171), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G5), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1961), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT99), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n485), .A2(G103), .A3(G2104), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT94), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT25), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n497), .A2(G139), .ZN(new_n711));
  NAND2_X1  g286(.A1(G115), .A2(G2104), .ZN(new_n712));
  INV_X1    g287(.A(G127), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n501), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(new_n486), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT95), .Z(new_n716));
  NAND3_X1  g291(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT96), .ZN(new_n718));
  MUX2_X1   g293(.A(G33), .B(new_n718), .S(G29), .Z(new_n719));
  AOI211_X1 g294(.A(new_n701), .B(new_n707), .C1(G2072), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(G2072), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT97), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G32), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n497), .A2(G141), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT26), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n462), .A2(G105), .ZN(new_n728));
  INV_X1    g303(.A(G129), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n727), .B(new_n728), .C1(new_n490), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n724), .B1(new_n731), .B2(new_n723), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT27), .ZN(new_n733));
  INV_X1    g308(.A(G1996), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT31), .B(G11), .Z(new_n736));
  INV_X1    g311(.A(G28), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT98), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n635), .B2(new_n723), .ZN(new_n742));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G164), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2078), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n723), .B1(new_n746), .B2(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n746), .B2(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G160), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2084), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n742), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n702), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n702), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n704), .A2(new_n705), .ZN(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT92), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n615), .B2(new_n702), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT93), .B(G1348), .Z(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n751), .A2(new_n755), .A3(new_n756), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n702), .A2(G19), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n574), .B2(new_n702), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1341), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n723), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  OAI221_X1 g342(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n485), .C2(G116), .ZN(new_n768));
  INV_X1    g343(.A(G128), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n490), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n497), .B2(G140), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n767), .B1(new_n771), .B2(new_n723), .ZN(new_n772));
  INV_X1    g347(.A(G2067), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n759), .A2(new_n760), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n765), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n735), .A2(new_n762), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT102), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n702), .A2(G20), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n620), .B2(new_n702), .ZN(new_n782));
  INV_X1    g357(.A(G1956), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n700), .A2(G2090), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT103), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n720), .A2(new_n722), .A3(new_n777), .A4(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G23), .B(G288), .S(G16), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n702), .A2(G6), .ZN(new_n792));
  INV_X1    g367(.A(G305), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n702), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT88), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(KEYINPUT88), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT32), .B(G1981), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n702), .B1(new_n534), .B2(new_n537), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G22), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT89), .B(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  OAI221_X1 g382(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n485), .C2(G107), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G119), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n490), .ZN(new_n812));
  INV_X1    g387(.A(G131), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n496), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G29), .ZN(new_n816));
  INV_X1    g391(.A(G25), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G29), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT87), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n816), .B(new_n822), .C1(new_n817), .C2(G29), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n821), .B1(new_n819), .B2(new_n823), .ZN(new_n825));
  MUX2_X1   g400(.A(G24), .B(G290), .S(G16), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1986), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n800), .A2(new_n829), .A3(new_n805), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT90), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT90), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n807), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n807), .B(new_n834), .C1(new_n831), .C2(new_n832), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n788), .B1(new_n836), .B2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  INV_X1    g414(.A(new_n788), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(G150));
  NAND2_X1  g416(.A1(new_n544), .A2(G93), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(new_n514), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n844), .C1(new_n571), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n573), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n846), .A2(new_n573), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n616), .A2(G559), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n853), .B(new_n854), .Z(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n856), .A2(new_n857), .A3(G860), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n848), .A2(new_n849), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n858), .A2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(new_n634), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n815), .A2(new_n641), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n497), .A2(G142), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n489), .A2(G130), .A3(new_n486), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT105), .ZN(new_n868));
  OAI221_X1 g443(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n485), .C2(G118), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n812), .A2(new_n641), .A3(new_n814), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n865), .A2(new_n866), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n871), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n866), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n771), .B(new_n510), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n731), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n725), .B2(new_n730), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n717), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n718), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n872), .B(new_n875), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n875), .A2(new_n872), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n878), .A2(new_n879), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n884), .B(new_n880), .C1(new_n885), .C2(new_n718), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n864), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n864), .A3(new_n886), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g469(.A(new_n626), .B1(new_n850), .B2(new_n851), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n850), .A2(new_n626), .A3(new_n851), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n615), .A2(G299), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n610), .A2(new_n614), .B1(new_n582), .B2(new_n586), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n899), .A2(new_n900), .A3(new_n898), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n896), .B(new_n897), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n899), .B2(new_n900), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n616), .A2(new_n620), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n615), .A2(G299), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n897), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n906), .B(new_n909), .C1(new_n910), .C2(new_n895), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n904), .A2(new_n911), .A3(KEYINPUT110), .ZN(new_n915));
  AOI21_X1  g490(.A(G305), .B1(new_n534), .B2(new_n537), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n534), .A2(new_n537), .A3(G305), .ZN(new_n918));
  OR2_X1    g493(.A1(G290), .A2(G288), .ZN(new_n919));
  NAND2_X1  g494(.A1(G290), .A2(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n917), .B(new_n918), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n918), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n926), .A2(new_n916), .B1(KEYINPUT108), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n928), .B2(KEYINPUT109), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n930), .A3(new_n927), .A4(new_n931), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n914), .A2(new_n915), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n929), .A2(new_n915), .A3(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n859), .A2(new_n605), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n937), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(new_n903), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n901), .ZN(new_n944));
  XNOR2_X1  g519(.A(G171), .B(G286), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n852), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G286), .B(G301), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n850), .A3(new_n851), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n946), .A2(new_n909), .A3(new_n906), .A4(new_n948), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n944), .A2(new_n949), .B1(new_n950), .B2(KEYINPUT112), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n950), .A2(KEYINPUT112), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n928), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n908), .A3(new_n907), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n928), .A3(new_n950), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n942), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n950), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n954), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(new_n957), .A3(new_n942), .A4(new_n958), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT44), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT113), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n928), .B1(new_n951), .B2(new_n952), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n967), .B2(new_n959), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT44), .A4(new_n964), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n942), .B1(new_n960), .B2(new_n963), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n967), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G40), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n977), .B(new_n475), .C1(new_n486), .C2(new_n482), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n510), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OR3_X1    g560(.A1(new_n985), .A2(G1986), .A3(G290), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n771), .B(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n731), .B(G1996), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n815), .A2(new_n821), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n815), .A2(new_n821), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n988), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n986), .A2(new_n987), .B1(new_n992), .B2(new_n985), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n986), .A2(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n988), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n990), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n773), .B2(new_n771), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n993), .A2(new_n994), .B1(new_n997), .B2(new_n985), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n984), .A2(new_n734), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n988), .A2(new_n731), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n985), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT126), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1002), .B(KEYINPUT47), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n998), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT60), .ZN(new_n1010));
  INV_X1    g585(.A(new_n760), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n510), .B2(new_n979), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n482), .A2(new_n486), .ZN(new_n1014));
  INV_X1    g589(.A(new_n475), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(G40), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n510), .A2(new_n1012), .A3(new_n979), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(G160), .A2(G40), .A3(new_n979), .A4(new_n510), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(G2067), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n616), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1021), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n510), .A2(new_n979), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n978), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1018), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n615), .B(new_n1023), .C1(new_n1028), .C2(new_n1011), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1010), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1024), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n978), .A3(new_n734), .A4(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(G1341), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1031), .B1(new_n1039), .B2(new_n574), .ZN(new_n1040));
  AOI211_X1 g615(.A(KEYINPUT59), .B(new_n573), .C1(new_n1035), .C2(new_n1038), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR4_X1   g617(.A1(new_n1019), .A2(new_n615), .A3(KEYINPUT60), .A4(new_n1021), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1030), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1025), .A2(KEYINPUT118), .A3(new_n978), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1048), .A3(new_n1018), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n783), .ZN(new_n1050));
  NAND2_X1  g625(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(G299), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n980), .A2(new_n1016), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT121), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1034), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n582), .A2(new_n1052), .A3(new_n1053), .A4(new_n586), .ZN(new_n1060));
  AND4_X1   g635(.A1(new_n1050), .A2(new_n1055), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1050), .A2(new_n1059), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1045), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1050), .A2(new_n1059), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1050), .A2(new_n1055), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1044), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1061), .A2(new_n1022), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1062), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n534), .A2(G8), .A3(new_n537), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n534), .A2(KEYINPUT55), .A3(G8), .A4(new_n537), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(G2090), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1033), .A2(new_n978), .A3(new_n1034), .ZN(new_n1081));
  INV_X1    g656(.A(G1971), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1078), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n590), .A2(KEYINPUT116), .A3(G1976), .A4(new_n591), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(G8), .A3(new_n1020), .ZN(new_n1087));
  OAI211_X1 g662(.A(G87), .B(new_n529), .C1(new_n525), .C2(new_n526), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n591), .A2(G1976), .A3(new_n588), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT52), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1024), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1078), .B1(new_n1095), .B2(new_n978), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .A4(new_n1086), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1020), .A2(G8), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n599), .A2(new_n598), .A3(new_n593), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G1981), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(G305), .B2(G1981), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1102), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT117), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n599), .A2(new_n598), .ZN(new_n1108));
  INV_X1    g683(.A(G1981), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n594), .A4(new_n596), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT49), .A4(new_n1102), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1099), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1083), .B1(new_n1049), .B2(G2090), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G8), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1085), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n705), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1119));
  INV_X1    g694(.A(G2078), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1033), .A2(new_n978), .A3(new_n1120), .A4(new_n1034), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1056), .A2(KEYINPUT53), .A3(new_n1120), .A4(new_n1034), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G171), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1119), .A2(new_n1123), .A3(G301), .A4(new_n1124), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1118), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1081), .A2(new_n754), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(G168), .C1(G2084), .C2(new_n1079), .ZN(new_n1134));
  NAND2_X1  g709(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1135));
  OR2_X1    g710(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(G8), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1133), .B1(G2084), .B2(new_n1079), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(G8), .A3(G286), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1134), .A2(G8), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1137), .B(new_n1139), .C1(new_n1140), .C2(new_n1135), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1134), .A2(G8), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT123), .A3(KEYINPUT51), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1145), .A2(KEYINPUT124), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1072), .A2(new_n1132), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1099), .A2(new_n1113), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G288), .A2(G1976), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1113), .A2(new_n1150), .B1(new_n1109), .B2(new_n793), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1085), .A2(new_n1149), .B1(new_n1151), .B2(new_n1100), .ZN(new_n1152));
  NOR4_X1   g727(.A1(new_n1027), .A2(new_n1013), .A3(new_n1016), .A4(G2084), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1966), .B1(new_n1056), .B2(new_n1034), .ZN(new_n1154));
  OAI211_X1 g729(.A(G8), .B(G168), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1138), .A2(new_n1157), .A3(G8), .A4(G168), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1085), .A2(new_n1114), .A3(new_n1117), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1085), .A4(new_n1114), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1152), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1148), .A2(new_n1166), .A3(KEYINPUT125), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT125), .B1(new_n1148), .B2(new_n1166), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1147), .A2(KEYINPUT62), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1118), .A2(new_n1126), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1167), .A2(new_n1168), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT115), .B1(G290), .B2(G1986), .ZN(new_n1175));
  NAND2_X1  g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1175), .B(new_n1176), .Z(new_n1177));
  AOI21_X1  g752(.A(new_n985), .B1(new_n992), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1009), .B1(new_n1174), .B2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g754(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1181), .B1(new_n694), .B2(new_n695), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1182), .A2(KEYINPUT127), .ZN(new_n1183));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n1184), .B(new_n1181), .C1(new_n694), .C2(new_n695), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g760(.A(new_n893), .B(new_n1186), .C1(new_n974), .C2(new_n973), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


