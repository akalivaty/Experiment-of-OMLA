//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(G116), .B(G119), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT2), .B(G113), .Z(new_n190));
  OR2_X1    g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n190), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT30), .ZN(new_n194));
  XOR2_X1   g008(.A(G134), .B(G137), .Z(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G128), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(G146), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n197), .A2(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .A4(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n196), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT11), .B1(new_n208), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n211), .B2(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(KEYINPUT65), .A3(G137), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n209), .A2(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n209), .A2(new_n212), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n215), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n207), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n221), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n217), .B1(new_n216), .B2(new_n218), .ZN(new_n228));
  AND4_X1   g042(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n218), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n201), .A2(new_n202), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT0), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(KEYINPUT64), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n201), .A2(new_n202), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT0), .B(G128), .Z(new_n240));
  AOI22_X1  g054(.A1(new_n237), .A2(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n224), .A2(new_n225), .B1(new_n230), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n223), .A2(new_n219), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT67), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT67), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n204), .B1(G143), .B2(new_n200), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n239), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n248), .A2(new_n205), .B1(G131), .B2(new_n195), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n194), .B1(new_n242), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n230), .A2(new_n241), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(new_n194), .A3(new_n250), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n193), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n193), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n249), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n253), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G237), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G210), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT26), .ZN(new_n265));
  INV_X1    g079(.A(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n259), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n256), .A2(new_n269), .A3(KEYINPUT70), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n223), .A2(new_n219), .B1(G131), .B2(new_n226), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n240), .A2(new_n239), .ZN(new_n276));
  INV_X1    g090(.A(new_n238), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT64), .B1(new_n231), .B2(new_n234), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n258), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n225), .B1(new_n243), .B2(new_n249), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT30), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n254), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n283), .A2(new_n193), .B1(new_n268), .B2(KEYINPUT69), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n271), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n274), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  INV_X1    g101(.A(new_n267), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n253), .A2(new_n250), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n193), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n291), .B2(new_n259), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n289), .B1(new_n290), .B2(new_n193), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n292), .B2(new_n293), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n288), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n286), .A2(new_n287), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n287), .B1(new_n286), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT32), .B(new_n187), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n256), .A2(new_n259), .ZN(new_n304));
  OR3_X1    g118(.A1(new_n304), .A2(KEYINPUT73), .A3(new_n267), .ZN(new_n305));
  OR3_X1    g119(.A1(new_n294), .A2(new_n296), .A3(new_n288), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT73), .B1(new_n304), .B2(new_n267), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT75), .B(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n193), .B1(new_n280), .B2(new_n281), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n259), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT28), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n314), .A2(new_n295), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n288), .A2(new_n307), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT74), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n311), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G472), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n302), .A2(new_n303), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n310), .B2(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n246), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G128), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n329), .A3(new_n332), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n328), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n331), .B2(G128), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n332), .B(new_n338), .C1(new_n330), .C2(new_n337), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G110), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n335), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n327), .B1(new_n342), .B2(new_n333), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n343), .B(new_n344), .C1(G110), .C2(new_n339), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G125), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G140), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT77), .A3(KEYINPUT16), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT16), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n347), .A3(G125), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n350), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(new_n353), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(new_n200), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n351), .A2(new_n200), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n346), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n334), .A2(new_n335), .A3(new_n328), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n339), .A2(G110), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n200), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n358), .A2(new_n200), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n364), .B(new_n365), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G137), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT79), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n361), .B1(new_n341), .B2(new_n345), .ZN(new_n376));
  INV_X1    g190(.A(new_n369), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n378), .A3(new_n310), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n326), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT81), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n326), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n378), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT82), .B1(new_n374), .B2(new_n378), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n326), .A2(G902), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT83), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n385), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n324), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G221), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT9), .B(G234), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G902), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G104), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT3), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n405));
  INV_X1    g219(.A(G107), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT85), .A2(G107), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT86), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT86), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n404), .A2(new_n407), .A3(new_n411), .A4(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(G104), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT3), .ZN(new_n414));
  AOI21_X1  g228(.A(G101), .B1(new_n403), .B2(G107), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n410), .A2(new_n412), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n409), .A2(KEYINPUT86), .B1(KEYINPUT3), .B2(new_n413), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(KEYINPUT87), .A3(new_n412), .A4(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n403), .A2(G107), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n410), .A2(new_n412), .A3(new_n414), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n424), .B2(G101), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n422), .A3(G101), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n241), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n407), .A2(new_n408), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n403), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n266), .B1(new_n430), .B2(new_n413), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n418), .B2(new_n420), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n248), .A2(new_n205), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT10), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n239), .B1(new_n247), .B2(new_n233), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n205), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT10), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n275), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n432), .B2(new_n433), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n437), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n432), .A2(new_n441), .A3(new_n433), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT88), .B(new_n230), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT12), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT90), .B(new_n230), .C1(new_n444), .C2(new_n445), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n440), .B(new_n448), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G140), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT84), .ZN(new_n457));
  INV_X1    g271(.A(G227), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n457), .B(new_n459), .Z(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n446), .A2(new_n447), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n451), .A3(new_n450), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n463), .A2(KEYINPUT91), .A3(new_n440), .A4(new_n448), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n440), .A2(new_n460), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT92), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n435), .A2(new_n468), .A3(new_n439), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n428), .A2(new_n434), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT93), .B1(new_n470), .B2(new_n438), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n275), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n440), .B2(new_n460), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n467), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n460), .B1(new_n453), .B2(new_n454), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n475), .B1(new_n480), .B2(new_n464), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT94), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(G469), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G469), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(new_n401), .ZN(new_n485));
  INV_X1    g299(.A(new_n466), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n463), .A2(new_n486), .A3(new_n448), .ZN(new_n487));
  INV_X1    g301(.A(new_n440), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n461), .B1(new_n472), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n311), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n490), .B2(new_n484), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n402), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n433), .A2(new_n349), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n279), .B2(new_n349), .ZN(new_n494));
  INV_X1    g308(.A(G224), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n496), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(KEYINPUT7), .B2(new_n496), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n427), .A2(new_n193), .ZN(new_n501));
  INV_X1    g315(.A(G116), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT5), .ZN(new_n504));
  OAI221_X1 g318(.A(G113), .B1(G119), .B2(new_n503), .C1(new_n188), .C2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(new_n192), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n426), .A2(new_n501), .B1(new_n432), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G122), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(KEYINPUT8), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n432), .A2(new_n506), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n432), .A2(new_n506), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n496), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n500), .A2(new_n509), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n401), .ZN(new_n516));
  INV_X1    g330(.A(new_n508), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n427), .A2(new_n193), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n421), .B2(new_n425), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n511), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT96), .B(KEYINPUT6), .Z(new_n521));
  OR2_X1    g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n507), .B2(new_n508), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n524), .A2(new_n525), .A3(new_n520), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(new_n524), .B2(new_n520), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n499), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n516), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G210), .B1(G237), .B2(G902), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n526), .A2(new_n527), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(KEYINPUT97), .A3(new_n499), .A4(new_n522), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT99), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n533), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n531), .B(KEYINPUT98), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT99), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n530), .A2(new_n539), .A3(new_n531), .A4(new_n533), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n260), .A2(new_n261), .A3(G214), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(new_n198), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT18), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(new_n218), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n351), .B(KEYINPUT101), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n360), .B1(new_n551), .B2(new_n200), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(KEYINPUT18), .A3(G131), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n553), .A2(KEYINPUT100), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(KEYINPUT100), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n550), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n548), .A2(new_n218), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n547), .A2(G131), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT19), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n351), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n551), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n359), .B(new_n559), .C1(new_n562), .C2(G146), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n564), .A2(KEYINPUT102), .ZN(new_n565));
  XNOR2_X1  g379(.A(G113), .B(G122), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n403), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n564), .B2(KEYINPUT102), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n547), .A2(KEYINPUT17), .A3(G131), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n559), .B2(KEYINPUT17), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT103), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n367), .B2(new_n368), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n359), .A2(KEYINPUT103), .A3(new_n366), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n556), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n565), .A2(new_n568), .B1(new_n576), .B2(new_n567), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT20), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n565), .A2(new_n568), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n567), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n578), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n576), .A2(new_n567), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n576), .A2(new_n567), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n401), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n580), .A2(new_n585), .B1(new_n588), .B2(G475), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n502), .A2(G122), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n406), .B1(new_n590), .B2(KEYINPUT14), .ZN(new_n591));
  XNOR2_X1  g405(.A(G116), .B(G122), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n593), .B2(KEYINPUT14), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n233), .A2(G143), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT104), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n246), .A2(G143), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n596), .A2(new_n208), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n208), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  OAI221_X1 g413(.A(new_n594), .B1(new_n429), .B2(new_n593), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT13), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n596), .A2(new_n601), .B1(G143), .B2(new_n246), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n208), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n429), .B(new_n592), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n600), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n399), .A2(new_n325), .A3(G953), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n600), .B(new_n608), .C1(new_n604), .C2(new_n606), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT105), .A3(new_n611), .ZN(new_n612));
  OR3_X1    g426(.A1(new_n607), .A2(KEYINPUT105), .A3(new_n609), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n310), .ZN(new_n614));
  OAI21_X1  g428(.A(G478), .B1(KEYINPUT106), .B2(KEYINPUT15), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(KEYINPUT106), .B2(KEYINPUT15), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n614), .B(new_n616), .Z(new_n617));
  NAND2_X1  g431(.A1(new_n589), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G952), .ZN(new_n619));
  AOI211_X1 g433(.A(G953), .B(new_n619), .C1(G234), .C2(G237), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n261), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT21), .B(G898), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n397), .A2(new_n492), .A3(new_n545), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n612), .A2(new_n613), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n610), .A2(KEYINPUT33), .A3(new_n611), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G478), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n311), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n631), .A2(new_n633), .B1(new_n632), .B2(new_n614), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n589), .A2(new_n634), .A3(new_n623), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n531), .B1(new_n530), .B2(new_n533), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n543), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT107), .ZN(new_n639));
  INV_X1    g453(.A(new_n531), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n536), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n534), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n543), .A4(new_n635), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n310), .B1(new_n298), .B2(new_n299), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G472), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n396), .A3(new_n300), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n492), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AOI21_X1  g466(.A(new_n544), .B1(new_n641), .B2(new_n534), .ZN(new_n653));
  INV_X1    g467(.A(new_n623), .ZN(new_n654));
  INV_X1    g468(.A(new_n617), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n589), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n492), .A2(new_n649), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  AND2_X1   g475(.A1(new_n647), .A2(new_n300), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n385), .A2(new_n387), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n363), .A2(new_n369), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n375), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n394), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n624), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n492), .A2(new_n545), .A3(new_n662), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AND2_X1   g486(.A1(new_n663), .A2(new_n667), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n402), .B(new_n673), .C1(new_n483), .C2(new_n491), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n621), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT108), .ZN(new_n677));
  INV_X1    g491(.A(new_n620), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(KEYINPUT108), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n656), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n324), .A2(new_n653), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XNOR2_X1  g499(.A(new_n680), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n492), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT40), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT38), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n541), .A2(KEYINPUT109), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n541), .A2(KEYINPUT109), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n541), .A2(KEYINPUT109), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(KEYINPUT38), .A3(new_n690), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n284), .A2(new_n271), .B1(new_n288), .B2(new_n313), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n302), .A2(new_n303), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n589), .A2(new_n617), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n668), .A2(new_n700), .A3(new_n544), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n695), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n688), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n198), .ZN(G45));
  INV_X1    g518(.A(new_n589), .ZN(new_n705));
  INV_X1    g519(.A(new_n634), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n681), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n324), .A2(new_n653), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n674), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(new_n402), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n490), .B2(new_n713), .ZN(new_n714));
  AOI211_X1 g528(.A(KEYINPUT110), .B(new_n311), .C1(new_n487), .C2(new_n489), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n487), .A2(new_n489), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n310), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT110), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n490), .A2(new_n713), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n719), .A2(new_n720), .A3(G469), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n490), .A2(new_n484), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n712), .A2(new_n716), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n397), .A2(new_n645), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT41), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G113), .ZN(G15));
  NAND3_X1  g541(.A1(new_n397), .A2(new_n724), .A3(new_n658), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NAND4_X1  g543(.A1(new_n724), .A2(new_n324), .A3(new_n653), .A4(new_n669), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NAND3_X1  g545(.A1(new_n653), .A2(new_n654), .A3(new_n699), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n286), .B1(new_n267), .B2(new_n315), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n187), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n647), .A2(new_n396), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n724), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  AND4_X1   g552(.A1(new_n647), .A2(new_n668), .A3(new_n708), .A4(new_n734), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n724), .A2(new_n739), .A3(new_n653), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NOR2_X1   g555(.A1(new_n402), .A2(new_n544), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n535), .A2(new_n538), .A3(new_n540), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n491), .B1(new_n477), .B2(new_n484), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n324), .A3(new_n396), .A4(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n708), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n745), .A2(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n397), .A3(new_n708), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n750), .B1(new_n752), .B2(new_n749), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(G131), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G33));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n397), .A3(new_n682), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n478), .B(new_n475), .C1(new_n480), .C2(new_n464), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT94), .B1(new_n465), .B2(new_n476), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n484), .B1(new_n481), .B2(KEYINPUT45), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n485), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n723), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n765), .B(new_n485), .C1(new_n761), .C2(new_n762), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n712), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n706), .A2(new_n589), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n705), .A2(KEYINPUT43), .A3(new_n634), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n668), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n662), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT44), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(KEYINPUT44), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n541), .A2(new_n544), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n768), .A2(new_n778), .A3(new_n686), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND2_X1  g594(.A1(new_n767), .A2(KEYINPUT47), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n712), .C1(new_n764), .C2(new_n766), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n777), .A2(new_n396), .A3(new_n324), .A4(new_n746), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n787));
  INV_X1    g601(.A(new_n724), .ZN(new_n788));
  INV_X1    g602(.A(new_n653), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n771), .A2(new_n620), .A3(new_n770), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n735), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n619), .B(G953), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n302), .A2(new_n396), .A3(new_n303), .A4(new_n697), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(new_n678), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n788), .A2(new_n795), .A3(new_n777), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n705), .A3(new_n706), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n788), .A2(new_n777), .A3(new_n791), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT48), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n798), .A2(new_n799), .A3(new_n397), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n798), .B2(new_n397), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n793), .B(new_n797), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n693), .A2(new_n695), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n792), .A2(new_n724), .A3(new_n544), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT50), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n705), .A2(new_n706), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n796), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n647), .A2(new_n668), .A3(new_n734), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n798), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n809), .A2(new_n814), .A3(KEYINPUT51), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n716), .A2(new_n722), .A3(new_n723), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n402), .ZN(new_n817));
  OAI21_X1  g631(.A(G469), .B1(new_n477), .B2(new_n758), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n479), .A2(new_n482), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n758), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n765), .B1(new_n820), .B2(new_n485), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n723), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n782), .B1(new_n823), .B2(new_n712), .ZN(new_n824));
  INV_X1    g638(.A(new_n783), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n817), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n792), .A2(new_n776), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n802), .B1(new_n815), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n809), .A2(new_n814), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n824), .B2(new_n825), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n781), .A2(new_n832), .A3(new_n783), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n833), .A3(new_n817), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n830), .B1(new_n834), .B2(new_n827), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n829), .B1(new_n835), .B2(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n829), .B(new_n838), .C1(new_n835), .C2(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n841));
  OAI21_X1  g655(.A(new_n674), .B1(new_n683), .B2(new_n709), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n789), .A2(new_n700), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n668), .A2(new_n402), .A3(new_n681), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n698), .A3(new_n744), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n740), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n842), .A2(KEYINPUT52), .A3(new_n740), .A4(new_n845), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n618), .A2(new_n681), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n776), .A2(new_n324), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n674), .A2(new_n852), .B1(new_n739), .B2(new_n751), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n753), .A2(new_n853), .A3(new_n756), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n623), .B1(new_n707), .B2(new_n656), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n492), .A2(new_n545), .A3(new_n649), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n625), .A2(new_n670), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n397), .B(new_n724), .C1(new_n645), .C2(new_n658), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n730), .A3(new_n737), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n730), .A3(KEYINPUT114), .A4(new_n737), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n854), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n841), .B1(new_n850), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n848), .A2(new_n866), .A3(new_n849), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n847), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n857), .A2(new_n859), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n854), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n865), .A3(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n850), .A2(new_n863), .A3(new_n841), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n859), .A2(new_n860), .ZN(new_n874));
  INV_X1    g688(.A(new_n857), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n862), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n753), .A2(new_n853), .A3(new_n756), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT115), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n854), .A2(new_n861), .A3(new_n879), .A4(new_n862), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n880), .A3(new_n868), .A4(new_n867), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n873), .B1(new_n881), .B2(new_n869), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n872), .B1(new_n882), .B2(new_n865), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n787), .B1(new_n840), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n872), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n869), .ZN(new_n886));
  INV_X1    g700(.A(new_n873), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n888), .B2(KEYINPUT54), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(KEYINPUT120), .A3(new_n837), .A4(new_n839), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n619), .A2(new_n261), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n816), .B(KEYINPUT49), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n794), .A2(new_n544), .A3(new_n402), .A4(new_n769), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n803), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(G75));
  NOR2_X1   g710(.A1(new_n261), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n310), .B1(new_n864), .B2(new_n871), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(new_n640), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n532), .A2(new_n522), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n499), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n898), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n899), .A2(new_n907), .A3(new_n537), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n899), .B2(new_n537), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT122), .B(new_n906), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(G51));
  AOI21_X1  g728(.A(new_n865), .B1(new_n864), .B2(new_n871), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n885), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n485), .B(KEYINPUT57), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n717), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n899), .A2(new_n820), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n897), .B1(new_n919), .B2(new_n920), .ZN(G54));
  AND3_X1   g735(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n898), .B1(new_n922), .B2(new_n583), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n583), .B2(new_n922), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  NOR2_X1   g740(.A1(new_n630), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n898), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n889), .A2(new_n926), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n630), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n864), .B2(new_n871), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n666), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n898), .C1(new_n391), .C2(new_n934), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g751(.A1(new_n876), .A2(new_n261), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n622), .B2(new_n495), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n901), .B1(G898), .B2(new_n261), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  XNOR2_X1  g757(.A(new_n283), .B(new_n562), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n707), .A2(new_n656), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n397), .A2(new_n776), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n687), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n842), .A2(new_n740), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n703), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n950), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(KEYINPUT62), .C1(new_n688), .C2(new_n702), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n948), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n779), .A3(new_n785), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n945), .B1(new_n955), .B2(new_n261), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n952), .A2(new_n753), .A3(new_n756), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n768), .A2(new_n397), .A3(new_n686), .A4(new_n843), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n959), .A2(new_n779), .A3(new_n785), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n261), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(G900), .B2(new_n261), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n945), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n957), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n458), .B2(new_n675), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT125), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n957), .A2(new_n958), .A3(new_n964), .A4(new_n967), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(G72));
  NOR2_X1   g785(.A1(new_n304), .A2(new_n288), .ZN(new_n972));
  INV_X1    g786(.A(new_n876), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n954), .A2(new_n779), .A3(new_n785), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  AND3_X1   g790(.A1(new_n974), .A2(KEYINPUT126), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT126), .B1(new_n974), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n972), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n961), .B2(new_n876), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n288), .A3(new_n304), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n898), .ZN(new_n985));
  INV_X1    g799(.A(new_n976), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n305), .A2(new_n308), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n284), .A2(new_n271), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n985), .B1(new_n888), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n980), .A2(new_n982), .A3(new_n990), .ZN(G57));
endmodule


