

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G164), .A2(G1384), .ZN(n751) );
  AND2_X2 U549 ( .A1(n710), .A2(G1996), .ZN(n687) );
  AND2_X2 U550 ( .A1(n543), .A2(n542), .ZN(G164) );
  XNOR2_X1 U551 ( .A(n517), .B(n516), .ZN(n856) );
  NOR2_X1 U552 ( .A1(n690), .A2(n938), .ZN(n696) );
  XNOR2_X1 U553 ( .A(n709), .B(KEYINPUT29), .ZN(n715) );
  NAND2_X1 U554 ( .A1(n686), .A2(n751), .ZN(n727) );
  INV_X1 U555 ( .A(KEYINPUT64), .ZN(n515) );
  NOR2_X1 U556 ( .A1(n633), .A2(G651), .ZN(n643) );
  XNOR2_X1 U557 ( .A(n515), .B(KEYINPUT17), .ZN(n516) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n514), .ZN(n850) );
  NOR2_X1 U559 ( .A1(n633), .A2(n527), .ZN(n649) );
  NOR2_X1 U560 ( .A1(n521), .A2(n520), .ZN(G160) );
  AND2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n851) );
  NAND2_X1 U562 ( .A1(n851), .A2(G113), .ZN(n513) );
  INV_X1 U563 ( .A(G2105), .ZN(n514) );
  AND2_X1 U564 ( .A1(n514), .A2(G2104), .ZN(n854) );
  NAND2_X1 U565 ( .A1(G101), .A2(n854), .ZN(n511) );
  XOR2_X1 U566 ( .A(KEYINPUT23), .B(n511), .Z(n512) );
  NAND2_X1 U567 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U568 ( .A1(G125), .A2(n850), .ZN(n519) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NAND2_X1 U570 ( .A1(G137), .A2(n856), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U572 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  INV_X1 U573 ( .A(G651), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n649), .A2(G76), .ZN(n522) );
  XNOR2_X1 U575 ( .A(KEYINPUT68), .B(n522), .ZN(n525) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n646) );
  NAND2_X1 U577 ( .A1(n646), .A2(G89), .ZN(n523) );
  XNOR2_X1 U578 ( .A(KEYINPUT4), .B(n523), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U580 ( .A(KEYINPUT5), .B(n526), .ZN(n535) );
  XNOR2_X1 U581 ( .A(KEYINPUT6), .B(KEYINPUT70), .ZN(n533) );
  NAND2_X1 U582 ( .A1(n643), .A2(G51), .ZN(n531) );
  NOR2_X1 U583 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n528), .Z(n645) );
  NAND2_X1 U585 ( .A1(n645), .A2(G63), .ZN(n529) );
  XOR2_X1 U586 ( .A(KEYINPUT69), .B(n529), .Z(n530) );
  NAND2_X1 U587 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U588 ( .A(n533), .B(n532), .Z(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U590 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  XOR2_X1 U591 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U592 ( .A1(n856), .A2(G138), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G102), .A2(n854), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G114), .A2(n851), .ZN(n537) );
  AND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n850), .A2(G126), .ZN(n539) );
  XNOR2_X1 U597 ( .A(n539), .B(KEYINPUT90), .ZN(n540) );
  AND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G85), .A2(n646), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G72), .A2(n649), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G60), .A2(n645), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G47), .A2(n643), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U605 ( .A1(n549), .A2(n548), .ZN(G290) );
  XNOR2_X1 U606 ( .A(G2451), .B(G2435), .ZN(n559) );
  XOR2_X1 U607 ( .A(G2446), .B(KEYINPUT107), .Z(n551) );
  XNOR2_X1 U608 ( .A(G2454), .B(G2430), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n551), .B(n550), .ZN(n555) );
  XOR2_X1 U610 ( .A(KEYINPUT106), .B(G2427), .Z(n553) );
  XNOR2_X1 U611 ( .A(G1341), .B(G1348), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U613 ( .A(n555), .B(n554), .Z(n557) );
  XNOR2_X1 U614 ( .A(G2443), .B(G2438), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U616 ( .A(n559), .B(n558), .ZN(n560) );
  AND2_X1 U617 ( .A1(n560), .A2(G14), .ZN(G401) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  NAND2_X1 U621 ( .A1(G64), .A2(n645), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G52), .A2(n643), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT65), .B(n563), .Z(n568) );
  NAND2_X1 U625 ( .A1(G90), .A2(n646), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G77), .A2(n649), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n566), .Z(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U632 ( .A(G223), .ZN(n824) );
  NAND2_X1 U633 ( .A1(n824), .A2(G567), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U635 ( .A1(G56), .A2(n645), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U637 ( .A1(n646), .A2(G81), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G68), .A2(n649), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n643), .A2(G43), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n938) );
  INV_X1 U645 ( .A(G860), .ZN(n600) );
  OR2_X1 U646 ( .A1(n938), .A2(n600), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U649 ( .A1(G66), .A2(n645), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G92), .A2(n646), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G79), .A2(n649), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G54), .A2(n643), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U656 ( .A(KEYINPUT67), .B(KEYINPUT15), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n587), .B(n586), .ZN(n931) );
  OR2_X1 U658 ( .A1(n931), .A2(G868), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G65), .A2(n645), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G53), .A2(n643), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G91), .A2(n646), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G78), .A2(n649), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n705) );
  INV_X1 U667 ( .A(n705), .ZN(G299) );
  INV_X1 U668 ( .A(G868), .ZN(n667) );
  NOR2_X1 U669 ( .A1(G286), .A2(n667), .ZN(n596) );
  XOR2_X1 U670 ( .A(KEYINPUT71), .B(n596), .Z(n599) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT72), .B(n597), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n601), .A2(n931), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT16), .ZN(n603) );
  XOR2_X1 U677 ( .A(KEYINPUT73), .B(n603), .Z(G148) );
  NAND2_X1 U678 ( .A1(n931), .A2(G868), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G559), .A2(n604), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT74), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n938), .A2(G868), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G99), .A2(n854), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G111), .A2(n851), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n850), .A2(G123), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G135), .A2(n856), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U690 ( .A(KEYINPUT75), .B(n613), .Z(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n984) );
  XOR2_X1 U692 ( .A(n984), .B(G2096), .Z(n617) );
  XNOR2_X1 U693 ( .A(G2100), .B(KEYINPUT76), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(KEYINPUT77), .B(n618), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G80), .A2(n649), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G55), .A2(n643), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT80), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n646), .A2(G93), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G67), .A2(n645), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n623), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n666) );
  NAND2_X1 U706 ( .A1(G559), .A2(n931), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n628), .B(n938), .ZN(n663) );
  NOR2_X1 U708 ( .A1(G860), .A2(n663), .ZN(n629) );
  XOR2_X1 U709 ( .A(n666), .B(n629), .Z(G145) );
  NAND2_X1 U710 ( .A1(G49), .A2(n643), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n645), .A2(n632), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n633), .A2(G87), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G62), .A2(n645), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G88), .A2(n646), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G50), .A2(n643), .ZN(n638) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(n638), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n649), .A2(G75), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(G303) );
  INV_X1 U724 ( .A(G303), .ZN(G166) );
  NAND2_X1 U725 ( .A1(n643), .A2(G48), .ZN(n644) );
  XNOR2_X1 U726 ( .A(KEYINPUT82), .B(n644), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G61), .A2(n645), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G86), .A2(n646), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U733 ( .A(KEYINPUT81), .B(n653), .Z(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(G305) );
  XNOR2_X1 U735 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n657) );
  XNOR2_X1 U736 ( .A(G288), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U737 ( .A(n657), .B(n656), .ZN(n660) );
  XNOR2_X1 U738 ( .A(G166), .B(G305), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(n666), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n662) );
  XNOR2_X1 U741 ( .A(G290), .B(n705), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n872) );
  XNOR2_X1 U743 ( .A(n872), .B(n663), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n664), .A2(G868), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(KEYINPUT86), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XOR2_X1 U753 ( .A(KEYINPUT66), .B(G82), .Z(G220) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U756 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G108), .A2(n675), .ZN(n829) );
  NAND2_X1 U758 ( .A1(G567), .A2(n829), .ZN(n683) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n677) );
  XNOR2_X1 U760 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n676) );
  XNOR2_X1 U761 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U762 ( .A1(n678), .A2(G218), .ZN(n679) );
  XNOR2_X1 U763 ( .A(KEYINPUT88), .B(n679), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n680), .A2(G96), .ZN(n828) );
  NAND2_X1 U765 ( .A1(G2106), .A2(n828), .ZN(n681) );
  XOR2_X1 U766 ( .A(KEYINPUT89), .B(n681), .Z(n682) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n903) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U769 ( .A1(n903), .A2(n684), .ZN(n827) );
  NAND2_X1 U770 ( .A1(n827), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n784) );
  NOR2_X1 U772 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U773 ( .A1(n784), .A2(n685), .ZN(n928) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n750) );
  INV_X1 U775 ( .A(n750), .ZN(n686) );
  INV_X1 U776 ( .A(n727), .ZN(n710) );
  XOR2_X1 U777 ( .A(n687), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U778 ( .A1(n727), .A2(G1341), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n696), .A2(n931), .ZN(n695) );
  AND2_X1 U781 ( .A1(n727), .A2(G1348), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT99), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n710), .A2(G2067), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n698) );
  OR2_X1 U786 ( .A1(n931), .A2(n696), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n710), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT27), .ZN(n701) );
  AND2_X1 U790 ( .A1(G1956), .A2(n727), .ZN(n700) );
  NOR2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U792 ( .A1(n705), .A2(n704), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U794 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U795 ( .A(n706), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U796 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n710), .A2(G1961), .ZN(n712) );
  XOR2_X1 U798 ( .A(KEYINPUT25), .B(G2078), .Z(n909) );
  NOR2_X1 U799 ( .A1(n727), .A2(n909), .ZN(n711) );
  NOR2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n720) );
  NOR2_X1 U801 ( .A1(n720), .A2(G301), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n713), .B(KEYINPUT98), .ZN(n714) );
  NOR2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n725) );
  NAND2_X1 U804 ( .A1(G8), .A2(n727), .ZN(n800) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n800), .ZN(n738) );
  NOR2_X1 U806 ( .A1(n727), .A2(G2084), .ZN(n740) );
  XNOR2_X1 U807 ( .A(n740), .B(KEYINPUT97), .ZN(n716) );
  NAND2_X1 U808 ( .A1(G8), .A2(n716), .ZN(n717) );
  NOR2_X1 U809 ( .A1(n738), .A2(n717), .ZN(n718) );
  XOR2_X1 U810 ( .A(KEYINPUT30), .B(n718), .Z(n719) );
  NOR2_X1 U811 ( .A1(G168), .A2(n719), .ZN(n722) );
  AND2_X1 U812 ( .A1(G301), .A2(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U814 ( .A(n723), .B(KEYINPUT31), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n737) );
  INV_X1 U816 ( .A(n737), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n726), .A2(G286), .ZN(n733) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n800), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U821 ( .A(KEYINPUT102), .B(n730), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n731), .A2(G303), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U824 ( .A(KEYINPUT103), .B(n734), .Z(n735) );
  NAND2_X1 U825 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U826 ( .A(KEYINPUT32), .B(n736), .ZN(n746) );
  NOR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U828 ( .A(KEYINPUT100), .B(n739), .ZN(n743) );
  XOR2_X1 U829 ( .A(KEYINPUT97), .B(n740), .Z(n741) );
  NAND2_X1 U830 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U832 ( .A(KEYINPUT101), .B(n744), .Z(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n796) );
  NAND2_X1 U834 ( .A1(n928), .A2(n796), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n747), .B(KEYINPUT104), .ZN(n790) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n927) );
  INV_X1 U837 ( .A(n927), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n800), .A2(n748), .ZN(n788) );
  XNOR2_X1 U839 ( .A(G1981), .B(KEYINPUT105), .ZN(n749) );
  XNOR2_X1 U840 ( .A(n749), .B(G305), .ZN(n941) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n819) );
  XNOR2_X1 U842 ( .A(G2067), .B(KEYINPUT37), .ZN(n817) );
  NAND2_X1 U843 ( .A1(n854), .A2(G104), .ZN(n752) );
  XOR2_X1 U844 ( .A(KEYINPUT91), .B(n752), .Z(n754) );
  NAND2_X1 U845 ( .A1(G140), .A2(n856), .ZN(n753) );
  NAND2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U847 ( .A(KEYINPUT34), .B(n755), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n851), .A2(G116), .ZN(n756) );
  XNOR2_X1 U849 ( .A(n756), .B(KEYINPUT92), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G128), .A2(n850), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U852 ( .A(KEYINPUT35), .B(n759), .ZN(n760) );
  XNOR2_X1 U853 ( .A(KEYINPUT93), .B(n760), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U855 ( .A(KEYINPUT36), .B(n763), .ZN(n847) );
  NOR2_X1 U856 ( .A1(n817), .A2(n847), .ZN(n993) );
  NAND2_X1 U857 ( .A1(n819), .A2(n993), .ZN(n815) );
  NAND2_X1 U858 ( .A1(G129), .A2(n850), .ZN(n765) );
  NAND2_X1 U859 ( .A1(G117), .A2(n851), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n854), .A2(G105), .ZN(n766) );
  XOR2_X1 U862 ( .A(KEYINPUT38), .B(n766), .Z(n767) );
  NOR2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G141), .A2(n856), .ZN(n769) );
  NAND2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n865) );
  NAND2_X1 U866 ( .A1(G1996), .A2(n865), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G119), .A2(n850), .ZN(n772) );
  NAND2_X1 U868 ( .A1(G107), .A2(n851), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n854), .A2(G95), .ZN(n773) );
  XOR2_X1 U871 ( .A(KEYINPUT94), .B(n773), .Z(n774) );
  NOR2_X1 U872 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U873 ( .A1(G131), .A2(n856), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n866) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n866), .ZN(n778) );
  XOR2_X1 U876 ( .A(KEYINPUT95), .B(n778), .Z(n779) );
  NAND2_X1 U877 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U878 ( .A(KEYINPUT96), .B(n781), .Z(n994) );
  INV_X1 U879 ( .A(n994), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n819), .A2(n782), .ZN(n809) );
  NAND2_X1 U881 ( .A1(n815), .A2(n809), .ZN(n804) );
  INV_X1 U882 ( .A(n804), .ZN(n783) );
  NAND2_X1 U883 ( .A1(n941), .A2(n783), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n784), .A2(KEYINPUT33), .ZN(n785) );
  NOR2_X1 U885 ( .A1(n800), .A2(n785), .ZN(n786) );
  NOR2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n791) );
  AND2_X1 U887 ( .A1(n788), .A2(n791), .ZN(n789) );
  AND2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n793) );
  AND2_X1 U889 ( .A1(n791), .A2(KEYINPUT33), .ZN(n792) );
  NOR2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n806) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n794) );
  NAND2_X1 U892 ( .A1(G8), .A2(n794), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n797), .A2(n800), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XOR2_X1 U896 ( .A(n798), .B(KEYINPUT24), .Z(n799) );
  OR2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X2 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n808) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n935) );
  NAND2_X1 U902 ( .A1(n935), .A2(n819), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n822) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n865), .ZN(n980) );
  INV_X1 U905 ( .A(n809), .ZN(n812) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n866), .ZN(n985) );
  NOR2_X1 U908 ( .A1(n810), .A2(n985), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n980), .A2(n813), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n814), .B(KEYINPUT39), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n817), .A2(n847), .ZN(n999) );
  NAND2_X1 U914 ( .A1(n818), .A2(n999), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U920 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(G188) );
  XOR2_X1 U923 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(G325) );
  XNOR2_X1 U925 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NAND2_X1 U929 ( .A1(n850), .A2(G124), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n830), .B(KEYINPUT44), .ZN(n832) );
  NAND2_X1 U931 ( .A1(G112), .A2(n851), .ZN(n831) );
  NAND2_X1 U932 ( .A1(n832), .A2(n831), .ZN(n836) );
  NAND2_X1 U933 ( .A1(G100), .A2(n854), .ZN(n834) );
  NAND2_X1 U934 ( .A1(G136), .A2(n856), .ZN(n833) );
  NAND2_X1 U935 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U936 ( .A1(n836), .A2(n835), .ZN(G162) );
  XOR2_X1 U937 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n838) );
  XNOR2_X1 U938 ( .A(G164), .B(KEYINPUT46), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n984), .B(n839), .ZN(n849) );
  NAND2_X1 U941 ( .A1(G103), .A2(n854), .ZN(n841) );
  NAND2_X1 U942 ( .A1(G139), .A2(n856), .ZN(n840) );
  NAND2_X1 U943 ( .A1(n841), .A2(n840), .ZN(n846) );
  NAND2_X1 U944 ( .A1(G127), .A2(n850), .ZN(n843) );
  NAND2_X1 U945 ( .A1(G115), .A2(n851), .ZN(n842) );
  NAND2_X1 U946 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(KEYINPUT47), .B(n844), .Z(n845) );
  NOR2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n988) );
  XNOR2_X1 U949 ( .A(n847), .B(n988), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n864) );
  NAND2_X1 U951 ( .A1(G130), .A2(n850), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G118), .A2(n851), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n862) );
  NAND2_X1 U954 ( .A1(n854), .A2(G106), .ZN(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT112), .B(n855), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G142), .A2(n856), .ZN(n857) );
  XOR2_X1 U957 ( .A(KEYINPUT113), .B(n857), .Z(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n860), .B(KEYINPUT45), .Z(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n864), .B(n863), .Z(n870) );
  XNOR2_X1 U962 ( .A(G162), .B(n865), .ZN(n867) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U964 ( .A(G160), .B(n868), .ZN(n869) );
  XNOR2_X1 U965 ( .A(n870), .B(n869), .ZN(n871) );
  NOR2_X1 U966 ( .A1(G37), .A2(n871), .ZN(G395) );
  XOR2_X1 U967 ( .A(n872), .B(G286), .Z(n874) );
  XNOR2_X1 U968 ( .A(n931), .B(G171), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U970 ( .A(n875), .B(n938), .ZN(n876) );
  NOR2_X1 U971 ( .A1(G37), .A2(n876), .ZN(G397) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(G1961), .Z(n878) );
  XNOR2_X1 U973 ( .A(G1986), .B(G1956), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U975 ( .A(n879), .B(G2474), .Z(n881) );
  XNOR2_X1 U976 ( .A(G1996), .B(G1991), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n885) );
  XOR2_X1 U978 ( .A(G1976), .B(G1981), .Z(n883) );
  XNOR2_X1 U979 ( .A(G1966), .B(G1971), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U981 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U982 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(G229) );
  XOR2_X1 U984 ( .A(G2100), .B(G2096), .Z(n889) );
  XNOR2_X1 U985 ( .A(KEYINPUT42), .B(G2678), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U987 ( .A(KEYINPUT43), .B(G2090), .Z(n891) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2072), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U991 ( .A(G2084), .B(G2078), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(G227) );
  NOR2_X1 U993 ( .A1(G229), .A2(G227), .ZN(n896) );
  XNOR2_X1 U994 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G397), .A2(n897), .ZN(n900) );
  NOR2_X1 U996 ( .A1(n903), .A2(G401), .ZN(n898) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n898), .Z(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  NOR2_X1 U999 ( .A1(G395), .A2(n901), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(KEYINPUT116), .B(n902), .ZN(G308) );
  INV_X1 U1001 ( .A(G308), .ZN(G225) );
  INV_X1 U1002 ( .A(n903), .ZN(G319) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1004 ( .A(G2090), .B(G35), .Z(n920) );
  XNOR2_X1 U1005 ( .A(G1991), .B(G25), .ZN(n915) );
  XNOR2_X1 U1006 ( .A(G2067), .B(KEYINPUT119), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(n904), .B(G26), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(G1996), .B(G32), .ZN(n906) );
  XNOR2_X1 U1009 ( .A(G33), .B(G2072), .ZN(n905) );
  NOR2_X1 U1010 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(G27), .B(n909), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT120), .B(n910), .ZN(n911) );
  NOR2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1015 ( .A(KEYINPUT121), .B(n913), .ZN(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n916), .A2(G28), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT122), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT53), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(G34), .B(G2084), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(KEYINPUT54), .B(n921), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1024 ( .A(KEYINPUT55), .B(n924), .Z(n925) );
  NOR2_X1 U1025 ( .A1(G29), .A2(n925), .ZN(n977) );
  XNOR2_X1 U1026 ( .A(G16), .B(KEYINPUT56), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n926), .B(KEYINPUT123), .ZN(n949) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(G1956), .B(G299), .ZN(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(n931), .B(G1348), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(G1971), .A2(G303), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n947) );
  XNOR2_X1 U1036 ( .A(n938), .B(G1341), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G301), .B(G1961), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G168), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(n943), .B(KEYINPUT57), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n974) );
  XNOR2_X1 U1045 ( .A(G1348), .B(KEYINPUT59), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n950), .B(G4), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G20), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G1981), .B(G6), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1051 ( .A(KEYINPUT125), .B(G1341), .Z(n955) );
  XNOR2_X1 U1052 ( .A(G19), .B(n955), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT60), .B(n958), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G21), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G1961), .B(G5), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n966) );
  XOR2_X1 U1062 ( .A(G1986), .B(G24), .Z(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n967), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1066 ( .A(KEYINPUT61), .B(n970), .Z(n972) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT124), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1070 ( .A(KEYINPUT126), .B(n975), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n978), .ZN(n1007) );
  XOR2_X1 U1073 ( .A(G160), .B(G2084), .Z(n983) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT51), .B(n981), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G2072), .B(n988), .Z(n990) );
  XOR2_X1 U1081 ( .A(G164), .B(G2078), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT50), .B(n991), .Z(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT117), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(KEYINPUT52), .B(n1001), .ZN(n1003) );
  INV_X1 U1090 ( .A(KEYINPUT55), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(G29), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(n1005), .B(KEYINPUT118), .Z(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(KEYINPUT127), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1009), .ZN(G311) );
  INV_X1 U1097 ( .A(G311), .ZN(G150) );
endmodule

