

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  INV_X1 U319 ( .A(n373), .ZN(n374) );
  XNOR2_X1 U320 ( .A(n409), .B(n408), .ZN(n504) );
  XNOR2_X1 U321 ( .A(n573), .B(KEYINPUT41), .ZN(n558) );
  INV_X1 U322 ( .A(n558), .ZN(n545) );
  AND2_X1 U323 ( .A1(G226GAT), .A2(G233GAT), .ZN(n287) );
  XNOR2_X1 U324 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n461) );
  XNOR2_X1 U325 ( .A(n462), .B(n461), .ZN(n564) );
  XNOR2_X1 U326 ( .A(n348), .B(G197GAT), .ZN(n373) );
  XNOR2_X1 U327 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U328 ( .A(n351), .B(n287), .ZN(n352) );
  XNOR2_X1 U329 ( .A(n407), .B(KEYINPUT100), .ZN(n408) );
  XNOR2_X1 U330 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U331 ( .A(n353), .B(n352), .ZN(n355) );
  INV_X1 U332 ( .A(G190GAT), .ZN(n467) );
  XNOR2_X1 U333 ( .A(KEYINPUT38), .B(n443), .ZN(n489) );
  XNOR2_X1 U334 ( .A(n467), .B(KEYINPUT58), .ZN(n468) );
  XNOR2_X1 U335 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U336 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n447), .B(n446), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n289) );
  XNOR2_X1 U339 ( .A(G211GAT), .B(G78GAT), .ZN(n288) );
  XNOR2_X1 U340 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U341 ( .A(n290), .B(G64GAT), .Z(n292) );
  XOR2_X1 U342 ( .A(G1GAT), .B(G8GAT), .Z(n413) );
  XNOR2_X1 U343 ( .A(n413), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n295) );
  XOR2_X1 U345 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n294) );
  XNOR2_X1 U346 ( .A(G71GAT), .B(G57GAT), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n429) );
  XOR2_X1 U348 ( .A(n295), .B(n429), .Z(n297) );
  XOR2_X1 U349 ( .A(G15GAT), .B(G127GAT), .Z(n338) );
  XOR2_X1 U350 ( .A(G22GAT), .B(G155GAT), .Z(n369) );
  XNOR2_X1 U351 ( .A(n338), .B(n369), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U353 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n299) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U356 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n303) );
  XNOR2_X1 U358 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n304), .B(KEYINPUT77), .ZN(n305) );
  XOR2_X1 U361 ( .A(n306), .B(n305), .Z(n562) );
  XOR2_X1 U362 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n308) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(KEYINPUT68), .B(n309), .Z(n423) );
  XOR2_X1 U366 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n311) );
  XNOR2_X1 U367 ( .A(KEYINPUT75), .B(KEYINPUT64), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n423), .B(n312), .ZN(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT10), .B(KEYINPUT76), .Z(n314) );
  XNOR2_X1 U371 ( .A(G218GAT), .B(G92GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U373 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n316) );
  XNOR2_X1 U374 ( .A(G134GAT), .B(G106GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U376 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U377 ( .A(G50GAT), .B(G162GAT), .Z(n370) );
  XOR2_X1 U378 ( .A(G99GAT), .B(G85GAT), .Z(n428) );
  XOR2_X1 U379 ( .A(G36GAT), .B(G190GAT), .Z(n351) );
  XOR2_X1 U380 ( .A(n428), .B(n351), .Z(n320) );
  NAND2_X1 U381 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n370), .B(n321), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U385 ( .A(n325), .B(n324), .Z(n532) );
  XOR2_X1 U386 ( .A(KEYINPUT36), .B(n532), .Z(n579) );
  XOR2_X1 U387 ( .A(KEYINPUT86), .B(G183GAT), .Z(n327) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n328) );
  XOR2_X1 U391 ( .A(n329), .B(n328), .Z(n354) );
  XOR2_X1 U392 ( .A(KEYINPUT85), .B(G99GAT), .Z(n331) );
  XNOR2_X1 U393 ( .A(G43GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U395 ( .A(G71GAT), .B(G176GAT), .Z(n333) );
  XNOR2_X1 U396 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n342) );
  XOR2_X1 U399 ( .A(G120GAT), .B(KEYINPUT0), .Z(n337) );
  XNOR2_X1 U400 ( .A(G113GAT), .B(G134GAT), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n398) );
  XOR2_X1 U402 ( .A(n398), .B(n338), .Z(n340) );
  NAND2_X1 U403 ( .A1(G227GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U406 ( .A(n354), .B(n343), .Z(n511) );
  XOR2_X1 U407 ( .A(G64GAT), .B(G92GAT), .Z(n345) );
  XNOR2_X1 U408 ( .A(G176GAT), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n432) );
  XOR2_X1 U410 ( .A(KEYINPUT95), .B(n432), .Z(n350) );
  XOR2_X1 U411 ( .A(G218GAT), .B(KEYINPUT21), .Z(n347) );
  XNOR2_X1 U412 ( .A(KEYINPUT88), .B(G211GAT), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U414 ( .A(G8GAT), .B(n373), .Z(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n353) );
  XOR2_X1 U416 ( .A(n355), .B(n354), .Z(n508) );
  OR2_X1 U417 ( .A1(n511), .A2(n508), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n356), .B(KEYINPUT96), .ZN(n376) );
  XOR2_X1 U419 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n358) );
  NAND2_X1 U420 ( .A1(G228GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U422 ( .A(n359), .B(G204GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(G106GAT), .B(G78GAT), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n360), .B(G148GAT), .ZN(n433) );
  XOR2_X1 U425 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n362) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n397) );
  XNOR2_X1 U428 ( .A(n433), .B(n397), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U430 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n366) );
  XNOR2_X1 U431 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U433 ( .A(n368), .B(n367), .Z(n372) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n375) );
  XOR2_X1 U436 ( .A(n375), .B(n374), .Z(n463) );
  NAND2_X1 U437 ( .A1(n376), .A2(n463), .ZN(n378) );
  INV_X1 U438 ( .A(KEYINPUT25), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n381) );
  INV_X1 U440 ( .A(n508), .ZN(n498) );
  XNOR2_X1 U441 ( .A(n498), .B(KEYINPUT27), .ZN(n402) );
  INV_X1 U442 ( .A(n511), .ZN(n521) );
  NOR2_X1 U443 ( .A1(n521), .A2(n463), .ZN(n379) );
  XOR2_X1 U444 ( .A(n379), .B(KEYINPUT26), .Z(n537) );
  INV_X1 U445 ( .A(n537), .ZN(n566) );
  NAND2_X1 U446 ( .A1(n402), .A2(n566), .ZN(n380) );
  NAND2_X1 U447 ( .A1(n381), .A2(n380), .ZN(n401) );
  XOR2_X1 U448 ( .A(G85GAT), .B(G162GAT), .Z(n383) );
  XNOR2_X1 U449 ( .A(G29GAT), .B(G148GAT), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U451 ( .A(KEYINPUT94), .B(G155GAT), .Z(n385) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(G127GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U454 ( .A(n387), .B(n386), .Z(n392) );
  XOR2_X1 U455 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n389) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U458 ( .A(KEYINPUT93), .B(n390), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U460 ( .A(G57GAT), .B(KEYINPUT92), .Z(n394) );
  XNOR2_X1 U461 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U463 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U465 ( .A(n400), .B(n399), .Z(n506) );
  NAND2_X1 U466 ( .A1(n401), .A2(n506), .ZN(n405) );
  INV_X1 U467 ( .A(n506), .ZN(n565) );
  NAND2_X1 U468 ( .A1(n565), .A2(n402), .ZN(n517) );
  NOR2_X1 U469 ( .A1(n521), .A2(n517), .ZN(n403) );
  XOR2_X1 U470 ( .A(n463), .B(KEYINPUT28), .Z(n520) );
  INV_X1 U471 ( .A(n520), .ZN(n514) );
  NAND2_X1 U472 ( .A1(n403), .A2(n514), .ZN(n404) );
  NAND2_X1 U473 ( .A1(n405), .A2(n404), .ZN(n472) );
  AND2_X1 U474 ( .A1(n579), .A2(n472), .ZN(n406) );
  AND2_X1 U475 ( .A1(n562), .A2(n406), .ZN(n409) );
  XNOR2_X1 U476 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n407) );
  XOR2_X1 U477 ( .A(G141GAT), .B(G22GAT), .Z(n411) );
  XNOR2_X1 U478 ( .A(G36GAT), .B(G50GAT), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U480 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U481 ( .A1(G229GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U483 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n417) );
  XNOR2_X1 U484 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U486 ( .A(n419), .B(n418), .Z(n425) );
  XOR2_X1 U487 ( .A(G15GAT), .B(G113GAT), .Z(n421) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(G197GAT), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U491 ( .A(n425), .B(n424), .Z(n540) );
  INV_X1 U492 ( .A(n540), .ZN(n568) );
  XOR2_X1 U493 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n427) );
  XNOR2_X1 U494 ( .A(G120GAT), .B(KEYINPUT74), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U496 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U500 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n435) );
  XNOR2_X1 U501 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n434) );
  XOR2_X1 U502 ( .A(n435), .B(n434), .Z(n436) );
  XOR2_X1 U503 ( .A(n441), .B(n440), .Z(n573) );
  NOR2_X1 U504 ( .A1(n568), .A2(n573), .ZN(n475) );
  NAND2_X1 U505 ( .A1(n504), .A2(n475), .ZN(n442) );
  XOR2_X1 U506 ( .A(KEYINPUT102), .B(n442), .Z(n443) );
  NAND2_X1 U507 ( .A1(n489), .A2(n521), .ZN(n447) );
  XOR2_X1 U508 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n445) );
  INV_X1 U509 ( .A(G43GAT), .ZN(n444) );
  XOR2_X1 U510 ( .A(KEYINPUT121), .B(n498), .Z(n460) );
  INV_X1 U511 ( .A(n562), .ZN(n576) );
  NOR2_X1 U512 ( .A1(n568), .A2(n558), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n448), .B(KEYINPUT46), .ZN(n449) );
  NOR2_X1 U514 ( .A1(n576), .A2(n449), .ZN(n450) );
  NAND2_X1 U515 ( .A1(n450), .A2(n532), .ZN(n452) );
  INV_X1 U516 ( .A(KEYINPUT47), .ZN(n451) );
  XNOR2_X1 U517 ( .A(n452), .B(n451), .ZN(n458) );
  NAND2_X1 U518 ( .A1(n579), .A2(n576), .ZN(n453) );
  XNOR2_X1 U519 ( .A(n453), .B(KEYINPUT110), .ZN(n454) );
  XNOR2_X1 U520 ( .A(n454), .B(KEYINPUT45), .ZN(n455) );
  NOR2_X1 U521 ( .A1(n573), .A2(n455), .ZN(n456) );
  NAND2_X1 U522 ( .A1(n456), .A2(n568), .ZN(n457) );
  NAND2_X1 U523 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n459), .B(KEYINPUT48), .ZN(n519) );
  NAND2_X1 U525 ( .A1(n460), .A2(n519), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n506), .A2(n463), .ZN(n464) );
  OR2_X1 U527 ( .A1(n564), .A2(n464), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n465), .B(KEYINPUT55), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n466), .A2(n521), .ZN(n561) );
  NOR2_X1 U530 ( .A1(n532), .A2(n561), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n532), .A2(n576), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT83), .ZN(n471) );
  XNOR2_X1 U533 ( .A(KEYINPUT16), .B(n471), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT97), .ZN(n492) );
  NAND2_X1 U536 ( .A1(n475), .A2(n492), .ZN(n483) );
  NOR2_X1 U537 ( .A1(n506), .A2(n483), .ZN(n476) );
  XOR2_X1 U538 ( .A(G1GAT), .B(n476), .Z(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT34), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n508), .A2(n483), .ZN(n478) );
  XOR2_X1 U541 ( .A(KEYINPUT98), .B(n478), .Z(n479) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n511), .A2(n483), .ZN(n481) );
  XNOR2_X1 U544 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n482), .Z(G1326GAT) );
  NOR2_X1 U547 ( .A1(n514), .A2(n483), .ZN(n484) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n484), .Z(G1327GAT) );
  NAND2_X1 U549 ( .A1(n489), .A2(n565), .ZN(n487) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n485), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U552 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n498), .A2(n489), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n488), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n520), .A2(n489), .ZN(n490) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(n490), .ZN(G1331GAT) );
  NOR2_X1 U557 ( .A1(n540), .A2(n558), .ZN(n491) );
  XOR2_X1 U558 ( .A(KEYINPUT105), .B(n491), .Z(n505) );
  NAND2_X1 U559 ( .A1(n492), .A2(n505), .ZN(n493) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(n493), .Z(n501) );
  NAND2_X1 U561 ( .A1(n501), .A2(n565), .ZN(n497) );
  XOR2_X1 U562 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n495) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n494) );
  XNOR2_X1 U564 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n501), .A2(n498), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n499), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n501), .A2(n521), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U571 ( .A1(n520), .A2(n501), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n505), .A2(n504), .ZN(n513) );
  NOR2_X1 U574 ( .A1(n506), .A2(n513), .ZN(n507) );
  XOR2_X1 U575 ( .A(G85GAT), .B(n507), .Z(G1336GAT) );
  NOR2_X1 U576 ( .A1(n508), .A2(n513), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(G1337GAT) );
  NOR2_X1 U579 ( .A1(n511), .A2(n513), .ZN(n512) );
  XOR2_X1 U580 ( .A(G99GAT), .B(n512), .Z(G1338GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(n515), .Z(n516) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT112), .ZN(n525) );
  INV_X1 U585 ( .A(n517), .ZN(n518) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n538) );
  NOR2_X1 U587 ( .A1(n520), .A2(n538), .ZN(n522) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT111), .B(n523), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n540), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT113), .Z(n527) );
  NAND2_X1 U593 ( .A1(n533), .A2(n545), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n576), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n535) );
  INV_X1 U601 ( .A(n532), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n533), .A2(n551), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n536), .Z(G1343GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(KEYINPUT116), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n552), .A2(n540), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n541), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U612 ( .A(KEYINPUT52), .B(n544), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n552), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n549) );
  NAND2_X1 U616 ( .A1(n576), .A2(n552), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n568), .A2(n561), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(n560) );
  NOR2_X1 U627 ( .A1(n558), .A2(n561), .ZN(n559) );
  XOR2_X1 U628 ( .A(n560), .B(n559), .Z(G1349GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n572) );
  NOR2_X1 U633 ( .A1(n568), .A2(n572), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U638 ( .A(n572), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U642 ( .A1(n580), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n582) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

