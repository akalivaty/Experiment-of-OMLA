//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G101), .B1(new_n190), .B2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT5), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT2), .B(G113), .Z(new_n202));
  AOI22_X1  g016(.A1(new_n196), .A2(new_n201), .B1(new_n202), .B2(new_n195), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT76), .A2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT76), .A2(G107), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(G104), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n191), .B2(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n192), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n194), .A2(new_n203), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT81), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n202), .A2(new_n195), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n195), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(new_n209), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G101), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n210), .B1(new_n207), .B2(new_n209), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n220), .A2(KEYINPUT77), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT77), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n218), .B2(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(KEYINPUT77), .A3(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(KEYINPUT80), .A3(new_n216), .A4(new_n219), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n213), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(G110), .B(G122), .Z(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n188), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n226), .A2(new_n231), .ZN(new_n236));
  INV_X1    g050(.A(new_n213), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n233), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n188), .A3(new_n233), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT0), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n251), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n242), .A2(G146), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT64), .B(G143), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n257), .B(new_n252), .C1(new_n258), .C2(new_n246), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT72), .B(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n242), .B2(G146), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n247), .A2(new_n248), .B1(G128), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n251), .A2(KEYINPUT1), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n257), .B(new_n266), .C1(new_n258), .C2(new_n246), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G125), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G224), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n275), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n262), .B2(new_n272), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n240), .A2(new_n241), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n275), .A2(KEYINPUT7), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n276), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n275), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR3_X1    g098(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n210), .B1(new_n285), .B2(new_n192), .ZN(new_n286));
  INV_X1    g100(.A(new_n211), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n203), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n233), .A2(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n233), .A2(KEYINPUT8), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n196), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n195), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n201), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G116), .ZN(new_n298));
  OAI21_X1  g112(.A(G113), .B1(new_n298), .B2(KEYINPUT5), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT83), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n215), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n286), .A2(new_n287), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n291), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n234), .B2(new_n232), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n284), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n280), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n280), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n187), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT11), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G137), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(G137), .ZN(new_n318));
  INV_X1    g132(.A(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT11), .A3(G134), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G131), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n317), .A2(new_n320), .A3(new_n323), .A4(new_n318), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n251), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n246), .B1(new_n243), .B2(new_n245), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(new_n256), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n267), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n211), .A3(new_n194), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n265), .B(new_n267), .C1(new_n286), .C2(new_n287), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n260), .B(new_n219), .C1(new_n222), .C2(new_n223), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n268), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n326), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G140), .ZN(new_n341));
  INV_X1    g155(.A(G953), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(G227), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n341), .B(new_n343), .Z(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n325), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n348), .B2(new_n340), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n313), .B(new_n314), .C1(new_n346), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(G469), .A2(G902), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(KEYINPUT79), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n340), .A2(new_n353), .A3(new_n344), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n344), .ZN(new_n356));
  INV_X1    g170(.A(new_n340), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n335), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n350), .B(new_n351), .C1(new_n359), .C2(new_n313), .ZN(new_n360));
  INV_X1    g174(.A(G221), .ZN(new_n361));
  XOR2_X1   g175(.A(KEYINPUT9), .B(G234), .Z(new_n362));
  AOI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(new_n314), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n312), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n258), .B2(new_n251), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n243), .A2(new_n245), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT92), .A3(G128), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n251), .A2(G143), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n372), .A2(new_n316), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n316), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n198), .A2(KEYINPUT14), .A3(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(G116), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(G107), .B(new_n375), .C1(new_n377), .C2(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n189), .A2(new_n376), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n316), .B1(new_n371), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n372), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n372), .A2(new_n382), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n189), .B(new_n376), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n362), .A2(G217), .A3(new_n342), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n388), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n380), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n395));
  OAI21_X1  g209(.A(G478), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT94), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(new_n314), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G902), .B1(new_n389), .B2(new_n391), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n396), .A2(KEYINPUT94), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT95), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n398), .B(new_n403), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G475), .ZN(new_n406));
  INV_X1    g220(.A(G237), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n407), .A2(new_n342), .A3(G143), .A4(G214), .ZN(new_n408));
  INV_X1    g222(.A(G214), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n409), .A2(G237), .A3(G953), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT85), .B(new_n408), .C1(new_n258), .C2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n408), .A2(KEYINPUT85), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(KEYINPUT86), .A3(new_n412), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n415), .A2(KEYINPUT18), .A3(new_n416), .A4(G131), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n413), .B1(new_n418), .B2(new_n323), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT87), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT73), .B1(new_n261), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(G125), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(G140), .C1(new_n270), .C2(new_n271), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G146), .ZN(new_n427));
  XOR2_X1   g241(.A(G125), .B(G140), .Z(new_n428));
  OR2_X1    g242(.A1(new_n428), .A2(G146), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n413), .B(new_n431), .C1(new_n418), .C2(new_n323), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n417), .A2(new_n420), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n411), .A2(G131), .A3(new_n412), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n413), .A2(new_n323), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT17), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n411), .A2(KEYINPUT88), .A3(G131), .A4(new_n412), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT90), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n437), .B2(new_n440), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT16), .A4(new_n423), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT16), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n261), .A2(new_n445), .A3(new_n421), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(G146), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(G146), .B1(new_n444), .B2(new_n446), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n443), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n434), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(G113), .B(G122), .Z(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT89), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(G104), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n451), .B(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n406), .B1(new_n456), .B2(new_n314), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n441), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n441), .A2(new_n458), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n450), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n455), .A3(new_n433), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n437), .A2(new_n440), .A3(new_n438), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n426), .A2(KEYINPUT19), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(KEYINPUT19), .B2(new_n428), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(new_n447), .C1(new_n465), .C2(G146), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n455), .B1(new_n466), .B2(new_n433), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n470));
  NOR2_X1   g284(.A1(G475), .A2(G902), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(KEYINPUT91), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n467), .B1(new_n451), .B2(new_n455), .ZN(new_n475));
  INV_X1    g289(.A(new_n471), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT20), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n478));
  AOI211_X1 g292(.A(KEYINPUT20), .B(new_n476), .C1(new_n462), .C2(new_n468), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n405), .B(new_n457), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G952), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  NAND2_X1  g297(.A1(G234), .A2(G237), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT21), .B(G898), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(G902), .A3(G953), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n366), .A2(new_n481), .A3(KEYINPUT96), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n490));
  INV_X1    g304(.A(new_n187), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n280), .A2(new_n308), .ZN(new_n492));
  INV_X1    g306(.A(new_n309), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n280), .A2(new_n308), .A3(new_n309), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n365), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n474), .A2(new_n480), .ZN(new_n499));
  INV_X1    g313(.A(new_n405), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n456), .A2(new_n314), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G475), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n499), .A2(new_n488), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n490), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT71), .B1(new_n297), .B2(G128), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(KEYINPUT23), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(KEYINPUT23), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n507), .C1(G119), .C2(new_n251), .ZN(new_n508));
  XNOR2_X1  g322(.A(G119), .B(G128), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT24), .B(G110), .Z(new_n510));
  AOI22_X1  g324(.A1(new_n508), .A2(G110), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n448), .B2(new_n449), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT74), .B(G110), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n508), .A2(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n447), .A3(new_n429), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT22), .B(G137), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT75), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n342), .A2(G221), .A3(G234), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n512), .A2(new_n515), .A3(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT25), .B1(new_n524), .B2(G902), .ZN(new_n525));
  INV_X1    g339(.A(G217), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(G234), .B2(new_n314), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n522), .A2(new_n528), .A3(new_n314), .A4(new_n523), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n527), .A2(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n407), .A2(new_n342), .A3(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n535), .A2(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n536), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n216), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n325), .A2(new_n255), .A3(new_n259), .ZN(new_n547));
  INV_X1    g361(.A(new_n318), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n316), .A2(G137), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n266), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n328), .A2(new_n256), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n324), .B(new_n550), .C1(new_n552), .C2(new_n264), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT65), .A3(KEYINPUT30), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT65), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(new_n553), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n546), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n547), .A2(new_n553), .A3(new_n546), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n545), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n546), .B1(new_n547), .B2(new_n553), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT28), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT68), .B1(new_n562), .B2(KEYINPUT28), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT67), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n544), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n540), .A2(new_n543), .A3(KEYINPUT67), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n547), .A2(new_n553), .A3(new_n546), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT68), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT28), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n565), .A2(new_n566), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT29), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n563), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n565), .A2(new_n566), .A3(new_n575), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n545), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n582), .B2(KEYINPUT29), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n563), .A2(new_n576), .A3(KEYINPUT69), .A4(new_n577), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G472), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n556), .B(new_n557), .C1(new_n547), .C2(new_n553), .ZN(new_n587));
  AND4_X1   g401(.A1(new_n547), .A2(new_n553), .A3(new_n558), .A4(new_n559), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n216), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n572), .A3(new_n544), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT31), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n570), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT31), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n589), .A2(new_n593), .A3(new_n572), .A4(new_n544), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n314), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n595), .A2(KEYINPUT32), .A3(new_n596), .A4(new_n314), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n586), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT70), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n586), .A2(new_n599), .A3(new_n603), .A4(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n534), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n489), .A2(new_n504), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n595), .A2(new_n314), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G472), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n597), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(new_n365), .A3(new_n534), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n187), .B(new_n488), .C1(new_n310), .C2(new_n311), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n399), .A2(G478), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n392), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n389), .A2(KEYINPUT97), .A3(new_n616), .A4(new_n391), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n615), .B1(new_n621), .B2(G478), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n499), .B2(new_n502), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  OAI21_X1  g440(.A(new_n502), .B1(new_n479), .B2(new_n473), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n500), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n614), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n516), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n532), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n530), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n610), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n489), .A2(new_n504), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT37), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(G110), .Z(G12));
  AOI21_X1  g453(.A(new_n635), .B1(new_n602), .B2(new_n604), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n487), .A2(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n485), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n627), .A2(new_n500), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n640), .A2(new_n366), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  AOI21_X1  g460(.A(new_n457), .B1(new_n474), .B2(new_n480), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n500), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n642), .B(KEYINPUT39), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n497), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n497), .A2(KEYINPUT98), .A3(new_n649), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n652), .A2(new_n655), .A3(new_n653), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n561), .A2(new_n562), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n562), .A2(new_n564), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n658), .A2(new_n544), .B1(new_n659), .B2(new_n570), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n660), .B2(G902), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n599), .A2(new_n600), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n657), .A2(new_n187), .A3(new_n635), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n494), .A2(new_n495), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT38), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  OR3_X1    g480(.A1(new_n656), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n258), .ZN(G45));
  AOI21_X1  g482(.A(new_n479), .B1(new_n477), .B2(new_n478), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n475), .A2(KEYINPUT91), .A3(KEYINPUT20), .A4(new_n476), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n502), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n622), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n642), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT99), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n671), .A2(new_n675), .A3(new_n672), .A4(new_n642), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n640), .A3(new_n366), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  OAI21_X1  g492(.A(new_n314), .B1(new_n346), .B2(new_n349), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n364), .A3(new_n350), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n612), .A2(new_n647), .A3(new_n622), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n605), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT100), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT41), .B(G113), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND2_X1  g500(.A1(new_n602), .A2(new_n604), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n612), .A2(new_n534), .ZN(new_n688));
  INV_X1    g502(.A(new_n681), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n312), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n628), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  INV_X1    g506(.A(new_n635), .ZN(new_n693));
  AOI22_X1  g507(.A1(G472), .A2(new_n585), .B1(new_n597), .B2(new_n598), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n603), .B1(new_n694), .B2(new_n600), .ZN(new_n695));
  INV_X1    g509(.A(new_n604), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n690), .B(new_n693), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT101), .B1(new_n697), .B2(new_n503), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n664), .A2(new_n187), .A3(new_n681), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n604), .B2(new_n602), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(new_n503), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n693), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n597), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n595), .A2(KEYINPUT102), .A3(new_n596), .A4(new_n314), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n608), .B2(G472), .ZN(new_n711));
  AOI211_X1 g525(.A(KEYINPUT103), .B(new_n596), .C1(new_n595), .C2(new_n314), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n688), .A2(new_n648), .A3(new_n713), .A4(new_n681), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR4_X1   g529(.A1(new_n709), .A2(new_n711), .A3(new_n712), .A4(new_n635), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n674), .A2(new_n676), .A3(new_n690), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n494), .A2(new_n187), .A3(new_n495), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n497), .A2(KEYINPUT104), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n365), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n605), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n674), .A2(new_n676), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n719), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n600), .A2(KEYINPUT105), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n600), .A2(KEYINPUT105), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n694), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n534), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n674), .A3(new_n724), .A4(new_n676), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT106), .B1(new_n727), .B2(new_n733), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  INV_X1    g553(.A(new_n644), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n725), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n316), .ZN(G36));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n671), .A2(new_n622), .B1(KEYINPUT107), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n647), .A2(new_n672), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n610), .A3(new_n693), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n720), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n359), .B(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G469), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n351), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(G469), .C1(new_n756), .C2(G902), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n350), .A3(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n761), .A2(new_n364), .A3(new_n649), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n750), .A2(KEYINPUT108), .A3(new_n751), .A4(new_n752), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n755), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  INV_X1    g579(.A(new_n726), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n364), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT47), .B1(new_n761), .B2(new_n364), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n687), .A2(new_n731), .A3(new_n720), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n769), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  AND2_X1   g590(.A1(new_n680), .A2(new_n350), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT49), .Z(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n534), .A3(new_n745), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n662), .A2(new_n363), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n187), .A3(new_n666), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n401), .B(KEYINPUT111), .Z(new_n784));
  AND3_X1   g598(.A1(new_n647), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n647), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n614), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n671), .A2(new_n672), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT110), .B1(new_n788), .B2(new_n612), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n613), .A2(new_n623), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n791), .A3(new_n611), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n606), .A2(new_n637), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n741), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n721), .A2(new_n723), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n674), .A2(new_n676), .A3(new_n713), .A4(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n627), .A2(new_n643), .A3(new_n784), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n687), .A2(new_n797), .A3(new_n497), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n693), .A3(new_n751), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n642), .A2(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n642), .A2(KEYINPUT113), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n635), .A2(new_n662), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n496), .A3(new_n497), .A4(new_n648), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n677), .A2(new_n717), .A3(new_n645), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n794), .B(new_n800), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n683), .A2(new_n691), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n704), .A2(new_n714), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n734), .B2(new_n736), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n782), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n794), .A2(new_n800), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n782), .B1(new_n727), .B2(new_n733), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n805), .B(new_n806), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n811), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n809), .A2(new_n812), .A3(new_n782), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n813), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n819), .B1(KEYINPUT54), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n751), .A2(new_n681), .ZN(new_n823));
  OR4_X1    g637(.A1(new_n534), .A2(new_n823), .A3(new_n485), .A4(new_n662), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n824), .A2(new_n788), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n824), .A2(new_n671), .A3(new_n672), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n666), .A2(new_n491), .A3(new_n681), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n747), .A2(new_n713), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n534), .A3(new_n485), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT50), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n827), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n823), .A2(new_n485), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n747), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n716), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT116), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n751), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n767), .A2(new_n768), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n777), .A2(new_n363), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT114), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n826), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n845), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n751), .A3(new_n832), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n837), .A2(new_n850), .A3(KEYINPUT51), .A4(new_n841), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n848), .A2(new_n483), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n822), .A2(new_n825), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n832), .A2(new_n690), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n730), .A2(new_n731), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n839), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT48), .Z(new_n857));
  NOR3_X1   g671(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(G952), .A2(G953), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n781), .B1(new_n858), .B2(new_n859), .ZN(G75));
  NAND2_X1  g674(.A1(new_n482), .A2(G953), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT118), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n314), .B1(new_n813), .B2(new_n817), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT117), .B1(new_n863), .B2(G210), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n240), .A2(new_n241), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n279), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  AOI221_X4 g684(.A(KEYINPUT56), .B1(KEYINPUT117), .B2(new_n868), .C1(new_n863), .C2(G210), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT119), .B(new_n862), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(G51));
  INV_X1    g690(.A(new_n862), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n819), .A2(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n818), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n351), .B(KEYINPUT57), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n346), .A2(new_n349), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n863), .A2(G469), .A3(new_n756), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(G54));
  NAND3_X1  g701(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(new_n469), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n469), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n877), .B1(new_n889), .B2(new_n890), .ZN(G60));
  NAND2_X1  g705(.A1(new_n619), .A2(new_n620), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(G478), .A2(G902), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT59), .Z(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n880), .A2(new_n881), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n822), .B2(new_n895), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n897), .A2(new_n862), .A3(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT60), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n818), .A2(new_n633), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n818), .A2(new_n901), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n862), .B(new_n902), .C1(new_n903), .C2(new_n531), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g719(.A(new_n342), .B1(new_n486), .B2(G224), .ZN(new_n906));
  INV_X1    g720(.A(new_n811), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(new_n793), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n342), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT121), .ZN(new_n910));
  INV_X1    g724(.A(G898), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n866), .B1(new_n911), .B2(G953), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n910), .B(new_n912), .ZN(G69));
  NAND2_X1  g727(.A1(new_n555), .A2(new_n560), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n465), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n677), .A2(new_n645), .A3(new_n717), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n667), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n667), .A2(KEYINPUT62), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OR3_X1    g736(.A1(new_n785), .A2(new_n786), .A3(new_n623), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n605), .A3(new_n654), .A4(new_n751), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n764), .A3(new_n775), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n916), .B1(new_n926), .B2(new_n342), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n762), .A2(new_n496), .A3(new_n648), .A4(new_n855), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n764), .A2(new_n775), .A3(new_n917), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n738), .B1(new_n740), .B2(new_n725), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n342), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n342), .A2(G900), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT123), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n927), .B1(new_n934), .B2(new_n916), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n342), .B1(G227), .B2(G900), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n935), .B(new_n936), .Z(G72));
  XNOR2_X1  g751(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n596), .A2(new_n314), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n938), .B(new_n939), .Z(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n926), .B2(new_n908), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n658), .ZN(new_n944));
  OAI211_X1 g758(.A(KEYINPUT125), .B(new_n940), .C1(new_n926), .C2(new_n908), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n943), .A2(new_n544), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n940), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n563), .B2(new_n590), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT127), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n821), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n929), .A2(new_n908), .A3(new_n930), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n545), .B(new_n658), .C1(new_n952), .C2(new_n947), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n862), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n953), .B2(new_n862), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(G57));
endmodule


