

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U322 ( .A(KEYINPUT103), .B(KEYINPUT25), .ZN(n407) );
  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n466) );
  XOR2_X1 U324 ( .A(n581), .B(KEYINPUT41), .Z(n551) );
  XNOR2_X1 U325 ( .A(n457), .B(KEYINPUT37), .ZN(n529) );
  XOR2_X1 U326 ( .A(G36GAT), .B(n450), .Z(n290) );
  XOR2_X1 U327 ( .A(KEYINPUT87), .B(n377), .Z(n291) );
  XOR2_X1 U328 ( .A(n379), .B(KEYINPUT84), .Z(n292) );
  XNOR2_X1 U329 ( .A(n468), .B(KEYINPUT115), .ZN(n469) );
  XNOR2_X1 U330 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U331 ( .A1(n581), .A2(n472), .ZN(n473) );
  XNOR2_X1 U332 ( .A(n467), .B(n466), .ZN(n475) );
  NOR2_X1 U333 ( .A1(n530), .A2(n413), .ZN(n414) );
  XNOR2_X1 U334 ( .A(n447), .B(G134GAT), .ZN(n448) );
  INV_X1 U335 ( .A(KEYINPUT55), .ZN(n492) );
  XNOR2_X1 U336 ( .A(n449), .B(n448), .ZN(n451) );
  AND2_X1 U337 ( .A1(n501), .A2(n456), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n385), .B(n384), .ZN(n478) );
  XNOR2_X1 U339 ( .A(n455), .B(n454), .ZN(n566) );
  XOR2_X1 U340 ( .A(n458), .B(KEYINPUT38), .Z(n514) );
  XNOR2_X1 U341 ( .A(n495), .B(G169GAT), .ZN(n496) );
  XNOR2_X1 U342 ( .A(n482), .B(G127GAT), .ZN(n483) );
  XNOR2_X1 U343 ( .A(n459), .B(G29GAT), .ZN(n460) );
  XNOR2_X1 U344 ( .A(n497), .B(n496), .ZN(G1348GAT) );
  XNOR2_X1 U345 ( .A(n461), .B(n460), .ZN(G1328GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT6), .B(G1GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(G148GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U349 ( .A(G141GAT), .B(G85GAT), .Z(n296) );
  XNOR2_X1 U350 ( .A(G29GAT), .B(G162GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n315) );
  XOR2_X1 U353 ( .A(G57GAT), .B(KEYINPUT93), .Z(n300) );
  XNOR2_X1 U354 ( .A(KEYINPUT97), .B(KEYINPUT1), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U356 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n302) );
  XNOR2_X1 U357 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U359 ( .A(n304), .B(n303), .Z(n313) );
  XOR2_X1 U360 ( .A(KEYINPUT81), .B(G134GAT), .Z(n306) );
  XNOR2_X1 U361 ( .A(G127GAT), .B(G113GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U363 ( .A(KEYINPUT0), .B(n307), .Z(n374) );
  XNOR2_X1 U364 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n308), .B(KEYINPUT2), .ZN(n358) );
  XOR2_X1 U366 ( .A(n358), .B(KEYINPUT4), .Z(n310) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n374), .B(n311), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n530) );
  XNOR2_X1 U372 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n316), .B(KEYINPUT68), .ZN(n433) );
  XOR2_X1 U374 ( .A(G120GAT), .B(G71GAT), .Z(n369) );
  XNOR2_X1 U375 ( .A(n433), .B(n369), .ZN(n318) );
  XOR2_X1 U376 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U378 ( .A(G204GAT), .B(KEYINPUT70), .Z(n320) );
  XNOR2_X1 U379 ( .A(G92GAT), .B(G176GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U381 ( .A(G64GAT), .B(n321), .Z(n394) );
  XNOR2_X1 U382 ( .A(n322), .B(n394), .ZN(n331) );
  XOR2_X1 U383 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n324) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U386 ( .A(n325), .B(KEYINPUT31), .Z(n329) );
  XNOR2_X1 U387 ( .A(G85GAT), .B(G99GAT), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n326), .B(KEYINPUT69), .ZN(n452) );
  XNOR2_X1 U389 ( .A(G148GAT), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n327), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U391 ( .A(n452), .B(n348), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n581) );
  XOR2_X1 U394 ( .A(G1GAT), .B(G15GAT), .Z(n434) );
  XOR2_X1 U395 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n333) );
  XNOR2_X1 U396 ( .A(KEYINPUT65), .B(KEYINPUT64), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n434), .B(n334), .ZN(n338) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G22GAT), .Z(n354) );
  XNOR2_X1 U400 ( .A(n354), .B(KEYINPUT29), .ZN(n336) );
  AND2_X1 U401 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U404 ( .A(n339), .B(G197GAT), .Z(n341) );
  XOR2_X1 U405 ( .A(G8GAT), .B(G169GAT), .Z(n391) );
  XNOR2_X1 U406 ( .A(G113GAT), .B(n391), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n341), .B(n340), .ZN(n347) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G50GAT), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n342), .B(KEYINPUT8), .ZN(n343) );
  XOR2_X1 U410 ( .A(KEYINPUT7), .B(n343), .Z(n345) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(G36GAT), .ZN(n344) );
  XNOR2_X1 U412 ( .A(n345), .B(n344), .ZN(n449) );
  INV_X1 U413 ( .A(n449), .ZN(n346) );
  XOR2_X1 U414 ( .A(n347), .B(n346), .Z(n516) );
  INV_X1 U415 ( .A(n516), .ZN(n574) );
  XNOR2_X1 U416 ( .A(KEYINPUT67), .B(n574), .ZN(n541) );
  OR2_X1 U417 ( .A1(n581), .A2(n541), .ZN(n502) );
  XOR2_X1 U418 ( .A(G162GAT), .B(KEYINPUT73), .Z(n453) );
  XOR2_X1 U419 ( .A(n453), .B(n348), .Z(n350) );
  NAND2_X1 U420 ( .A1(G228GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U421 ( .A(n350), .B(n349), .ZN(n362) );
  XOR2_X1 U422 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n352) );
  XNOR2_X1 U423 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U425 ( .A(n353), .B(KEYINPUT22), .Z(n356) );
  XNOR2_X1 U426 ( .A(G50GAT), .B(n354), .ZN(n355) );
  XNOR2_X1 U427 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U428 ( .A(n357), .B(KEYINPUT90), .Z(n360) );
  XNOR2_X1 U429 ( .A(n358), .B(KEYINPUT23), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U432 ( .A(KEYINPUT91), .B(G197GAT), .Z(n364) );
  XNOR2_X1 U433 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U435 ( .A(G211GAT), .B(n365), .ZN(n386) );
  XNOR2_X1 U436 ( .A(n366), .B(n386), .ZN(n491) );
  XOR2_X1 U437 ( .A(KEYINPUT20), .B(G169GAT), .Z(n368) );
  XNOR2_X1 U438 ( .A(G190GAT), .B(G15GAT), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U440 ( .A(n370), .B(n369), .Z(n372) );
  XNOR2_X1 U441 ( .A(G43GAT), .B(G99GAT), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n374), .B(n373), .ZN(n385) );
  XOR2_X1 U444 ( .A(KEYINPUT88), .B(KEYINPUT83), .Z(n376) );
  XNOR2_X1 U445 ( .A(KEYINPUT82), .B(KEYINPUT85), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  NAND2_X1 U447 ( .A1(G227GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n291), .B(n378), .ZN(n379) );
  XOR2_X1 U449 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n381) );
  XNOR2_X1 U450 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U452 ( .A(G183GAT), .B(n382), .Z(n404) );
  XNOR2_X1 U453 ( .A(n404), .B(G176GAT), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n292), .B(n383), .ZN(n384) );
  INV_X1 U455 ( .A(n478), .ZN(n534) );
  INV_X1 U456 ( .A(n386), .ZN(n390) );
  XOR2_X1 U457 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n388) );
  XNOR2_X1 U458 ( .A(KEYINPUT99), .B(KEYINPUT101), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n390), .B(n389), .ZN(n398) );
  XOR2_X1 U461 ( .A(n391), .B(KEYINPUT75), .Z(n392) );
  XOR2_X1 U462 ( .A(G190GAT), .B(KEYINPUT74), .Z(n450) );
  XNOR2_X1 U463 ( .A(n392), .B(n290), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n396) );
  NAND2_X1 U465 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n398), .A2(n397), .ZN(n402) );
  INV_X1 U468 ( .A(n397), .ZN(n400) );
  INV_X1 U469 ( .A(n398), .ZN(n399) );
  NAND2_X1 U470 ( .A1(n400), .A2(n399), .ZN(n401) );
  NAND2_X1 U471 ( .A1(n402), .A2(n401), .ZN(n403) );
  XOR2_X1 U472 ( .A(n404), .B(n403), .Z(n486) );
  AND2_X1 U473 ( .A1(n534), .A2(n486), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n405), .B(KEYINPUT102), .ZN(n406) );
  NOR2_X1 U475 ( .A1(n491), .A2(n406), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n411) );
  BUF_X1 U477 ( .A(n486), .Z(n532) );
  XOR2_X1 U478 ( .A(KEYINPUT27), .B(n532), .Z(n415) );
  NAND2_X1 U479 ( .A1(n478), .A2(n491), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n409), .B(KEYINPUT26), .ZN(n571) );
  NOR2_X1 U481 ( .A1(n415), .A2(n571), .ZN(n410) );
  NOR2_X1 U482 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U483 ( .A(n412), .B(KEYINPUT104), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n414), .B(KEYINPUT105), .ZN(n418) );
  INV_X1 U485 ( .A(n530), .ZN(n489) );
  NOR2_X1 U486 ( .A1(n415), .A2(n489), .ZN(n477) );
  XNOR2_X1 U487 ( .A(KEYINPUT28), .B(n491), .ZN(n537) );
  NOR2_X1 U488 ( .A1(n534), .A2(n537), .ZN(n416) );
  NAND2_X1 U489 ( .A1(n477), .A2(n416), .ZN(n417) );
  NAND2_X1 U490 ( .A1(n418), .A2(n417), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n419), .B(KEYINPUT106), .ZN(n501) );
  XOR2_X1 U492 ( .A(G71GAT), .B(G78GAT), .Z(n421) );
  XNOR2_X1 U493 ( .A(G127GAT), .B(G155GAT), .ZN(n420) );
  XNOR2_X1 U494 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U495 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n423) );
  XNOR2_X1 U496 ( .A(G183GAT), .B(KEYINPUT77), .ZN(n422) );
  XNOR2_X1 U497 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U498 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U499 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n427) );
  NAND2_X1 U500 ( .A1(G231GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U501 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U502 ( .A(KEYINPUT12), .B(n428), .ZN(n429) );
  XNOR2_X1 U503 ( .A(n430), .B(n429), .ZN(n440) );
  XOR2_X1 U504 ( .A(KEYINPUT75), .B(G64GAT), .Z(n432) );
  XNOR2_X1 U505 ( .A(KEYINPUT79), .B(G8GAT), .ZN(n431) );
  XNOR2_X1 U506 ( .A(n432), .B(n431), .ZN(n438) );
  XOR2_X1 U507 ( .A(n434), .B(n433), .Z(n436) );
  XNOR2_X1 U508 ( .A(G211GAT), .B(G22GAT), .ZN(n435) );
  XNOR2_X1 U509 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U510 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U511 ( .A(n440), .B(n439), .ZN(n584) );
  XOR2_X1 U512 ( .A(G106GAT), .B(G92GAT), .Z(n442) );
  NAND2_X1 U513 ( .A1(G232GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U514 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U515 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n444) );
  XNOR2_X1 U516 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n443) );
  XNOR2_X1 U517 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U518 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U519 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U521 ( .A(KEYINPUT36), .B(n566), .ZN(n588) );
  NOR2_X1 U522 ( .A1(n584), .A2(n588), .ZN(n456) );
  OR2_X1 U523 ( .A1(n502), .A2(n529), .ZN(n458) );
  NAND2_X1 U524 ( .A1(n530), .A2(n514), .ZN(n461) );
  XOR2_X1 U525 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n459) );
  INV_X1 U526 ( .A(n584), .ZN(n564) );
  NAND2_X1 U527 ( .A1(n574), .A2(n551), .ZN(n462) );
  XOR2_X1 U528 ( .A(KEYINPUT46), .B(n462), .Z(n463) );
  NOR2_X1 U529 ( .A1(n584), .A2(n463), .ZN(n464) );
  XOR2_X1 U530 ( .A(KEYINPUT113), .B(n464), .Z(n465) );
  NAND2_X1 U531 ( .A1(n465), .A2(n566), .ZN(n467) );
  NOR2_X1 U532 ( .A1(n564), .A2(n588), .ZN(n470) );
  INV_X1 U533 ( .A(KEYINPUT45), .ZN(n468) );
  NAND2_X1 U534 ( .A1(n471), .A2(n541), .ZN(n472) );
  XNOR2_X1 U535 ( .A(KEYINPUT116), .B(n473), .ZN(n474) );
  NOR2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U537 ( .A(n476), .B(KEYINPUT48), .Z(n485) );
  NAND2_X1 U538 ( .A1(n477), .A2(n485), .ZN(n548) );
  NOR2_X1 U539 ( .A1(n478), .A2(n548), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT117), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n537), .A2(n480), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT118), .B(n481), .Z(n545) );
  NOR2_X1 U543 ( .A1(n564), .A2(n545), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1342GAT) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n488) );
  INV_X1 U547 ( .A(KEYINPUT54), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n490) );
  NAND2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n572) );
  NOR2_X1 U550 ( .A1(n491), .A2(n572), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n494), .A2(n534), .ZN(n567) );
  NOR2_X1 U553 ( .A1(n541), .A2(n567), .ZN(n497) );
  INV_X1 U554 ( .A(KEYINPUT122), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n499) );
  NAND2_X1 U556 ( .A1(n566), .A2(n584), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U558 ( .A1(n501), .A2(n500), .ZN(n517) );
  NOR2_X1 U559 ( .A1(n502), .A2(n517), .ZN(n509) );
  NAND2_X1 U560 ( .A1(n530), .A2(n509), .ZN(n503) );
  XNOR2_X1 U561 ( .A(KEYINPUT34), .B(n503), .ZN(n504) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(n504), .ZN(G1324GAT) );
  XOR2_X1 U563 ( .A(G8GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U564 ( .A1(n509), .A2(n532), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT35), .Z(n508) );
  NAND2_X1 U567 ( .A1(n509), .A2(n534), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(G1326GAT) );
  NAND2_X1 U569 ( .A1(n509), .A2(n537), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n510), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U571 ( .A1(n514), .A2(n532), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G36GAT), .B(n511), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n514), .A2(n534), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n512), .B(KEYINPUT40), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n537), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n520) );
  NAND2_X1 U579 ( .A1(n551), .A2(n516), .ZN(n528) );
  NOR2_X1 U580 ( .A1(n528), .A2(n517), .ZN(n518) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(n518), .Z(n525) );
  NAND2_X1 U582 ( .A1(n525), .A2(n530), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n521), .Z(G1332GAT) );
  XOR2_X1 U585 ( .A(G64GAT), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U586 ( .A1(n525), .A2(n532), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n534), .A2(n525), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U591 ( .A1(n525), .A2(n537), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n530), .A2(n538), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n538), .A2(n532), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n538), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT112), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n536), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(KEYINPUT44), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U604 ( .A1(n545), .A2(n541), .ZN(n542) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  INV_X1 U606 ( .A(n551), .ZN(n560) );
  NOR2_X1 U607 ( .A1(n545), .A2(n560), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n566), .A2(n545), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n548), .A2(n571), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT120), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n574), .A2(n557), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n553) );
  NAND2_X1 U618 ( .A1(n551), .A2(n557), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n584), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U624 ( .A(n566), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n567), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n564), .A2(n567), .ZN(n565) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U634 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT124), .ZN(n587) );
  NAND2_X1 U639 ( .A1(n574), .A2(n587), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n578) );
  INV_X1 U642 ( .A(KEYINPUT125), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n587), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n589) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

