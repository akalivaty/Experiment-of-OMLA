//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969;
  XOR2_X1   g000(.A(KEYINPUT75), .B(KEYINPUT6), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n206), .A2(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n211), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n205), .A2(KEYINPUT72), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n213), .A2(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT71), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n204), .B(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n212), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G113gat), .B(G120gat), .Z(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT67), .B1(new_n227), .B2(G134gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n226), .B(new_n228), .C1(new_n224), .C2(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n223), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n231), .A2(new_n227), .A3(KEYINPUT68), .A4(G134gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n221), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n221), .A2(new_n237), .A3(new_n233), .A4(new_n225), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n206), .A2(new_n207), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n213), .ZN(new_n241));
  XNOR2_X1  g040(.A(G141gat), .B(G148gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n207), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n204), .B(KEYINPUT71), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n233), .A2(new_n225), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n249), .B(new_n241), .C1(new_n244), .C2(new_n245), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n239), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n253));
  AND2_X1   g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n234), .A2(KEYINPUT73), .A3(KEYINPUT4), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n252), .A2(new_n253), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n238), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n251), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n248), .A2(new_n246), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n234), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n254), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(KEYINPUT5), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n239), .A2(new_n251), .A3(new_n256), .ZN(new_n265));
  INV_X1    g064(.A(new_n255), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT74), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n257), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G57gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n257), .A2(new_n264), .A3(new_n267), .A4(new_n272), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n203), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n202), .B1(new_n268), .B2(new_n273), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G8gat), .B(G36gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G64gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G92gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT65), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(KEYINPUT23), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n299), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n295), .A2(new_n301), .A3(KEYINPUT25), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n298), .A2(new_n303), .A3(new_n302), .A4(new_n300), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n285), .A3(new_n286), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312));
  AND2_X1   g111(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n284), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n297), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(new_n284), .C1(new_n313), .C2(new_n314), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n311), .A2(new_n312), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n324), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n322), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n318), .A2(new_n319), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(KEYINPUT66), .A3(new_n316), .A4(new_n321), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n336), .A2(new_n338), .B1(new_n305), .B2(new_n310), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n312), .A2(KEYINPUT29), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n323), .B(new_n334), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n312), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n292), .B(KEYINPUT65), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n306), .B1(new_n345), .B2(new_n287), .ZN(new_n346));
  INV_X1    g145(.A(new_n307), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n304), .A2(new_n308), .A3(new_n298), .A4(new_n300), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n346), .A2(new_n347), .B1(new_n348), .B2(new_n306), .ZN(new_n349));
  INV_X1    g148(.A(new_n322), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n334), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n282), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n311), .A2(new_n322), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n312), .A2(new_n339), .B1(new_n354), .B2(new_n340), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n281), .B(new_n342), .C1(new_n355), .C2(new_n334), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n343), .A2(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n281), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n278), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n336), .A2(new_n338), .ZN(new_n364));
  INV_X1    g163(.A(new_n248), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n311), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n311), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n248), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n339), .A2(new_n370), .A3(new_n365), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n367), .A2(new_n369), .A3(new_n373), .A4(new_n371), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT70), .ZN(new_n379));
  XNOR2_X1  g178(.A(G15gat), .B(G43gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n378), .A2(KEYINPUT70), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT33), .B1(new_n372), .B2(new_n374), .ZN(new_n385));
  INV_X1    g184(.A(new_n382), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT34), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT32), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n383), .A2(new_n387), .A3(new_n390), .A4(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT31), .B(G50gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT76), .B(G22gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n331), .B2(new_n332), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n246), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n407), .B(new_n246), .C1(new_n404), .C2(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G228gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n250), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n416), .B2(new_n334), .ZN(new_n417));
  AOI211_X1 g216(.A(KEYINPUT78), .B(new_n333), .C1(new_n250), .C2(new_n415), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n403), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n413), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n334), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT78), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(new_n414), .A3(new_n334), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(KEYINPUT79), .A3(new_n409), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n413), .B1(new_n422), .B2(new_n405), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n402), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n428), .B(new_n401), .C1(new_n420), .C2(new_n426), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n398), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n410), .A2(new_n419), .A3(new_n403), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT79), .B1(new_n425), .B2(new_n409), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n401), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(new_n429), .A3(new_n402), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n397), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n396), .A2(new_n439), .A3(KEYINPUT85), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT85), .B1(new_n396), .B2(new_n439), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n363), .B(KEYINPUT35), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n265), .A2(new_n254), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n262), .A2(new_n254), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT39), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n265), .A2(new_n446), .A3(new_n254), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(KEYINPUT40), .A3(new_n272), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n447), .A2(new_n272), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(KEYINPUT80), .A3(KEYINPUT40), .A4(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT40), .B1(new_n451), .B2(new_n445), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(new_n361), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n455), .A3(new_n274), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n457));
  AOI21_X1  g256(.A(new_n281), .B1(new_n358), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n358), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT38), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n276), .B2(new_n277), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n344), .A2(new_n351), .A3(new_n334), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n355), .A2(KEYINPUT82), .A3(new_n334), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n323), .B1(new_n339), .B2(new_n341), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n333), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT81), .B1(new_n468), .B2(new_n333), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n459), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n458), .B1(new_n473), .B2(KEYINPUT83), .ZN(new_n474));
  INV_X1    g273(.A(new_n471), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(new_n465), .A3(new_n466), .A4(new_n469), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(KEYINPUT83), .A3(KEYINPUT37), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n356), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n439), .B(new_n456), .C1(new_n462), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n439), .ZN(new_n482));
  INV_X1    g281(.A(new_n277), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n274), .A2(new_n275), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n203), .ZN(new_n485));
  INV_X1    g284(.A(new_n361), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n394), .A2(KEYINPUT36), .A3(new_n395), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT36), .B1(new_n394), .B2(new_n395), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n481), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n396), .A2(new_n439), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n362), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n442), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G85gat), .ZN(new_n499));
  AND2_X1   g298(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT8), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n498), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT98), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G99gat), .ZN(new_n509));
  INV_X1    g308(.A(G106gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT98), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n503), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n505), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT97), .B(G92gat), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n515), .A2(new_n499), .B1(KEYINPUT8), .B2(new_n503), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n513), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n498), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT99), .A4(new_n498), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G57gat), .B(G64gat), .Z(new_n523));
  OR2_X1    g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT9), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n525), .B(new_n524), .C1(new_n530), .C2(new_n527), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n522), .A2(KEYINPUT10), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT102), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n522), .A2(KEYINPUT102), .A3(KEYINPUT10), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n531), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n537), .A3(new_n521), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT101), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n518), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n532), .A2(KEYINPUT101), .A3(new_n514), .A4(new_n518), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n538), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n535), .A2(new_n536), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G230gat), .A2(G233gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n538), .A2(new_n541), .A3(new_n543), .ZN(new_n548));
  INV_X1    g347(.A(new_n546), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G120gat), .B(G148gat), .ZN(new_n552));
  INV_X1    g351(.A(G176gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(G204gat), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n547), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(G29gat), .A2(G36gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G29gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT88), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(KEYINPUT88), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(G36gat), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT15), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n570), .A4(new_n566), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n522), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT41), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(KEYINPUT100), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n520), .A2(new_n521), .B1(new_n573), .B2(new_n576), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n577), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT17), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n577), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n589), .A2(new_n591), .A3(new_n521), .A4(new_n520), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n579), .A2(new_n580), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n587), .B2(new_n592), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n563), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n594), .A3(new_n562), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT96), .B(G211gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(G1gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT16), .ZN(new_n609));
  AND2_X1   g408(.A1(G15gat), .A2(G22gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(G15gat), .A2(G22gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G15gat), .ZN(new_n613));
  INV_X1    g412(.A(G22gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G15gat), .A2(G22gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n608), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G8gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT91), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(KEYINPUT89), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n615), .A2(new_n623), .A3(new_n608), .A4(new_n616), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n612), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT90), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n625), .A2(new_n626), .A3(G8gat), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n625), .B2(G8gat), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n620), .B(new_n621), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G183gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(G8gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT90), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n626), .A3(G8gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(new_n283), .A3(new_n620), .A4(new_n621), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n630), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n630), .B2(new_n635), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n607), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n619), .B(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n632), .B2(new_n633), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n283), .B1(new_n643), .B2(new_n621), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n629), .A2(G183gat), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n636), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n607), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n635), .A3(new_n637), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G127gat), .B(G155gat), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n640), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n640), .B2(new_n649), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n606), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n639), .A3(new_n607), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n649), .A3(new_n651), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n605), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n559), .B(new_n600), .C1(new_n654), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G229gat), .A2(G233gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n589), .A2(new_n643), .A3(new_n591), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n663), .A2(KEYINPUT92), .A3(new_n577), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT92), .B1(new_n663), .B2(new_n577), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n661), .B(new_n662), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n643), .A2(new_n588), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n664), .B2(new_n665), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n661), .B(KEYINPUT93), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT13), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT92), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n643), .B2(new_n588), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n663), .A2(KEYINPUT92), .A3(new_n577), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n677), .A2(KEYINPUT18), .A3(new_n661), .A4(new_n662), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n668), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n680));
  XOR2_X1   g479(.A(G113gat), .B(G141gat), .Z(new_n681));
  XNOR2_X1  g480(.A(G169gat), .B(G197gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT12), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n679), .A2(KEYINPUT87), .A3(new_n686), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n660), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n495), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n278), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT103), .B(G1gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1324gat));
  AND2_X1   g495(.A1(new_n495), .A2(new_n692), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(G8gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT16), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n486), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G8gat), .B1(new_n693), .B2(new_n361), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT105), .Z(G1325gat));
  NAND3_X1  g505(.A1(new_n697), .A2(new_n613), .A3(new_n396), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n693), .B2(new_n490), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT106), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n439), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT107), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(new_n713), .ZN(G1327gat));
  NAND2_X1  g513(.A1(new_n654), .A2(new_n659), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n690), .A3(new_n559), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n495), .A2(new_n600), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n568), .A2(new_n569), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n485), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n495), .A2(new_n600), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n495), .A2(KEYINPUT44), .A3(new_n600), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n716), .B(KEYINPUT108), .Z(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n485), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n720), .B1(new_n728), .B2(new_n718), .ZN(G1328gat));
  INV_X1    g528(.A(G36gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n717), .A2(new_n730), .A3(new_n486), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT46), .Z(new_n732));
  AND2_X1   g531(.A1(new_n727), .A2(new_n486), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n730), .ZN(G1329gat));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n717), .A2(new_n735), .A3(new_n396), .ZN(new_n736));
  INV_X1    g535(.A(new_n490), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n725), .A2(new_n726), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(G43gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g539(.A(new_n716), .ZN(new_n741));
  NOR4_X1   g540(.A1(new_n721), .A2(G50gat), .A3(new_n439), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n726), .A3(new_n482), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(G50gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g544(.A(new_n715), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n600), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n495), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n559), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n691), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n485), .B(KEYINPUT109), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n486), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(G1333gat));
  INV_X1    g558(.A(G71gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n396), .B(KEYINPUT110), .ZN(new_n761));
  AND4_X1   g560(.A1(new_n760), .A2(new_n748), .A3(new_n750), .A4(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n495), .A2(new_n737), .A3(new_n747), .A4(new_n750), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G71gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT111), .B1(new_n762), .B2(new_n765), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(KEYINPUT50), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n751), .A2(new_n482), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n691), .A2(new_n715), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n723), .A2(new_n559), .A3(new_n724), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(new_n499), .A3(new_n278), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n495), .A2(new_n600), .A3(new_n775), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT51), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n495), .A2(new_n780), .A3(new_n600), .A4(new_n775), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n559), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n485), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n777), .B1(new_n784), .B2(new_n499), .ZN(G1336gat));
  NOR2_X1   g584(.A1(new_n361), .A2(G92gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n779), .A2(new_n559), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT113), .ZN(new_n790));
  INV_X1    g589(.A(new_n515), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n776), .B2(new_n361), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n787), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(new_n794), .A3(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n787), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n788), .B2(KEYINPUT52), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT113), .B(new_n799), .C1(new_n787), .C2(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n776), .B2(new_n490), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n396), .A2(new_n509), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n782), .B2(new_n804), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n510), .A3(new_n482), .ZN(new_n806));
  OAI21_X1  g605(.A(G106gat), .B1(new_n776), .B2(new_n439), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n806), .B(new_n807), .C1(new_n810), .C2(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1339gat));
  NAND4_X1  g613(.A1(new_n668), .A2(new_n673), .A3(new_n678), .A4(new_n686), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n670), .A2(new_n672), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n661), .B1(new_n677), .B2(new_n662), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n685), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n535), .A2(new_n549), .A3(new_n544), .A4(new_n536), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n547), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n545), .A2(new_n823), .A3(new_n546), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n555), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n820), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n547), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n555), .A4(new_n824), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n819), .A2(new_n558), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n715), .B1(new_n829), .B2(new_n600), .ZN(new_n830));
  INV_X1    g629(.A(new_n600), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n819), .A2(new_n559), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(new_n558), .A3(new_n828), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n831), .B(new_n832), .C1(new_n690), .C2(new_n833), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n830), .A2(new_n834), .B1(new_n660), .B2(new_n690), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(new_n752), .A3(new_n486), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n440), .A2(new_n441), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(G113gat), .A3(new_n690), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n835), .A2(new_n482), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n278), .A2(new_n486), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n396), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT115), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n690), .ZN(new_n845));
  INV_X1    g644(.A(G113gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n847), .B(new_n848), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n844), .B2(new_n749), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n838), .A2(G120gat), .A3(new_n749), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1341gat));
  NOR3_X1   g651(.A1(new_n844), .A2(new_n227), .A3(new_n746), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n715), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n227), .B2(new_n854), .ZN(G1342gat));
  NOR3_X1   g654(.A1(new_n838), .A2(G134gat), .A3(new_n831), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT56), .ZN(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n844), .B2(new_n831), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n830), .A2(new_n834), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n660), .A2(new_n690), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n482), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n835), .B2(new_n439), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n490), .A2(new_n842), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n691), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(G141gat), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n737), .A2(new_n439), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n836), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(G141gat), .A3(new_n690), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n866), .A2(new_n868), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n691), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(G141gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(new_n874), .ZN(G1344gat));
  AOI211_X1 g684(.A(KEYINPUT59), .B(new_n208), .C1(new_n882), .C2(new_n559), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT119), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n864), .C1(new_n835), .C2(new_n439), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n888), .A2(new_n559), .A3(new_n890), .A4(new_n868), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n208), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n559), .A2(new_n208), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n886), .A2(new_n895), .B1(new_n876), .B2(new_n896), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n876), .A2(new_n746), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n715), .ZN(new_n899));
  MUX2_X1   g698(.A(new_n898), .B(new_n899), .S(G155gat), .Z(G1346gat));
  NOR2_X1   g699(.A1(new_n876), .A2(new_n831), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n600), .ZN(new_n902));
  MUX2_X1   g701(.A(new_n901), .B(new_n902), .S(G162gat), .Z(G1347gat));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n752), .A2(new_n486), .A3(new_n761), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(KEYINPUT121), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(KEYINPUT121), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n841), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(new_n691), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n835), .A2(new_n485), .A3(new_n361), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n837), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(G169gat), .A3(new_n690), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n909), .A2(new_n912), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n908), .A2(G176gat), .A3(new_n559), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n553), .B1(new_n911), .B2(new_n749), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(G1349gat));
  OAI21_X1  g715(.A(new_n715), .B1(new_n314), .B2(new_n313), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n906), .A2(new_n715), .A3(new_n841), .A4(new_n907), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(G183gat), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT122), .B1(new_n921), .B2(KEYINPUT60), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n921), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n922), .A2(new_n923), .B1(new_n924), .B2(new_n927), .ZN(G1350gat));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n908), .A2(new_n600), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(G190gat), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT61), .B(new_n284), .C1(new_n908), .C2(new_n600), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n600), .A2(new_n284), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n931), .A2(new_n932), .B1(new_n911), .B2(new_n933), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n888), .A2(new_n890), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n888), .A2(KEYINPUT124), .A3(new_n890), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n753), .A2(new_n737), .A3(new_n361), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n691), .A4(new_n941), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n937), .A2(new_n691), .A3(new_n941), .A4(new_n938), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT125), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(G197gat), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n910), .A2(new_n875), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n946), .A2(G197gat), .A3(new_n690), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1352gat));
  NAND4_X1  g747(.A1(new_n937), .A2(new_n559), .A3(new_n941), .A4(new_n938), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n946), .A2(G204gat), .A3(new_n749), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n950), .A2(KEYINPUT126), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1353gat));
  OR3_X1    g756(.A1(new_n946), .A2(G211gat), .A3(new_n746), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n888), .A2(new_n715), .A3(new_n890), .A4(new_n941), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT127), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n959), .A2(new_n962), .ZN(new_n964));
  AND4_X1   g763(.A1(KEYINPUT63), .A2(new_n963), .A3(G211gat), .A4(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n958), .B1(new_n961), .B2(new_n965), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n939), .A2(new_n600), .A3(new_n941), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G218gat), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n831), .A2(G218gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n946), .B2(new_n969), .ZN(G1355gat));
endmodule


