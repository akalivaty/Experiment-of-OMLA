

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n565), .A2(n537), .ZN(n787) );
  XNOR2_X1 U549 ( .A(n518), .B(KEYINPUT17), .ZN(n520) );
  NAND2_X1 U550 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U551 ( .A(G2104), .B(KEYINPUT66), .ZN(n517) );
  INV_X1 U552 ( .A(KEYINPUT13), .ZN(n607) );
  XNOR2_X1 U553 ( .A(n524), .B(KEYINPUT67), .ZN(n591) );
  NOR2_X1 U554 ( .A1(n610), .A2(n609), .ZN(n612) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NOR2_X1 U556 ( .A1(n739), .A2(n515), .ZN(n513) );
  AND2_X1 U557 ( .A1(n705), .A2(n704), .ZN(n514) );
  AND2_X1 U558 ( .A1(n1020), .A2(n754), .ZN(n515) );
  AND2_X1 U559 ( .A1(G1976), .A2(G288), .ZN(n516) );
  XNOR2_X1 U560 ( .A(n616), .B(KEYINPUT65), .ZN(n631) );
  INV_X1 U561 ( .A(KEYINPUT97), .ZN(n638) );
  XNOR2_X1 U562 ( .A(n639), .B(n638), .ZN(n643) );
  INV_X1 U563 ( .A(KEYINPUT100), .ZN(n647) );
  XNOR2_X1 U564 ( .A(n647), .B(KEYINPUT29), .ZN(n648) );
  INV_X1 U565 ( .A(KEYINPUT103), .ZN(n672) );
  NAND2_X1 U566 ( .A1(n725), .A2(n600), .ZN(n625) );
  NOR2_X1 U567 ( .A1(n703), .A2(n516), .ZN(n687) );
  INV_X1 U568 ( .A(n1005), .ZN(n693) );
  OR2_X1 U569 ( .A1(n693), .A2(n692), .ZN(n694) );
  INV_X1 U570 ( .A(KEYINPUT68), .ZN(n518) );
  INV_X1 U571 ( .A(KEYINPUT70), .ZN(n531) );
  INV_X1 U572 ( .A(G651), .ZN(n537) );
  XNOR2_X1 U573 ( .A(n531), .B(KEYINPUT1), .ZN(n532) );
  NOR2_X1 U574 ( .A1(G651), .A2(n565), .ZN(n793) );
  NAND2_X1 U575 ( .A1(n612), .A2(n611), .ZN(n1017) );
  AND2_X1 U576 ( .A1(n594), .A2(n593), .ZN(n760) );
  INV_X1 U577 ( .A(G2105), .ZN(n595) );
  INV_X1 U578 ( .A(n517), .ZN(n523) );
  INV_X1 U579 ( .A(n523), .ZN(n597) );
  AND2_X1 U580 ( .A1(n595), .A2(n597), .ZN(n877) );
  NAND2_X1 U581 ( .A1(n877), .A2(G102), .ZN(n522) );
  XNOR2_X2 U582 ( .A(n520), .B(n519), .ZN(n713) );
  NAND2_X1 U583 ( .A1(G138), .A2(n713), .ZN(n521) );
  NAND2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n523), .A2(G2105), .ZN(n524) );
  NAND2_X1 U586 ( .A1(n591), .A2(G126), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT88), .ZN(n528) );
  AND2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U589 ( .A1(G114), .A2(n881), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT89), .B(n526), .Z(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n530), .A2(n529), .ZN(G164) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n565) );
  NAND2_X1 U594 ( .A1(n793), .A2(G53), .ZN(n535) );
  NOR2_X1 U595 ( .A1(G543), .A2(n537), .ZN(n533) );
  XNOR2_X2 U596 ( .A(n533), .B(n532), .ZN(n789) );
  NAND2_X1 U597 ( .A1(G65), .A2(n789), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(KEYINPUT71), .B(n536), .ZN(n541) );
  NOR2_X2 U600 ( .A1(G651), .A2(G543), .ZN(n792) );
  NAND2_X1 U601 ( .A1(G91), .A2(n792), .ZN(n539) );
  NAND2_X1 U602 ( .A1(G78), .A2(n787), .ZN(n538) );
  AND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(G299) );
  NAND2_X1 U605 ( .A1(n793), .A2(G52), .ZN(n543) );
  NAND2_X1 U606 ( .A1(G64), .A2(n789), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G90), .A2(n792), .ZN(n545) );
  NAND2_X1 U609 ( .A1(G77), .A2(n787), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(G171) );
  NAND2_X1 U613 ( .A1(n792), .A2(G89), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G76), .A2(n787), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n793), .A2(G51), .ZN(n554) );
  NAND2_X1 U619 ( .A1(G63), .A2(n789), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G88), .A2(n792), .ZN(n560) );
  NAND2_X1 U626 ( .A1(G75), .A2(n787), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n793), .A2(G50), .ZN(n562) );
  NAND2_X1 U629 ( .A1(G62), .A2(n789), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(G166) );
  XOR2_X1 U632 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U633 ( .A1(G87), .A2(n565), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n789), .A2(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n793), .A2(G49), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(G288) );
  NAND2_X1 U639 ( .A1(n792), .A2(G86), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G61), .A2(n789), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n787), .A2(G73), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n793), .A2(G48), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(G305) );
  AND2_X1 U647 ( .A1(G60), .A2(n789), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G85), .A2(n792), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G72), .A2(n787), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n793), .A2(G47), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(G290) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n725) );
  NAND2_X1 U655 ( .A1(G137), .A2(n713), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n881), .A2(G113), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n586), .A2(KEYINPUT69), .ZN(n590) );
  INV_X1 U659 ( .A(n586), .ZN(n588) );
  INV_X1 U660 ( .A(KEYINPUT69), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n594) );
  INV_X1 U663 ( .A(n591), .ZN(n592) );
  INV_X1 U664 ( .A(n592), .ZN(n880) );
  NAND2_X1 U665 ( .A1(G125), .A2(n880), .ZN(n593) );
  AND2_X1 U666 ( .A1(n595), .A2(G101), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT23), .B(n598), .Z(n759) );
  AND2_X1 U669 ( .A1(G40), .A2(n759), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n760), .A2(n599), .ZN(n726) );
  INV_X1 U671 ( .A(n726), .ZN(n600) );
  INV_X1 U672 ( .A(G1996), .ZN(n927) );
  NOR2_X1 U673 ( .A1(n625), .A2(n927), .ZN(n602) );
  XOR2_X1 U674 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n601) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(n615) );
  AND2_X1 U676 ( .A1(n625), .A2(G1341), .ZN(n613) );
  NAND2_X1 U677 ( .A1(n789), .A2(G56), .ZN(n603) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(n603), .Z(n610) );
  NAND2_X1 U679 ( .A1(G68), .A2(n787), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n792), .A2(G81), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n793), .A2(G43), .ZN(n611) );
  NOR2_X1 U685 ( .A1(n613), .A2(n1017), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n792), .A2(G92), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G66), .A2(n789), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(KEYINPUT74), .B(n619), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G79), .A2(n787), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G54), .A2(n793), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U694 ( .A(KEYINPUT15), .B(n624), .Z(n1010) );
  NAND2_X1 U695 ( .A1(n631), .A2(n1010), .ZN(n629) );
  BUF_X2 U696 ( .A(n625), .Z(n665) );
  INV_X1 U697 ( .A(n665), .ZN(n651) );
  NOR2_X1 U698 ( .A1(n651), .A2(G1348), .ZN(n627) );
  NOR2_X1 U699 ( .A1(G2067), .A2(n665), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(KEYINPUT98), .ZN(n633) );
  OR2_X1 U703 ( .A1(n1010), .A2(n631), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n641) );
  INV_X1 U705 ( .A(G2072), .ZN(n926) );
  NOR2_X1 U706 ( .A1(n665), .A2(n926), .ZN(n635) );
  XOR2_X1 U707 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n634) );
  XNOR2_X1 U708 ( .A(n635), .B(n634), .ZN(n637) );
  XNOR2_X1 U709 ( .A(G1956), .B(KEYINPUT96), .ZN(n953) );
  NAND2_X1 U710 ( .A1(n665), .A2(n953), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n639) );
  OR2_X1 U712 ( .A1(G299), .A2(n643), .ZN(n640) );
  AND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(KEYINPUT99), .ZN(n646) );
  NAND2_X1 U715 ( .A1(G299), .A2(n643), .ZN(n644) );
  XNOR2_X1 U716 ( .A(KEYINPUT28), .B(n644), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n655) );
  NOR2_X1 U719 ( .A1(n651), .A2(G1961), .ZN(n650) );
  XOR2_X1 U720 ( .A(KEYINPUT94), .B(n650), .Z(n653) );
  XNOR2_X1 U721 ( .A(KEYINPUT25), .B(G2078), .ZN(n925) );
  NAND2_X1 U722 ( .A1(n651), .A2(n925), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n659), .A2(G171), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n664) );
  NOR2_X1 U726 ( .A1(G2084), .A2(n665), .ZN(n676) );
  NAND2_X1 U727 ( .A1(G8), .A2(n665), .ZN(n703) );
  NOR2_X1 U728 ( .A1(G1966), .A2(n703), .ZN(n679) );
  NOR2_X1 U729 ( .A1(n676), .A2(n679), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G8), .A2(n656), .ZN(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT30), .B(n657), .ZN(n658) );
  NOR2_X1 U732 ( .A1(G168), .A2(n658), .ZN(n661) );
  NOR2_X1 U733 ( .A1(G171), .A2(n659), .ZN(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT31), .B(n662), .Z(n663) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n677) );
  NAND2_X1 U737 ( .A1(n677), .A2(G286), .ZN(n671) );
  NOR2_X1 U738 ( .A1(G1971), .A2(n703), .ZN(n667) );
  NOR2_X1 U739 ( .A1(G2090), .A2(n665), .ZN(n666) );
  NOR2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT102), .B(n668), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(G303), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n674), .A2(G8), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT32), .ZN(n684) );
  NAND2_X1 U747 ( .A1(G8), .A2(n676), .ZN(n682) );
  INV_X1 U748 ( .A(n677), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U750 ( .A(KEYINPUT101), .B(n680), .Z(n681) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n699) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n690) );
  NOR2_X1 U754 ( .A1(G303), .A2(G1971), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n690), .A2(n685), .ZN(n1009) );
  NAND2_X1 U756 ( .A1(n699), .A2(n1009), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT104), .ZN(n688) );
  AND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U759 ( .A1(KEYINPUT33), .A2(n689), .ZN(n695) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n1005) );
  NAND2_X1 U761 ( .A1(n690), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U762 ( .A1(n691), .A2(n703), .ZN(n692) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  INV_X1 U764 ( .A(n696), .ZN(n706) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U766 ( .A1(G8), .A2(n697), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n700), .A2(n703), .ZN(n705) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n701) );
  XOR2_X1 U770 ( .A(n701), .B(KEYINPUT24), .Z(n702) );
  OR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n706), .A2(n514), .ZN(n740) );
  NAND2_X1 U773 ( .A1(G117), .A2(n881), .ZN(n708) );
  NAND2_X1 U774 ( .A1(G129), .A2(n880), .ZN(n707) );
  NAND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n877), .A2(G105), .ZN(n709) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n712), .B(KEYINPUT92), .ZN(n715) );
  NAND2_X1 U780 ( .A1(G141), .A2(n713), .ZN(n714) );
  NAND2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n894) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n894), .ZN(n716) );
  XNOR2_X1 U783 ( .A(n716), .B(KEYINPUT93), .ZN(n724) );
  INV_X1 U784 ( .A(G1991), .ZN(n923) );
  NAND2_X1 U785 ( .A1(n877), .A2(G95), .ZN(n718) );
  NAND2_X1 U786 ( .A1(G131), .A2(n713), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G107), .A2(n881), .ZN(n720) );
  NAND2_X1 U789 ( .A1(G119), .A2(n880), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U791 ( .A1(n722), .A2(n721), .ZN(n889) );
  NOR2_X1 U792 ( .A1(n923), .A2(n889), .ZN(n723) );
  NOR2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n993) );
  NOR2_X1 U794 ( .A1(n725), .A2(n726), .ZN(n754) );
  INV_X1 U795 ( .A(n754), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n993), .A2(n727), .ZN(n745) );
  INV_X1 U797 ( .A(n745), .ZN(n738) );
  XNOR2_X1 U798 ( .A(G2067), .B(KEYINPUT37), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n877), .A2(G104), .ZN(n729) );
  NAND2_X1 U800 ( .A1(G140), .A2(n713), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n731) );
  XOR2_X1 U802 ( .A(KEYINPUT91), .B(KEYINPUT34), .Z(n730) );
  XNOR2_X1 U803 ( .A(n731), .B(n730), .ZN(n736) );
  NAND2_X1 U804 ( .A1(G116), .A2(n881), .ZN(n733) );
  NAND2_X1 U805 ( .A1(G128), .A2(n880), .ZN(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U807 ( .A(KEYINPUT35), .B(n734), .Z(n735) );
  NOR2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U809 ( .A(KEYINPUT36), .B(n737), .ZN(n897) );
  NOR2_X1 U810 ( .A1(n751), .A2(n897), .ZN(n984) );
  NAND2_X1 U811 ( .A1(n754), .A2(n984), .ZN(n749) );
  NAND2_X1 U812 ( .A1(n738), .A2(n749), .ZN(n739) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n1020) );
  NAND2_X1 U814 ( .A1(n740), .A2(n513), .ZN(n757) );
  XOR2_X1 U815 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n748) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n894), .ZN(n981) );
  AND2_X1 U817 ( .A1(n923), .A2(n889), .ZN(n741) );
  XNOR2_X1 U818 ( .A(KEYINPUT106), .B(n741), .ZN(n983) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n742) );
  XOR2_X1 U820 ( .A(n742), .B(KEYINPUT105), .Z(n743) );
  NOR2_X1 U821 ( .A1(n983), .A2(n743), .ZN(n744) );
  NOR2_X1 U822 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U823 ( .A1(n981), .A2(n746), .ZN(n747) );
  XNOR2_X1 U824 ( .A(n748), .B(n747), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n751), .A2(n897), .ZN(n992) );
  NAND2_X1 U827 ( .A1(n752), .A2(n992), .ZN(n753) );
  XNOR2_X1 U828 ( .A(KEYINPUT108), .B(n753), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U831 ( .A(n758), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U832 ( .A1(n760), .A2(n759), .ZN(G160) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U834 ( .A1(G123), .A2(n880), .ZN(n761) );
  XNOR2_X1 U835 ( .A(n761), .B(KEYINPUT18), .ZN(n769) );
  NAND2_X1 U836 ( .A1(G135), .A2(n713), .ZN(n762) );
  XNOR2_X1 U837 ( .A(n762), .B(KEYINPUT78), .ZN(n764) );
  NAND2_X1 U838 ( .A1(G111), .A2(n881), .ZN(n763) );
  NAND2_X1 U839 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U840 ( .A1(G99), .A2(n877), .ZN(n765) );
  XNOR2_X1 U841 ( .A(KEYINPUT79), .B(n765), .ZN(n766) );
  NOR2_X1 U842 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U843 ( .A1(n769), .A2(n768), .ZN(n985) );
  XNOR2_X1 U844 ( .A(G2096), .B(n985), .ZN(n770) );
  OR2_X1 U845 ( .A1(G2100), .A2(n770), .ZN(G156) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  INV_X1 U847 ( .A(G108), .ZN(G238) );
  INV_X1 U848 ( .A(G132), .ZN(G219) );
  INV_X1 U849 ( .A(G82), .ZN(G220) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U851 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U852 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n773) );
  INV_X1 U853 ( .A(G223), .ZN(n830) );
  NAND2_X1 U854 ( .A1(G567), .A2(n830), .ZN(n772) );
  XNOR2_X1 U855 ( .A(n773), .B(n772), .ZN(G234) );
  INV_X1 U856 ( .A(G860), .ZN(n780) );
  OR2_X1 U857 ( .A1(n1017), .A2(n780), .ZN(G153) );
  XNOR2_X1 U858 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NOR2_X1 U859 ( .A1(n1010), .A2(G868), .ZN(n774) );
  XNOR2_X1 U860 ( .A(n774), .B(KEYINPUT75), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(G284) );
  INV_X1 U863 ( .A(G868), .ZN(n811) );
  XNOR2_X1 U864 ( .A(KEYINPUT76), .B(n811), .ZN(n777) );
  NOR2_X1 U865 ( .A1(G286), .A2(n777), .ZN(n779) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n781), .A2(n1010), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n782), .B(KEYINPUT77), .ZN(n783) );
  XOR2_X1 U871 ( .A(KEYINPUT16), .B(n783), .Z(G148) );
  NOR2_X1 U872 ( .A1(G868), .A2(n1017), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G868), .A2(n1010), .ZN(n784) );
  NOR2_X1 U874 ( .A1(G559), .A2(n784), .ZN(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G80), .A2(n787), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n788), .B(KEYINPUT80), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G67), .A2(n789), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G93), .A2(n792), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  OR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n810) );
  NAND2_X1 U884 ( .A1(G559), .A2(n1010), .ZN(n798) );
  XNOR2_X1 U885 ( .A(n798), .B(n1017), .ZN(n808) );
  NOR2_X1 U886 ( .A1(G860), .A2(n808), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT81), .B(n799), .Z(n800) );
  XOR2_X1 U888 ( .A(n810), .B(n800), .Z(G145) );
  XNOR2_X1 U889 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n802) );
  XNOR2_X1 U890 ( .A(G288), .B(KEYINPUT19), .ZN(n801) );
  XNOR2_X1 U891 ( .A(n802), .B(n801), .ZN(n805) );
  XOR2_X1 U892 ( .A(n810), .B(G299), .Z(n803) );
  XNOR2_X1 U893 ( .A(n803), .B(G305), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n805), .B(n804), .ZN(n807) );
  XNOR2_X1 U895 ( .A(G290), .B(G166), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n807), .B(n806), .ZN(n903) );
  XNOR2_X1 U897 ( .A(n808), .B(n903), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n809), .A2(G868), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n813), .A2(n812), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2084), .A2(G2078), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n814) );
  XNOR2_X1 U903 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XOR2_X1 U905 ( .A(KEYINPUT21), .B(n817), .Z(n818) );
  NOR2_X1 U906 ( .A1(n926), .A2(n818), .ZN(n819) );
  XNOR2_X1 U907 ( .A(KEYINPUT85), .B(n819), .ZN(G158) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U909 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U910 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U911 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U912 ( .A1(G96), .A2(n822), .ZN(n835) );
  NAND2_X1 U913 ( .A1(n835), .A2(G2106), .ZN(n828) );
  NAND2_X1 U914 ( .A1(G120), .A2(G69), .ZN(n823) );
  NOR2_X1 U915 ( .A1(G237), .A2(n823), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT86), .B(n824), .Z(n825) );
  NOR2_X1 U917 ( .A1(G238), .A2(n825), .ZN(n826) );
  XNOR2_X1 U918 ( .A(KEYINPUT87), .B(n826), .ZN(n834) );
  NAND2_X1 U919 ( .A1(n834), .A2(G567), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n837) );
  NAND2_X1 U921 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n837), .A2(n829), .ZN(n833) );
  NAND2_X1 U923 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(KEYINPUT111), .ZN(G261) );
  INV_X1 U935 ( .A(G261), .ZN(G325) );
  INV_X1 U936 ( .A(n837), .ZN(G319) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(G2084), .B(G2078), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT113), .B(G1961), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n848), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1981), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1956), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U955 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT112), .B(G2474), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U958 ( .A1(n880), .A2(G124), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G136), .A2(n713), .ZN(n858) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(KEYINPUT114), .B(n860), .Z(n862) );
  NAND2_X1 U963 ( .A1(n881), .A2(G112), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G100), .A2(n877), .ZN(n863) );
  XNOR2_X1 U966 ( .A(KEYINPUT115), .B(n863), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U968 ( .A1(n877), .A2(G106), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G142), .A2(n713), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n868), .B(KEYINPUT45), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G130), .A2(n880), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n881), .A2(G118), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT116), .B(n871), .Z(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n985), .B(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(G164), .B(G160), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n893) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n891) );
  NAND2_X1 U981 ( .A1(n877), .A2(G103), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G139), .A2(n713), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n888) );
  XNOR2_X1 U984 ( .A(KEYINPUT118), .B(KEYINPUT47), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n880), .A2(G127), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n881), .A2(G115), .ZN(n882) );
  XOR2_X1 U987 ( .A(KEYINPUT117), .B(n882), .Z(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U989 ( .A(n886), .B(n885), .Z(n887) );
  NOR2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n975) );
  XNOR2_X1 U991 ( .A(n889), .B(n975), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n894), .B(G162), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n898) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U998 ( .A(n1017), .B(G286), .ZN(n901) );
  XNOR2_X1 U999 ( .A(G171), .B(n1010), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n903), .B(n902), .Z(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G397) );
  XNOR2_X1 U1003 ( .A(G2451), .B(G2427), .ZN(n914) );
  XOR2_X1 U1004 ( .A(G2430), .B(G2443), .Z(n906) );
  XNOR2_X1 U1005 ( .A(G2435), .B(G2438), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1007 ( .A(G2454), .B(KEYINPUT109), .Z(n908) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1010 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1011 ( .A(G2446), .B(KEYINPUT110), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n915), .A2(G14), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n921), .ZN(G401) );
  INV_X1 U1023 ( .A(KEYINPUT55), .ZN(n1000) );
  XNOR2_X1 U1024 ( .A(G2084), .B(G34), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(n922), .B(KEYINPUT54), .ZN(n938) );
  XNOR2_X1 U1026 ( .A(G25), .B(n923), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n924), .A2(G28), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(G27), .B(n925), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n926), .B(G33), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n927), .B(G32), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G26), .B(G2067), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(n936), .B(KEYINPUT53), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n941) );
  XOR2_X1 U1038 ( .A(G2090), .B(KEYINPUT122), .Z(n939) );
  XNOR2_X1 U1039 ( .A(G35), .B(n939), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(n1000), .B(n942), .ZN(n944) );
  INV_X1 U1042 ( .A(G29), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(G11), .A2(n945), .ZN(n974) );
  XOR2_X1 U1045 ( .A(G1961), .B(G5), .Z(n958) );
  XNOR2_X1 U1046 ( .A(KEYINPUT123), .B(G1341), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(n946), .B(G19), .ZN(n952) );
  XOR2_X1 U1048 ( .A(KEYINPUT124), .B(G4), .Z(n948) );
  XNOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT59), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(n948), .B(n947), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(G1981), .B(G6), .ZN(n949) );
  NOR2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(G20), .B(n953), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(KEYINPUT60), .B(n956), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(G21), .B(G1966), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1060 ( .A(KEYINPUT125), .B(n961), .Z(n968) );
  XOR2_X1 U1061 ( .A(G1986), .B(G24), .Z(n963) );
  XOR2_X1 U1062 ( .A(G1971), .B(G22), .Z(n962) );
  NAND2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n964) );
  NOR2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(n969), .B(KEYINPUT126), .ZN(n970) );
  XNOR2_X1 U1069 ( .A(KEYINPUT61), .B(n970), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(G16), .A2(n971), .ZN(n972) );
  XOR2_X1 U1071 ( .A(KEYINPUT127), .B(n972), .Z(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n1004) );
  XNOR2_X1 U1073 ( .A(G2072), .B(n975), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(n976), .B(KEYINPUT121), .ZN(n978) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1077 ( .A(KEYINPUT50), .B(n979), .Z(n998) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n980) );
  NOR2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1080 ( .A(KEYINPUT51), .B(n982), .Z(n991) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G2084), .B(G160), .ZN(n987) );
  XNOR2_X1 U1084 ( .A(KEYINPUT119), .B(n987), .ZN(n988) );
  NOR2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1089 ( .A(KEYINPUT120), .B(n996), .Z(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1028) );
  XOR2_X1 U1095 ( .A(KEYINPUT56), .B(G16), .Z(n1026) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G168), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT57), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(G1956), .B(G299), .Z(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(n1010), .B(G1348), .Z(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1024) );
  XNOR2_X1 U1104 ( .A(G171), .B(G1961), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(G1971), .A2(G303), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G1341), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n516), .A2(n1020), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

