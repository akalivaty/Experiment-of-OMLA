//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n463), .B1(new_n464), .B2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  AOI21_X1  g054(.A(new_n476), .B1(new_n471), .B2(new_n473), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  OR3_X1    g057(.A1(new_n481), .A2(KEYINPUT68), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n474), .B2(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT68), .B1(new_n481), .B2(new_n482), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n476), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n498));
  AOI22_X1  g073(.A1(G126), .A2(new_n480), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT4), .B1(new_n465), .B2(new_n466), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n476), .A2(G138), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n474), .B2(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT70), .A2(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n507), .B(KEYINPUT6), .C1(new_n508), .C2(KEYINPUT71), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n511), .A2(G543), .A3(new_n512), .A4(new_n513), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n508), .ZN(new_n526));
  OR3_X1    g101(.A1(new_n524), .A2(KEYINPUT73), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT73), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  AND4_X1   g104(.A1(new_n519), .A2(new_n511), .A3(new_n512), .A4(new_n513), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n523), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G168));
  XOR2_X1   g113(.A(KEYINPUT74), .B(G90), .Z(new_n539));
  NOR2_X1   g114(.A1(new_n520), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n508), .A2(new_n541), .B1(new_n523), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AND2_X1   g119(.A1(new_n530), .A2(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n508), .A2(new_n546), .B1(new_n523), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT75), .Z(G188));
  AND3_X1   g131(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n558));
  OAI21_X1  g133(.A(G65), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n564), .A3(G651), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n563), .A2(new_n565), .B1(G91), .B2(new_n530), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n514), .A2(new_n567), .A3(G53), .A4(G543), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n523), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n566), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND2_X1  g150(.A1(new_n536), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n520), .ZN(G288));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n520), .A2(new_n580), .B1(new_n508), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n536), .A2(G48), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AND2_X1   g160(.A1(new_n530), .A2(G85), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n508), .A2(new_n587), .B1(new_n523), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n520), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n519), .A2(G66), .ZN(new_n595));
  INV_X1    g170(.A(G79), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n516), .ZN(new_n597));
  AOI22_X1  g172(.A1(G54), .A2(new_n536), .B1(new_n597), .B2(G651), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT10), .B1(new_n520), .B2(new_n593), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT77), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G284));
  XOR2_X1   g177(.A(G284), .B(KEYINPUT78), .Z(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT79), .Z(G148));
  NAND2_X1  g185(.A1(new_n601), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g189(.A(new_n474), .ZN(new_n615));
  INV_X1    g190(.A(G135), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n615), .A2(KEYINPUT80), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(G111), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G2105), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n480), .B2(G123), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT80), .B1(new_n615), .B2(new_n616), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2100), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT15), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2435), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT81), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n645), .B(KEYINPUT17), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(new_n649), .B2(new_n646), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT82), .ZN(new_n651));
  INV_X1    g226(.A(new_n645), .ZN(new_n652));
  INV_X1    g227(.A(new_n646), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(new_n644), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n644), .A3(new_n646), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n671), .B(new_n672), .C1(new_n670), .C2(new_n669), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G21), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G168), .B2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(G1966), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(G29), .A2(G32), .ZN(new_n686));
  NAND3_X1  g261(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT26), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  AOI22_X1  g265(.A1(new_n474), .A2(G141), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n480), .A2(G129), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n476), .A2(G105), .A3(G2104), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT93), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n686), .B1(new_n703), .B2(G29), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n681), .A2(G20), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT97), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT23), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G299), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1956), .ZN(new_n711));
  INV_X1    g286(.A(new_n467), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n712), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(new_n476), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n474), .A2(G139), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT25), .Z(new_n717));
  AND3_X1   g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G29), .B2(G33), .ZN(new_n720));
  INV_X1    g295(.A(G2072), .ZN(new_n721));
  NOR2_X1   g296(.A1(G27), .A2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G164), .B2(G29), .ZN(new_n723));
  OAI22_X1  g298(.A1(new_n720), .A2(new_n721), .B1(G2078), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n623), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G11), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(KEYINPUT31), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(KEYINPUT31), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n706), .A2(new_n711), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n733), .A2(new_n734), .A3(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n478), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT94), .B(KEYINPUT30), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G28), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n738), .B1(G29), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n736), .A2(new_n737), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n725), .A2(G26), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n480), .A2(G128), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n474), .A2(G140), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n725), .ZN(new_n750));
  MUX2_X1   g325(.A(new_n743), .B(new_n750), .S(KEYINPUT28), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT89), .B(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n731), .A2(new_n741), .A3(new_n742), .A4(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n601), .B2(G16), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT86), .B(G1348), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G171), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G5), .B2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(G2078), .B2(new_n723), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n725), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n725), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n765), .B(new_n766), .S(KEYINPUT96), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT29), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G2090), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(G2090), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n720), .A2(new_n721), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT91), .Z(new_n772));
  NOR4_X1   g347(.A1(new_n764), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n755), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT85), .Z(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G24), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n590), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1986), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT34), .ZN(new_n781));
  NAND2_X1  g356(.A1(G288), .A2(G16), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n681), .A2(G23), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT83), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G22), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G166), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1971), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n787), .B(new_n788), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n584), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G6), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT32), .B(G1981), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n781), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n787), .A2(new_n788), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n792), .A2(new_n793), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n801), .A2(KEYINPUT34), .A3(new_n802), .A4(new_n798), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n780), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n480), .A2(G119), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n474), .A2(G131), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n476), .A2(G107), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G25), .B(new_n809), .S(G29), .Z(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT35), .B(G1991), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n810), .B(new_n811), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n777), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n777), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n814), .B(new_n817), .C1(new_n804), .C2(new_n812), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n685), .B(new_n775), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n761), .A2(new_n762), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  INV_X1    g396(.A(G19), .ZN(new_n822));
  OAI21_X1  g397(.A(KEYINPUT87), .B1(new_n822), .B2(G16), .ZN(new_n823));
  OR3_X1    g398(.A1(new_n822), .A2(KEYINPUT87), .A3(G16), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n823), .B(new_n824), .C1(new_n549), .C2(new_n681), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT88), .Z(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1341), .Z(new_n827));
  NOR3_X1   g402(.A1(new_n819), .A2(new_n821), .A3(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n813), .A2(new_n815), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n817), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n813), .A2(new_n815), .A3(new_n777), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n774), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n821), .ZN(new_n833));
  INV_X1    g408(.A(new_n827), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n685), .ZN(G150));
  XNOR2_X1  g410(.A(KEYINPUT98), .B(G93), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n520), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n838), .A2(new_n508), .B1(new_n523), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n601), .A2(G559), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT38), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n549), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT99), .B1(new_n545), .B2(new_n548), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n842), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n841), .A2(new_n848), .A3(new_n549), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n844), .B1(new_n854), .B2(G860), .ZN(G145));
  INV_X1    g430(.A(new_n718), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n700), .B2(new_n702), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n699), .A2(new_n718), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n480), .A2(G130), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n474), .A2(G142), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n476), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n626), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n748), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n505), .B(new_n809), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n748), .A3(new_n867), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n859), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n857), .A2(new_n858), .B1(new_n872), .B2(new_n873), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G162), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n875), .A2(new_n876), .A3(new_n489), .A4(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n623), .B(new_n478), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT101), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n884), .A2(new_n889), .A3(new_n885), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g467(.A1(new_n842), .A2(new_n604), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  NOR2_X1   g469(.A1(G303), .A2(G305), .ZN(new_n895));
  NOR2_X1   g470(.A1(G166), .A2(new_n584), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n590), .B(G288), .Z(new_n898));
  AND2_X1   g473(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI22_X1  g476(.A1(new_n895), .A2(new_n896), .B1(KEYINPUT103), .B2(new_n898), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n905), .B(KEYINPUT42), .C1(new_n894), .C2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(KEYINPUT42), .B2(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(new_n600), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n908), .B2(G299), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(G299), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n600), .A2(new_n566), .A3(new_n571), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n909), .B1(new_n912), .B2(KEYINPUT102), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(new_n916), .A3(new_n911), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n611), .B(new_n853), .ZN(new_n919));
  MUX2_X1   g494(.A(new_n918), .B(new_n913), .S(new_n919), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n907), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n893), .B1(new_n921), .B2(new_n604), .ZN(G295));
  OAI21_X1  g497(.A(new_n893), .B1(new_n921), .B2(new_n604), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  XNOR2_X1  g499(.A(G301), .B(G168), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n853), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n851), .A3(new_n852), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(KEYINPUT106), .A3(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n928), .A2(KEYINPUT106), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n915), .A2(new_n929), .A3(new_n917), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n928), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT107), .B1(new_n932), .B2(new_n913), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n914), .A2(new_n934), .A3(new_n928), .A4(new_n927), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n903), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n885), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n932), .B(new_n940), .C1(new_n914), .C2(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n901), .B2(new_n902), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n901), .A2(new_n944), .A3(new_n902), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n924), .B(new_n937), .C1(new_n943), .C2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n948), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n936), .A2(new_n885), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n953), .A3(KEYINPUT110), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n946), .A3(new_n947), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n924), .A4(new_n937), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n937), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n924), .B1(new_n951), .B2(new_n952), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT3), .B1(new_n472), .B2(G2104), .ZN(new_n968));
  OAI211_X1 g543(.A(G138), .B(new_n476), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n969), .A2(KEYINPUT4), .B1(new_n501), .B2(new_n500), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n494), .A2(new_n498), .ZN(new_n971));
  OAI211_X1 g546(.A(G126), .B(G2105), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n470), .A2(G40), .A3(new_n475), .A4(new_n477), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT111), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT46), .Z(new_n982));
  INV_X1    g557(.A(KEYINPUT125), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n978), .B(KEYINPUT112), .Z(new_n984));
  INV_X1    g559(.A(G2067), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n748), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n699), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n982), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n983), .B2(new_n987), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  OR2_X1    g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  INV_X1    g566(.A(new_n978), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT127), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n984), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n986), .B1(new_n699), .B2(new_n979), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n997), .A2(new_n998), .B1(new_n981), .B2(new_n703), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n809), .A2(new_n811), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n809), .A2(new_n811), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n999), .A2(new_n1001), .B1(new_n985), .B2(new_n749), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n996), .A2(new_n1003), .B1(new_n1004), .B2(new_n984), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n990), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n977), .B1(new_n974), .B2(new_n975), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(KEYINPUT116), .ZN(new_n1010));
  INV_X1    g585(.A(new_n977), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n976), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1966), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n505), .A2(new_n1017), .A3(new_n966), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1018), .A3(new_n1011), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G2084), .ZN(new_n1020));
  OAI21_X1  g595(.A(G8), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT120), .B1(G168), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(G8), .C1(new_n535), .C2(new_n537), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(KEYINPUT121), .A3(new_n1025), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n684), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1020), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1026), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1030), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1035), .B2(new_n1026), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1031), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G2078), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT53), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1032), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(G171), .B(KEYINPUT54), .Z(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1019), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1016), .A2(new_n1018), .A3(new_n1011), .A4(KEYINPUT117), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n762), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1049));
  NAND2_X1  g624(.A1(new_n1009), .A2(new_n1007), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(G2078), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1042), .A2(new_n1043), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  OR3_X1    g627(.A1(new_n1050), .A2(KEYINPUT123), .A3(new_n1041), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT123), .B1(new_n1050), .B2(new_n1041), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n1043), .ZN(new_n1056));
  INV_X1    g631(.A(G1956), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1019), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n568), .A2(new_n570), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n530), .A2(G91), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n564), .B1(new_n561), .B2(G651), .ZN(new_n1062));
  AOI211_X1 g637(.A(KEYINPUT76), .B(new_n508), .C1(new_n559), .C2(new_n560), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1059), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n566), .A2(KEYINPUT57), .A3(new_n571), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1009), .A2(new_n1007), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1058), .B2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1058), .A2(new_n1067), .A3(new_n1069), .A4(KEYINPUT119), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1073), .A2(KEYINPUT61), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1058), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1071), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n974), .A2(new_n977), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT58), .B(G1341), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1050), .A2(G1996), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n549), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(KEYINPUT59), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1084), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(KEYINPUT59), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1081), .A2(new_n549), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1078), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1348), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1047), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1079), .A2(new_n985), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n908), .A2(KEYINPUT60), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n908), .A2(KEYINPUT60), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1348), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1092), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT60), .B(new_n908), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1075), .A2(new_n1089), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1071), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1070), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n600), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1039), .B(new_n1056), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT113), .B(G1981), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n584), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n677), .B2(new_n584), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1079), .A2(new_n1022), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(KEYINPUT49), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1109), .B(new_n1110), .C1(new_n1107), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G288), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1022), .B(new_n1079), .C1(new_n1114), .C2(G1976), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1115), .B(new_n1116), .C1(G1976), .C2(new_n1114), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1113), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n527), .A2(G8), .A3(new_n528), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT55), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1050), .A2(new_n791), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(G2090), .B2(new_n1019), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G8), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1120), .A2(KEYINPUT63), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1035), .A2(G8), .A3(G168), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1026), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1021), .A2(new_n1027), .B1(new_n1132), .B2(new_n1030), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1021), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT62), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1136), .B(new_n1031), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1042), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1135), .A2(new_n1137), .A3(G171), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1104), .A2(new_n1131), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1141), .A2(new_n1127), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1127), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1119), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT63), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1126), .A2(new_n1119), .ZN(new_n1147));
  INV_X1    g722(.A(G1976), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1113), .A2(new_n1148), .A3(new_n1114), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1106), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1110), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n992), .B1(new_n991), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1003), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1152), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1157), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1006), .B1(new_n1158), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g738(.A(G319), .ZN(new_n1165));
  OR2_X1    g739(.A1(G229), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1166), .B1(new_n888), .B2(new_n890), .ZN(new_n1167));
  AOI21_X1  g741(.A(G227), .B1(new_n641), .B2(G14), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n954), .A2(new_n1167), .A3(new_n959), .A4(new_n1168), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


