//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n455), .A2(new_n448), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n469), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n464), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT70), .Z(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n470), .ZN(new_n479));
  NAND3_X1  g054(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G137), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n475), .A2(new_n483), .ZN(G160));
  AND2_X1   g059(.A1(new_n481), .A2(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n480), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  AOI211_X1 g067(.A(new_n485), .B(new_n488), .C1(new_n492), .C2(G124), .ZN(G162));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n464), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI22_X1  g071(.A1(new_n491), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n467), .B2(new_n472), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n464), .B1(new_n489), .B2(new_n490), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n501), .B2(new_n498), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(G62), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT73), .A3(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n504), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n517), .A2(KEYINPUT6), .A3(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT6), .B1(new_n517), .B2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n526), .B1(new_n504), .B2(KEYINPUT72), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(KEYINPUT6), .A3(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(new_n528), .B1(new_n512), .B2(new_n513), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n511), .B1(new_n527), .B2(new_n528), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n530), .A2(new_n535), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n505), .A2(new_n506), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n536), .A2(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n529), .A2(G90), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n529), .A2(G81), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n512), .B2(new_n513), .ZN(new_n551));
  AND2_X1   g126(.A1(G68), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n536), .A2(G43), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT75), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(new_n541), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G651), .B1(G91), .B2(new_n529), .ZN(new_n565));
  OAI211_X1 g140(.A(G53), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n536), .A2(new_n569), .A3(G53), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n568), .B1(new_n567), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n509), .A2(new_n515), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  AOI22_X1  g150(.A1(G88), .A2(new_n529), .B1(new_n536), .B2(G50), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G303));
  NAND2_X1  g152(.A1(new_n529), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n536), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(G86), .A2(new_n529), .B1(new_n536), .B2(G48), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n505), .B2(new_n506), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n583), .B1(new_n586), .B2(G651), .ZN(new_n587));
  AOI211_X1 g162(.A(KEYINPUT76), .B(new_n504), .C1(new_n584), .C2(new_n585), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n582), .B1(new_n587), .B2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n529), .A2(G85), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n512), .B2(new_n513), .ZN(new_n592));
  AND2_X1   g167(.A1(G72), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT77), .B(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n536), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT78), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n590), .A2(new_n594), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n520), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n541), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n536), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT79), .Z(new_n614));
  AOI21_X1  g189(.A(new_n603), .B1(new_n614), .B2(new_n602), .ZN(G284));
  AOI21_X1  g190(.A(new_n603), .B1(new_n614), .B2(new_n602), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  XOR2_X1   g194(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n469), .A2(new_n471), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT68), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n465), .A2(new_n466), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n630), .A2(G2104), .A3(new_n464), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT82), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n492), .A2(G123), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n639), .A2(new_n640), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n481), .A2(G135), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  OAI211_X1 g221(.A(new_n637), .B(new_n646), .C1(new_n635), .C2(new_n634), .ZN(G156));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT85), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2427), .B(G2430), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n658), .B2(new_n659), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n649), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  INV_X1    g241(.A(new_n649), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(new_n662), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT16), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n648), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n675), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(KEYINPUT87), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(KEYINPUT87), .B2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n678), .A3(new_n675), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT18), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n677), .A2(new_n681), .A3(new_n679), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2096), .B(G2100), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1971), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT20), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(new_n702), .B(new_n701), .S(new_n695), .Z(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n700), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n700), .B2(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT89), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n708), .A2(new_n710), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n693), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n715), .A2(new_n692), .A3(new_n711), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(G229));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n481), .A2(G131), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G107), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G2105), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n720), .B(new_n723), .C1(new_n492), .C2(G119), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1986), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n598), .A2(new_n600), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n727), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n728), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(G166), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G16), .B2(G22), .ZN(new_n736));
  INV_X1    g311(.A(G1971), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT32), .B(G1981), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n730), .A2(G6), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G305), .B2(G16), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n736), .A2(new_n737), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n737), .B2(new_n736), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n730), .A2(G23), .ZN(new_n745));
  INV_X1    g320(.A(G288), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n730), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT33), .B(G1976), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n742), .A2(new_n739), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n744), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT34), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n734), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(KEYINPUT36), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT36), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n757), .B(new_n758), .Z(new_n759));
  NOR2_X1   g334(.A1(G168), .A2(new_n730), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n730), .B2(G21), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT94), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n730), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n730), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n555), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G16), .B2(G19), .ZN(new_n769));
  INV_X1    g344(.A(G1341), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n767), .A2(G1961), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n764), .B(new_n771), .C1(new_n770), .C2(new_n769), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n718), .B1(KEYINPUT24), .B2(G34), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(G34), .ZN(new_n774));
  INV_X1    g349(.A(G160), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n492), .A2(G129), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT26), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n780), .B(new_n782), .C1(G141), .C2(new_n481), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n718), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n718), .B2(G32), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n778), .B1(new_n767), .B2(G1961), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n787), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n630), .A2(G127), .ZN(new_n792));
  NAND2_X1  g367(.A1(G115), .A2(G2104), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n464), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT25), .Z(new_n796));
  INV_X1    g371(.A(G139), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n501), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n718), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n718), .B2(G33), .ZN(new_n801));
  INV_X1    g376(.A(G2072), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(G28), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n718), .B1(new_n804), .B2(G28), .ZN(new_n806));
  AND2_X1   g381(.A1(KEYINPUT31), .A2(G11), .ZN(new_n807));
  NOR2_X1   g382(.A1(KEYINPUT31), .A2(G11), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n761), .B2(new_n762), .ZN(new_n810));
  NAND2_X1  g385(.A1(G164), .A2(G29), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G27), .B2(G29), .ZN(new_n812));
  INV_X1    g387(.A(G2078), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n791), .A2(new_n803), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n772), .A2(new_n790), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n788), .A2(new_n789), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n718), .A2(G35), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G162), .B2(new_n718), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT29), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2090), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n730), .A2(G4), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n614), .B2(new_n730), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT91), .B(G1348), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n645), .A2(new_n718), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT95), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(KEYINPUT95), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(new_n813), .B2(new_n812), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n830), .B1(new_n802), .B2(new_n801), .C1(new_n777), .C2(new_n776), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n730), .A2(G20), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT23), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n618), .B2(new_n730), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(G1956), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n481), .A2(G140), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT92), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n492), .A2(G128), .ZN(new_n839));
  OR2_X1    g414(.A1(G104), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT93), .Z(new_n842));
  NAND3_X1  g417(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G29), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n718), .A2(G26), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT28), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G2067), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n831), .A2(new_n836), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n816), .A2(new_n817), .A3(new_n826), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n759), .A2(new_n850), .ZN(G311));
  INV_X1    g426(.A(G311), .ZN(G150));
  NAND2_X1  g427(.A1(new_n614), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n529), .A2(G93), .ZN(new_n855));
  OAI211_X1 g430(.A(G55), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n856));
  OAI21_X1  g431(.A(G67), .B1(new_n505), .B2(new_n506), .ZN(new_n857));
  NAND2_X1  g432(.A1(G80), .A2(G543), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G651), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n855), .B(new_n856), .C1(new_n860), .C2(KEYINPUT98), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(KEYINPUT98), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n856), .B1(new_n520), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g441(.A(KEYINPUT98), .B(new_n504), .C1(new_n857), .C2(new_n858), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(KEYINPUT98), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n555), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n854), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n861), .A2(new_n862), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(new_n874), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(G145));
  NOR2_X1   g455(.A1(new_n495), .A2(new_n496), .ZN(new_n881));
  INV_X1    g456(.A(new_n491), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(G126), .ZN(new_n883));
  INV_X1    g458(.A(new_n499), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n628), .B2(new_n629), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT4), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n481), .B2(G138), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n843), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n843), .A2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n492), .A2(G130), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  INV_X1    g470(.A(G118), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(G2105), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n481), .B2(G142), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n894), .B(new_n898), .C1(new_n889), .C2(new_n890), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n632), .A2(new_n724), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n632), .A2(new_n724), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n784), .A2(new_n799), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n779), .A2(new_n783), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n907), .A2(new_n794), .A3(new_n798), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n903), .B(new_n904), .C1(new_n908), .C2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n645), .B(G160), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(G162), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n900), .A2(new_n910), .A3(new_n901), .A4(new_n911), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n913), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(KEYINPUT100), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n922));
  AOI211_X1 g497(.A(new_n922), .B(new_n915), .C1(new_n913), .C2(new_n916), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g500(.A(new_n871), .B(KEYINPUT101), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(new_n623), .ZN(new_n927));
  INV_X1    g502(.A(new_n613), .ZN(new_n928));
  NAND2_X1  g503(.A1(G299), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n613), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(G299), .A2(new_n928), .A3(KEYINPUT102), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n935), .A3(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n927), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n933), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n937), .B(KEYINPUT103), .C1(new_n927), .C2(new_n938), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n927), .A2(KEYINPUT103), .A3(new_n938), .ZN(new_n940));
  NAND2_X1  g515(.A1(G305), .A2(new_n746), .ZN(new_n941));
  OAI211_X1 g516(.A(G288), .B(new_n582), .C1(new_n587), .C2(new_n588), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n516), .B2(new_n524), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n575), .A2(KEYINPUT104), .A3(new_n576), .ZN(new_n947));
  NAND3_X1  g522(.A1(G290), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G290), .B1(new_n946), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n729), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n943), .A3(new_n948), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT42), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n953), .A2(new_n943), .A3(new_n948), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n943), .B1(new_n953), .B2(new_n948), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(KEYINPUT105), .A3(new_n954), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n961), .B2(KEYINPUT42), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n939), .A2(new_n940), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n939), .B2(new_n940), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(G868), .B2(new_n877), .ZN(G295));
  OAI21_X1  g542(.A(new_n966), .B1(G868), .B2(new_n877), .ZN(G331));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  AOI21_X1  g544(.A(G286), .B1(G171), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n863), .B1(new_n861), .B2(new_n862), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n868), .A2(new_n555), .A3(new_n869), .ZN(new_n973));
  NAND2_X1  g548(.A1(G301), .A2(KEYINPUT106), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n974), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n864), .B2(new_n870), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n970), .A3(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n934), .A2(new_n936), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n938), .A2(new_n977), .A3(new_n981), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n960), .B(new_n959), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n934), .A2(new_n936), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n938), .A2(new_n977), .A3(new_n981), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n961), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n989), .A3(new_n918), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n975), .A2(new_n976), .A3(new_n971), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT41), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n938), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n929), .A2(new_n931), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n986), .A2(KEYINPUT41), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n961), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n984), .A3(new_n1000), .A4(new_n918), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n991), .A2(new_n992), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n984), .A3(new_n918), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n987), .A2(new_n988), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n959), .A2(new_n960), .ZN(new_n1009));
  AOI21_X1  g584(.A(G37), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n1000), .A3(new_n989), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT108), .B(new_n1002), .C1(new_n1012), .C2(KEYINPUT44), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1000), .B1(new_n1010), .B2(new_n999), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1015), .B2(KEYINPUT107), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1007), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1002), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1013), .A2(new_n1020), .ZN(G397));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(G164), .B2(G1384), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n477), .A2(new_n482), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n630), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1024), .B(G40), .C1(new_n1025), .C2(new_n464), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n843), .B(G2067), .Z(new_n1029));
  INV_X1    g604(.A(G1996), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n907), .B(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT109), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n724), .A2(new_n726), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n724), .A2(new_n726), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1027), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G290), .B(G1986), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1027), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G40), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n475), .A2(new_n1040), .A3(new_n483), .ZN(new_n1041));
  INV_X1    g616(.A(G1384), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1023), .A3(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT56), .B(G2072), .Z(new_n1045));
  OR2_X1    g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n888), .A2(new_n1048), .A3(new_n1042), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT116), .B(G1956), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n567), .A2(new_n570), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n565), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT117), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n618), .A2(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(KEYINPUT117), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(G160), .A2(G40), .A3(new_n1042), .A4(new_n888), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G2067), .ZN(new_n1065));
  INV_X1    g640(.A(G1348), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1050), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n613), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1046), .A2(new_n1061), .A3(new_n1052), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1063), .A2(KEYINPUT61), .A3(new_n1069), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n613), .B1(new_n1067), .B2(KEYINPUT60), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(KEYINPUT60), .B2(new_n1067), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT58), .B(G1341), .Z(new_n1078));
  NAND2_X1  g653(.A1(new_n1064), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(G1996), .B2(new_n1044), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n555), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT59), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1067), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1070), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1041), .A2(new_n1023), .A3(new_n1043), .A4(new_n813), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1041), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(G1961), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1024), .B(KEYINPUT121), .ZN(new_n1092));
  NOR4_X1   g667(.A1(new_n475), .A2(new_n1088), .A3(new_n1040), .A4(G2078), .ZN(new_n1093));
  AND4_X1   g668(.A1(new_n1023), .A2(new_n1092), .A3(new_n1043), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1087), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n1096), .A2(KEYINPUT123), .A3(G301), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT123), .B1(new_n1096), .B2(G301), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1086), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1088), .B1(new_n1100), .B2(KEYINPUT119), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(KEYINPUT119), .B2(new_n1100), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1102), .A3(G301), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1097), .A2(new_n1098), .A3(KEYINPUT54), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G86), .ZN(new_n1105));
  INV_X1    g680(.A(G48), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n520), .A2(new_n1105), .B1(new_n522), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n504), .B1(new_n584), .B2(new_n585), .ZN(new_n1108));
  OAI21_X1  g683(.A(G1981), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(G305), .B2(G1981), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT49), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1109), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1064), .A3(G8), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n746), .A2(G1976), .ZN(new_n1115));
  INV_X1    g690(.A(G1976), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(G288), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1064), .A2(G8), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1064), .A2(KEYINPUT112), .A3(G8), .A4(new_n1115), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n888), .A2(new_n1042), .ZN(new_n1122));
  OAI211_X1 g697(.A(G8), .B(new_n1115), .C1(new_n1026), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(G8), .B1(new_n516), .B2(new_n524), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT55), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT111), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT110), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT111), .ZN(new_n1131));
  NAND4_X1  g706(.A1(G303), .A2(new_n1131), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1130), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G2090), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1090), .A2(new_n1137), .B1(new_n1044), .B2(new_n737), .ZN(new_n1138));
  INV_X1    g713(.A(G8), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1133), .B(new_n1136), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1044), .A2(new_n737), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1041), .A2(new_n1047), .A3(new_n1049), .A4(new_n1137), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1136), .A2(new_n1133), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1126), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT122), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1126), .A2(new_n1140), .A3(new_n1148), .A4(new_n1145), .ZN(new_n1149));
  NAND2_X1  g724(.A1(G286), .A2(G8), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1090), .A2(new_n777), .B1(new_n1044), .B2(new_n762), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT51), .B(new_n1150), .C1(new_n1151), .C2(new_n1139), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1044), .A2(new_n762), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1041), .A2(new_n1047), .A3(new_n1049), .A4(new_n777), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1153), .B(G8), .C1(new_n1156), .C2(G286), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1150), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT118), .B(new_n1150), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1152), .B(new_n1157), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1147), .A2(new_n1149), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1096), .A2(G301), .ZN(new_n1165));
  AOI21_X1  g740(.A(G301), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1085), .A2(new_n1104), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1147), .A2(new_n1166), .A3(new_n1149), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1170), .A2(KEYINPUT62), .A3(new_n1152), .A4(new_n1157), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1169), .A2(KEYINPUT124), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT124), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1168), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1125), .A2(new_n1120), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1151), .A2(new_n1139), .A3(G286), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(KEYINPUT63), .A3(new_n1140), .A4(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1126), .A2(new_n1140), .A3(new_n1182), .A4(new_n1145), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT63), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1183), .A2(new_n1186), .A3(KEYINPUT114), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1114), .A2(new_n1116), .A3(new_n746), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(G1981), .B2(G305), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT113), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1064), .A2(G8), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1192), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1191), .A2(new_n1193), .B1(new_n1126), .B2(new_n1178), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT114), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1184), .A2(new_n1195), .A3(new_n1185), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT115), .B1(new_n1187), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1183), .A2(new_n1186), .A3(KEYINPUT114), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT115), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1199), .A2(new_n1200), .A3(new_n1196), .A4(new_n1194), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1039), .B1(new_n1177), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1028), .B1(new_n1029), .B2(new_n784), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT46), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1208));
  XOR2_X1   g783(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1209));
  XNOR2_X1  g784(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1211));
  OR2_X1    g786(.A1(new_n843), .A2(G2067), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1028), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1027), .A2(new_n728), .A3(new_n729), .ZN(new_n1214));
  XOR2_X1   g789(.A(new_n1214), .B(KEYINPUT48), .Z(new_n1215));
  NOR2_X1   g790(.A1(new_n1037), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1210), .A2(new_n1213), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1203), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g793(.A1(G227), .A2(new_n462), .ZN(new_n1220));
  NOR2_X1   g794(.A1(G229), .A2(new_n1220), .ZN(new_n1221));
  AND3_X1   g795(.A1(new_n924), .A2(new_n673), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n991), .A2(new_n1001), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  NAND2_X1  g801(.A1(new_n1222), .A2(new_n1224), .ZN(G225));
endmodule


