//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(G20), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n224), .A2(new_n225), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n215), .B(new_n221), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n219), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n209), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G77), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n255), .A2(new_n257), .B1(G77), .B2(new_n250), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT8), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT8), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(KEYINPUT68), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT15), .B(G87), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n268), .A2(new_n271), .B1(new_n210), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n253), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT69), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n275), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n258), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n283), .A2(G232), .B1(G107), .B2(new_n282), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G238), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT66), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT66), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n209), .C1(G41), .C2(G45), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n291), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n298), .A2(G244), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n290), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n278), .B1(new_n279), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT70), .B(G200), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n290), .B2(new_n302), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n258), .ZN(new_n308));
  INV_X1    g0108(.A(new_n277), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n274), .A2(new_n275), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n290), .A2(new_n312), .A3(new_n302), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n303), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n271), .B2(new_n272), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n320), .A2(new_n253), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT11), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n251), .A2(new_n318), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(KEYINPUT11), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n254), .A2(G68), .A3(new_n256), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n322), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n301), .A2(new_n294), .A3(G274), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n292), .A2(G238), .A3(new_n294), .A4(new_n296), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n269), .A2(new_n205), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G226), .A2(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G232), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(G1698), .ZN(new_n333));
  OR2_X1    g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n330), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n328), .B(new_n329), .C1(new_n337), .C2(new_n294), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n332), .A2(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G226), .B2(G1698), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n343), .A2(new_n282), .B1(new_n269), .B2(new_n205), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n289), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n345), .A2(new_n328), .A3(new_n329), .A4(new_n339), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n327), .B1(new_n347), .B2(G200), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n338), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT72), .B1(new_n338), .B2(KEYINPUT13), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n338), .A2(new_n340), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G190), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n317), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n283), .A2(G222), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT67), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n356), .B(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n286), .A2(G223), .B1(G77), .B2(new_n282), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n294), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G226), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n328), .B1(new_n297), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n312), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n254), .A2(G50), .A3(new_n256), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n263), .A2(new_n270), .B1(G150), .B2(new_n264), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n203), .A2(G20), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n253), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n365), .B1(G50), .B2(new_n250), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n314), .B1(new_n360), .B2(new_n362), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n363), .A2(G190), .ZN(new_n374));
  INV_X1    g0174(.A(new_n305), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n360), .B2(new_n362), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT9), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n370), .A2(new_n377), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n374), .A2(new_n376), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n379), .A2(new_n378), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT10), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n374), .A4(new_n376), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n373), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n347), .A2(G169), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n350), .A2(new_n351), .ZN(new_n388));
  INV_X1    g0188(.A(new_n349), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G179), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n314), .B1(new_n341), .B2(new_n346), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT73), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n387), .B(new_n390), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n327), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n263), .A2(new_n256), .ZN(new_n398));
  INV_X1    g0198(.A(new_n263), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n398), .A2(new_n254), .B1(new_n251), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n282), .B2(new_n210), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NOR4_X1   g0203(.A1(new_n280), .A2(new_n281), .A3(new_n403), .A4(G20), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n259), .A2(new_n318), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n201), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n264), .A2(G159), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n369), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n401), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n292), .A2(G232), .A3(new_n294), .A4(new_n296), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n328), .ZN(new_n417));
  OR2_X1    g0217(.A1(G223), .A2(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n361), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n280), .C2(new_n281), .ZN(new_n420));
  INV_X1    g0220(.A(G87), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n269), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n294), .B1(new_n424), .B2(KEYINPUT74), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  AOI211_X1 g0227(.A(G190), .B(new_n417), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(KEYINPUT74), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n289), .A3(new_n427), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n416), .A2(new_n328), .ZN(new_n431));
  AOI21_X1  g0231(.A(G200), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n415), .B(KEYINPUT17), .C1(new_n428), .C2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n334), .A2(new_n210), .A3(new_n335), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n403), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n318), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n412), .B1(new_n437), .B2(new_n409), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n414), .A3(new_n253), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n400), .C1(new_n428), .C2(new_n432), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n433), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(G223), .A2(G1698), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n361), .B2(G1698), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n422), .B1(new_n445), .B2(new_n336), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n289), .B1(new_n446), .B2(new_n426), .ZN(new_n447));
  INV_X1    g0247(.A(new_n427), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n312), .B(new_n431), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n417), .B1(new_n425), .B2(new_n427), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G169), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT18), .B1(new_n415), .B2(new_n451), .ZN(new_n452));
  AOI211_X1 g0252(.A(G179), .B(new_n417), .C1(new_n425), .C2(new_n427), .ZN(new_n453));
  AOI21_X1  g0253(.A(G169), .B1(new_n430), .B2(new_n431), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n439), .A2(new_n400), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n443), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n355), .A2(new_n385), .A3(new_n397), .A4(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(G244), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT77), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT77), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n336), .A2(new_n464), .A3(G244), .A4(new_n285), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G250), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT4), .A2(G244), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n285), .B(new_n472), .C1(new_n280), .C2(new_n281), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n336), .A2(KEYINPUT78), .A3(new_n285), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n467), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n289), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n289), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G257), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n209), .A2(G45), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n482), .B2(new_n483), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n300), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n479), .A2(G190), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT75), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n494), .B1(new_n498), .B2(new_n206), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n207), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT76), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT75), .B(G97), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT6), .B1(new_n504), .B2(G107), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n501), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n507), .A3(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n435), .A2(new_n436), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(G107), .B1(G77), .B2(new_n264), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n369), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n251), .A2(new_n205), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n209), .A2(G33), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n250), .A2(new_n513), .A3(new_n219), .A4(new_n252), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(new_n205), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n490), .B1(new_n478), .B2(new_n289), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(G190), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n294), .B1(new_n520), .B2(new_n467), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n521), .B2(new_n490), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n493), .A2(new_n516), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n479), .A2(new_n312), .A3(new_n491), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n314), .B1(new_n521), .B2(new_n490), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n511), .C2(new_n515), .ZN(new_n526));
  INV_X1    g0326(.A(new_n268), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n250), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n514), .A2(new_n421), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G87), .A2(G107), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n504), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n210), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n336), .A2(new_n210), .A3(G68), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n504), .B2(new_n271), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  AOI211_X1 g0338(.A(new_n528), .B(new_n529), .C1(new_n538), .C2(new_n253), .ZN(new_n539));
  OAI211_X1 g0339(.A(G244), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n540));
  OAI211_X1 g0340(.A(G238), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n289), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n294), .A2(G250), .A3(new_n487), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n294), .A2(G274), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n487), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n375), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n547), .B1(new_n543), .B2(new_n289), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n539), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n538), .A2(new_n253), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n514), .A2(new_n268), .ZN(new_n555));
  INV_X1    g0355(.A(new_n528), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n549), .A2(new_n314), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n312), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n523), .A2(new_n526), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g0363(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n206), .A2(G20), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT82), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n568), .B(new_n565), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n565), .A2(KEYINPUT23), .B1(G20), .B2(new_n542), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n567), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n210), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n336), .A2(new_n579), .A3(new_n210), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n576), .B1(new_n575), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n253), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT25), .B1(new_n251), .B2(new_n206), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n206), .B2(new_n514), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n591));
  OAI211_X1 g0391(.A(G250), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n289), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n485), .A2(G264), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n489), .ZN(new_n597));
  INV_X1    g0397(.A(G200), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n289), .A2(new_n594), .B1(new_n485), .B2(G264), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n279), .A3(new_n489), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n585), .A2(new_n590), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT83), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n597), .A2(new_n604), .A3(new_n312), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n597), .A2(G169), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT83), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(G179), .A3(new_n489), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n573), .B1(new_n610), .B2(KEYINPUT82), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n581), .A2(new_n611), .A3(new_n572), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT24), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n582), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n589), .B1(new_n614), .B2(new_n253), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n603), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n485), .A2(G270), .B1(new_n300), .B2(new_n488), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n619));
  INV_X1    g0419(.A(G303), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n336), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n289), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n314), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  MUX2_X1   g0423(.A(new_n250), .B(new_n514), .S(G116), .Z(new_n624));
  OAI211_X1 g0424(.A(new_n210), .B(new_n469), .C1(new_n504), .C2(G33), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n252), .A2(new_n219), .B1(G20), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT20), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(G33), .B1(new_n495), .B2(new_n497), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n469), .A2(new_n210), .ZN(new_n630));
  OAI211_X1 g0430(.A(KEYINPUT20), .B(new_n627), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n624), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n623), .A2(new_n633), .A3(KEYINPUT21), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT80), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n623), .A2(new_n633), .A3(KEYINPUT80), .A4(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n623), .A2(new_n633), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n617), .A2(new_n622), .A3(G179), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n639), .A2(new_n640), .B1(new_n642), .B2(new_n633), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n617), .A2(new_n622), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n633), .B1(G200), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n279), .B2(new_n644), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n638), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n461), .A2(new_n563), .A3(new_n616), .A4(new_n647), .ZN(G372));
  NOR3_X1   g0448(.A1(new_n415), .A2(KEYINPUT18), .A3(new_n451), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n457), .B1(new_n455), .B2(new_n456), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n440), .B(KEYINPUT17), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n316), .B1(new_n353), .B2(new_n348), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n327), .B2(new_n396), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI211_X1 g0456(.A(KEYINPUT86), .B(new_n653), .C1(new_n327), .C2(new_n396), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n381), .A2(new_n384), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n373), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT85), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n561), .B1(new_n526), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n516), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(KEYINPUT85), .A3(new_n524), .A4(new_n525), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT26), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n526), .A2(new_n561), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n560), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT84), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n638), .A2(new_n643), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n609), .A2(new_n615), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n603), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n669), .B1(new_n672), .B2(new_n563), .ZN(new_n673));
  INV_X1    g0473(.A(new_n603), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n638), .A2(new_n643), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n609), .A2(new_n615), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n563), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(KEYINPUT84), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n668), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n660), .B1(new_n461), .B2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n633), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n675), .A2(new_n646), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n675), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n616), .ZN(new_n692));
  INV_X1    g0492(.A(new_n687), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n615), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n676), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n675), .A2(new_n616), .A3(new_n687), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n671), .B2(new_n693), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n213), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n209), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n531), .A2(G116), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n702), .A2(new_n703), .B1(new_n218), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT87), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n662), .A2(new_n664), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .ZN(new_n709));
  INV_X1    g0509(.A(new_n560), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n526), .A2(new_n561), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n666), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n709), .B(new_n712), .C1(new_n563), .C2(new_n672), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n707), .B1(new_n713), .B2(new_n693), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n679), .A2(new_n673), .ZN(new_n715));
  INV_X1    g0515(.A(new_n668), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n687), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n714), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n544), .A2(new_n595), .A3(new_n548), .A4(new_n596), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n641), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n517), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n644), .A2(new_n597), .A3(new_n312), .A4(new_n549), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n517), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n517), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT31), .B1(new_n729), .B2(new_n687), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n647), .A2(new_n616), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n678), .A2(new_n733), .A3(new_n693), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n719), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n706), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G20), .A3(new_n279), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n336), .B1(new_n742), .B2(G329), .ZN(new_n743));
  INV_X1    g0543(.A(G326), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n210), .A2(new_n312), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n279), .A3(G200), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  INV_X1    g0549(.A(G294), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n210), .B1(new_n740), .B2(G190), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n210), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n375), .A2(new_n279), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT90), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n745), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT90), .B1(new_n210), .B2(new_n312), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n758), .A2(G190), .A3(new_n598), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G283), .A2(new_n756), .B1(new_n761), .B2(G322), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n758), .A2(new_n279), .A3(new_n598), .A4(new_n759), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n753), .B(new_n762), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n375), .A2(G190), .A3(new_n754), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT94), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n769), .B1(G303), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G77), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n751), .B(KEYINPUT95), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n205), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n336), .B1(new_n748), .B2(new_n318), .C1(new_n202), .C2(new_n746), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n760), .A2(new_n259), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n755), .A2(new_n206), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n742), .A2(G159), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT93), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n775), .A2(G87), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n781), .A2(new_n788), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT96), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n776), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n219), .B1(G20), .B2(new_n314), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n210), .A2(G13), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT88), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G45), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n702), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n700), .A2(new_n282), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G355), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G116), .B2(new_n213), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n700), .A2(new_n336), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n480), .B2(new_n218), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n245), .A2(new_n480), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n797), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n803), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT89), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n798), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  INV_X1    g0620(.A(new_n814), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n690), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n691), .A2(new_n803), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(G330), .B2(new_n690), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NOR2_X1   g0626(.A1(new_n797), .A2(new_n812), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n803), .B1(G77), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n748), .ZN(new_n830));
  INV_X1    g0630(.A(new_n746), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n830), .A2(G150), .B1(new_n831), .B2(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G143), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n760), .C1(new_n779), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n755), .A2(new_n318), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n336), .B1(new_n741), .B2(new_n838), .C1(new_n259), .C2(new_n751), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n837), .B(new_n839), .C1(new_n775), .C2(G50), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n336), .B1(new_n742), .B2(G311), .ZN(new_n842));
  INV_X1    g0642(.A(G283), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n748), .C1(new_n620), .C2(new_n746), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n755), .A2(new_n421), .B1(new_n760), .B2(new_n750), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n784), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n206), .B2(new_n774), .C1(new_n779), .C2(new_n626), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n829), .B1(new_n848), .B2(new_n797), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n304), .A2(new_n306), .B1(new_n278), .B2(new_n693), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n316), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n316), .A2(new_n687), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n849), .A2(KEYINPUT98), .B1(new_n812), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(KEYINPUT98), .B2(new_n849), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n307), .A2(new_n316), .A3(new_n693), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n680), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n852), .B1(new_n850), .B2(new_n316), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n737), .C1(new_n717), .C2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(KEYINPUT99), .A3(new_n802), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n858), .B1(new_n717), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n736), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT99), .B1(new_n860), .B2(new_n802), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(G384));
  NOR3_X1   g0666(.A1(new_n219), .A2(new_n210), .A3(new_n626), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n503), .A2(new_n507), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT35), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT36), .ZN(new_n872));
  OR3_X1    g0672(.A1(new_n217), .A2(new_n272), .A3(new_n406), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n202), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n209), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n685), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n456), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n652), .B2(new_n651), .ZN(new_n879));
  NOR2_X1   g0679(.A1(KEYINPUT101), .A2(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n440), .ZN(new_n881));
  NAND2_X1  g0681(.A1(KEYINPUT101), .A2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n415), .B2(new_n451), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n455), .A2(new_n456), .B1(KEYINPUT101), .B2(KEYINPUT37), .ZN(new_n885));
  INV_X1    g0685(.A(new_n880), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(new_n440), .A3(new_n878), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT38), .B1(new_n879), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n884), .A2(new_n887), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n456), .B(new_n877), .C1(new_n443), .C2(new_n459), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT39), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT102), .A4(KEYINPUT39), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n890), .B(new_n891), .C1(KEYINPUT103), .C2(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n884), .A2(new_n887), .A3(KEYINPUT103), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n892), .B(new_n899), .C1(new_n879), .C2(new_n888), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n896), .B(new_n897), .C1(KEYINPUT39), .C2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n327), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n347), .A2(new_n393), .A3(G169), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT73), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n352), .A2(G179), .B1(new_n386), .B2(KEYINPUT14), .ZN(new_n908));
  AOI211_X1 g0708(.A(KEYINPUT100), .B(new_n903), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT100), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n396), .B2(new_n327), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n687), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n853), .B1(new_n680), .B2(new_n857), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n397), .A2(KEYINPUT100), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n396), .A2(new_n910), .A3(new_n327), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n327), .A2(new_n687), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n354), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n919), .B1(new_n354), .B2(new_n396), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n889), .A2(new_n893), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n924), .A2(new_n925), .B1(new_n651), .B2(new_n877), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n461), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n719), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n660), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n927), .B(new_n930), .Z(new_n931));
  INV_X1    g0731(.A(G330), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n854), .B1(new_n732), .B2(new_n734), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n901), .A2(new_n923), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n922), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n912), .B2(new_n920), .ZN(new_n936));
  NOR4_X1   g0736(.A1(new_n563), .A2(new_n647), .A3(new_n616), .A4(new_n687), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT31), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n517), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT30), .B1(new_n721), .B2(new_n517), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n939), .A2(new_n940), .A3(new_n726), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n938), .B1(new_n941), .B2(new_n693), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n859), .B1(new_n937), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n936), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n889), .A2(new_n893), .A3(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n934), .A2(KEYINPUT40), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n461), .B1(new_n734), .B2(new_n732), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n932), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n931), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n209), .B2(new_n800), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n931), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n876), .B1(new_n955), .B2(new_n956), .ZN(G367));
  NAND2_X1  g0757(.A1(new_n807), .A2(new_n241), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n816), .B1(new_n700), .B2(new_n527), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n802), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n539), .A2(new_n693), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n710), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n561), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT107), .B1(new_n774), .B2(new_n626), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n780), .A2(G283), .B1(KEYINPUT46), .B2(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n755), .A2(new_n504), .B1(new_n760), .B2(new_n620), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n336), .B1(new_n742), .B2(G317), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n206), .B2(new_n751), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n748), .A2(new_n750), .B1(new_n746), .B2(new_n768), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n965), .B(new_n970), .C1(KEYINPUT46), .C2(new_n964), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT108), .Z(new_n972));
  INV_X1    g0772(.A(G150), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n755), .A2(new_n272), .B1(new_n760), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n282), .B1(new_n742), .B2(G137), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n833), .B2(new_n746), .C1(new_n834), .C2(new_n748), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(G68), .C2(new_n782), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n259), .B2(new_n774), .C1(new_n779), .C2(new_n202), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(KEYINPUT47), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n797), .B1(new_n980), .B2(KEYINPUT47), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n960), .B1(new_n821), .B2(new_n963), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n696), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n523), .B(new_n526), .C1(new_n516), .C2(new_n693), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n526), .B2(new_n693), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n697), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT42), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n985), .A2(new_n676), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n687), .B1(new_n991), .B2(new_n526), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n988), .A2(new_n989), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n993), .A2(new_n994), .B1(KEYINPUT43), .B2(new_n963), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT104), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n996), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n987), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n987), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n801), .A2(G1), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n698), .A2(new_n986), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n698), .A2(new_n1012), .A3(new_n986), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n698), .B2(new_n986), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT105), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT106), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT106), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT105), .B1(new_n984), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1018), .A2(new_n984), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n697), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n675), .A2(new_n687), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n695), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(new_n691), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n738), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n738), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n701), .B(KEYINPUT41), .Z(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1008), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n983), .B1(new_n1007), .B2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n1008), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1025), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n695), .A2(new_n821), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n808), .B1(new_n238), .B2(G45), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n703), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n804), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n399), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n480), .B1(new_n318), .B2(new_n272), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n263), .B2(new_n202), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1038), .A2(new_n1043), .B1(G107), .B2(new_n213), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n802), .B(new_n1035), .C1(new_n815), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n782), .A2(new_n527), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n775), .A2(G77), .B1(G68), .B2(new_n766), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n336), .B1(new_n973), .B2(new_n741), .C1(new_n399), .C2(new_n748), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G159), .B2(new_n831), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G97), .A2(new_n756), .B1(new_n761), .B2(G50), .ZN(new_n1050));
  AND4_X1   g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n774), .A2(new_n750), .B1(new_n843), .B2(new_n751), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n780), .A2(G303), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT110), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT109), .B(G322), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n768), .A2(new_n748), .B1(new_n746), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n761), .B2(G317), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n779), .B2(new_n620), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT110), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OAI211_X1 g0863(.A(KEYINPUT111), .B(new_n1053), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT111), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n1052), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1064), .A2(new_n1067), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n282), .B1(new_n744), .B2(new_n741), .C1(new_n755), .C2(new_n626), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1068), .B2(KEYINPUT49), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1051), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n797), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1045), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(KEYINPUT112), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n1045), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1034), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1025), .B1(new_n719), .B2(new_n737), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1027), .A2(new_n1079), .A3(new_n701), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(G393));
  XNOR2_X1  g0881(.A(new_n1016), .B(new_n984), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1027), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1083), .B(new_n701), .C1(new_n1027), .C2(new_n1021), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1082), .A2(new_n1033), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n815), .B1(new_n213), .B2(new_n504), .C1(new_n808), .C2(new_n248), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n803), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT113), .Z(new_n1088));
  NOR2_X1   g0888(.A1(new_n986), .A2(new_n821), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n779), .A2(new_n399), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n336), .B1(new_n741), .B2(new_n833), .C1(new_n748), .C2(new_n202), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n783), .A2(new_n272), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G87), .C2(new_n756), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n760), .A2(new_n834), .B1(new_n973), .B2(new_n746), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n318), .C2(new_n774), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n748), .A2(new_n620), .B1(new_n751), .B2(new_n626), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n766), .B2(G294), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT114), .Z(new_n1099));
  OAI21_X1  g0899(.A(new_n282), .B1(new_n1056), .B2(new_n741), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n787), .B(new_n1100), .C1(new_n775), .C2(G283), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n761), .A2(G311), .B1(G317), .B2(new_n831), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1090), .A2(new_n1096), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1088), .B(new_n1089), .C1(new_n797), .C2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1085), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1084), .A2(new_n1107), .ZN(G390));
  OAI21_X1  g0908(.A(new_n712), .B1(new_n672), .B2(new_n563), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n666), .B1(new_n662), .B2(new_n664), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n693), .B(new_n851), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n853), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n923), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n901), .C1(new_n687), .C2(new_n912), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n913), .B1(new_n915), .B2(new_n923), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n902), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n859), .C1(new_n937), .C2(new_n944), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n936), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n933), .A2(new_n923), .A3(G330), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1114), .B(new_n1120), .C1(new_n1115), .C2(new_n902), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1118), .A2(new_n1112), .ZN(new_n1123));
  OAI211_X1 g0923(.A(KEYINPUT115), .B(G330), .C1(new_n937), .C2(new_n944), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n859), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT115), .B1(new_n735), .B2(G330), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n936), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1117), .A2(new_n936), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1123), .A2(new_n1127), .B1(new_n1129), .B2(new_n915), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n737), .A2(new_n928), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n660), .B(new_n1131), .C1(new_n718), .C2(new_n461), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1122), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1119), .A2(new_n1133), .A3(new_n1121), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n701), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1119), .A2(new_n1008), .A3(new_n1121), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n802), .B1(new_n399), .B2(new_n827), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n780), .A2(new_n498), .B1(G107), .B2(new_n830), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT116), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n282), .B1(new_n741), .B2(new_n750), .C1(new_n746), .C2(new_n843), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n760), .A2(new_n626), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1092), .A2(new_n837), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n792), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1141), .A2(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n775), .A2(G150), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n755), .A2(new_n202), .B1(new_n760), .B2(new_n838), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n282), .B1(new_n742), .B2(G125), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  INV_X1    g0952(.A(G137), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n746), .C1(new_n1153), .C2(new_n748), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1150), .B(new_n1154), .C1(G159), .C2(new_n782), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n779), .B2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1146), .A2(new_n1147), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT117), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n797), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1139), .B1(new_n1161), .B2(new_n1162), .C1(new_n813), .C2(new_n902), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1137), .A2(new_n1138), .A3(new_n1163), .ZN(G378));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n949), .B2(new_n932), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n947), .B1(new_n946), .B2(new_n901), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n889), .A2(new_n893), .A3(new_n947), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1168), .A2(new_n936), .A3(new_n945), .ZN(new_n1169));
  OAI211_X1 g0969(.A(KEYINPUT120), .B(G330), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n370), .A2(new_n877), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n385), .B(new_n1171), .Z(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1166), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1173), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1172), .B(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1177), .A2(new_n950), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n927), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n927), .A3(new_n1178), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n1008), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n803), .B1(G50), .B2(new_n828), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1185));
  INV_X1    g0985(.A(G41), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n282), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n755), .A2(new_n259), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n282), .B(new_n1186), .C1(new_n741), .C2(new_n843), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n775), .C2(G77), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT118), .Z(new_n1191));
  AOI22_X1  g0991(.A1(new_n830), .A2(G97), .B1(new_n831), .B2(G116), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n206), .B2(new_n760), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G68), .B2(new_n782), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1191), .B(new_n1194), .C1(new_n268), .C2(new_n767), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1187), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1156), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n775), .A2(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT119), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT119), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n830), .A2(G132), .B1(new_n831), .B2(G125), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n1152), .B2(new_n760), .C1(new_n783), .C2(new_n973), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G137), .B2(new_n766), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n756), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n742), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1197), .B1(new_n1196), .B2(new_n1195), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1184), .B1(new_n1211), .B2(new_n797), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1174), .B2(new_n813), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1183), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1132), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1136), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(new_n1181), .A3(KEYINPUT57), .A4(new_n1182), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n701), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1175), .A2(new_n927), .A3(new_n1178), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n927), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1221), .B2(new_n1216), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1214), .B1(new_n1218), .B2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1134), .A2(new_n1030), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n936), .A2(new_n812), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n828), .A2(G68), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n779), .A2(new_n206), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n775), .A2(G97), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n282), .B1(new_n741), .B2(new_n620), .C1(new_n748), .C2(new_n626), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G294), .B2(new_n831), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G77), .A2(new_n756), .B1(new_n761), .B2(G283), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1046), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n282), .B(new_n1188), .C1(G128), .C2(new_n742), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n202), .B2(new_n783), .C1(new_n834), .C2(new_n774), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G132), .A2(new_n831), .B1(new_n830), .B2(new_n1198), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1153), .B2(new_n760), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(KEYINPUT121), .A2(new_n1237), .B1(new_n766), .B2(G150), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(KEYINPUT121), .B2(new_n1237), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1228), .A2(new_n1233), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n802), .B(new_n1227), .C1(new_n1240), .C2(new_n797), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1226), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1130), .B2(new_n1033), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1225), .A2(new_n1244), .ZN(G381));
  XNOR2_X1  g1045(.A(G375), .B(KEYINPUT122), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1078), .A2(new_n825), .A3(new_n1080), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1247), .A2(G390), .A3(G384), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1248), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT123), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1246), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1251), .A2(new_n1252), .ZN(G407));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT124), .Z(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G378), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1246), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G407), .A2(new_n1259), .ZN(G409));
  OAI211_X1 g1060(.A(G378), .B(new_n1214), .C1(new_n1218), .C2(new_n1222), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1216), .A2(new_n1181), .A3(new_n1030), .A4(new_n1182), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1183), .A3(new_n1213), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(new_n1256), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1130), .A2(new_n1132), .A3(KEYINPUT60), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n701), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1224), .B1(new_n1133), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1272), .A2(new_n1244), .B1(new_n1273), .B2(G384), .ZN(new_n1274));
  OAI211_X1 g1074(.A(KEYINPUT125), .B(new_n856), .C1(new_n864), .C2(new_n865), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1243), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n865), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n863), .A3(new_n861), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n856), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1277), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1255), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1283), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1283), .A2(G2897), .A3(new_n1255), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1283), .B1(G2897), .B2(new_n1256), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1266), .A2(new_n1255), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G390), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1247), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n825), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n983), .B(G390), .C1(new_n1007), .C2(new_n1031), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1299), .A2(new_n1300), .A3(KEYINPUT61), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1284), .A2(new_n1289), .A3(new_n1292), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1303), .B1(new_n1267), .B2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1278), .A2(new_n1281), .A3(new_n1277), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1310), .A2(new_n1285), .A3(new_n1257), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1287), .A2(new_n1309), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1312), .B2(KEYINPUT126), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1287), .A2(new_n1314), .A3(new_n1309), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1305), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1299), .A2(new_n1300), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1297), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT127), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1302), .B1(new_n1316), .B2(new_n1324), .ZN(G405));
  AND2_X1   g1125(.A1(G375), .A2(new_n1262), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1261), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1283), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1324), .ZN(G402));
endmodule


