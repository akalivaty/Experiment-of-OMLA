//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT0), .A3(G128), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT0), .B(G128), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT64), .A2(G131), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n201), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n194), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(G128), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n190), .B2(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n209), .A2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(G128), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n210), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n216), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n218), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  INV_X1    g044(.A(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n201), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n198), .A2(G134), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n200), .A3(G131), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n230), .A3(new_n234), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT30), .B(new_n205), .C1(new_n229), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT66), .B(G116), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G119), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT2), .B(G113), .Z(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n226), .A2(new_n227), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n232), .A2(new_n234), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n205), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n239), .A2(new_n245), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G237), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G210), .ZN(new_n255));
  INV_X1    g069(.A(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n257), .B(new_n258), .Z(new_n259));
  XNOR2_X1  g073(.A(new_n201), .B(new_n202), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n193), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT68), .B1(new_n215), .B2(new_n216), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n226), .A2(new_n218), .A3(new_n227), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n232), .A2(new_n230), .A3(new_n234), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(new_n235), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n261), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT66), .A2(G116), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT66), .A2(G116), .ZN(new_n269));
  OAI21_X1  g083(.A(G119), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n241), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(new_n244), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n252), .A2(new_n259), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT31), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n252), .A2(new_n277), .A3(new_n259), .A4(new_n274), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n273), .B1(new_n205), .B2(new_n248), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n267), .B2(new_n273), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n283), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n245), .B(new_n261), .C1(new_n264), .C2(new_n266), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT70), .B(new_n285), .C1(new_n286), .C2(new_n281), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n286), .B2(KEYINPUT28), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n284), .A2(new_n287), .A3(new_n289), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n259), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n189), .B1(new_n279), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT73), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n298));
  INV_X1    g112(.A(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n276), .A2(new_n278), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n293), .B2(new_n292), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n298), .B(new_n299), .C1(new_n301), .C2(new_n189), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n252), .A2(new_n274), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n303), .B(new_n305), .C1(new_n292), .C2(new_n293), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n289), .A2(new_n291), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n267), .A2(new_n273), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT28), .B1(new_n308), .B2(new_n286), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n307), .A2(KEYINPUT29), .A3(new_n259), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n188), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n297), .A2(new_n302), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n188), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n319), .B2(G128), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n320), .A2(KEYINPUT23), .B1(new_n319), .B2(G128), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT75), .B(new_n322), .C1(new_n319), .C2(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G110), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n206), .A3(G119), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT74), .B1(new_n319), .B2(G128), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n319), .A2(G128), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT24), .B(G110), .Z(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G125), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT16), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT76), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n337), .A3(G140), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n339), .A2(new_n341), .B1(G125), .B2(new_n333), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n207), .B(new_n336), .C1(new_n342), .C2(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n340), .B1(new_n337), .B2(G140), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n333), .A2(KEYINPUT76), .A3(G125), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n334), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT16), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n207), .B1(new_n348), .B2(new_n336), .ZN(new_n349));
  OAI221_X1 g163(.A(new_n325), .B1(new_n330), .B2(new_n332), .C1(new_n344), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n330), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n324), .B2(G110), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT77), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n336), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G146), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n351), .B(new_n356), .C1(new_n324), .C2(G110), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n334), .A2(new_n338), .A3(new_n207), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n353), .A2(new_n355), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G137), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n350), .A2(new_n359), .A3(new_n363), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n318), .B1(new_n367), .B2(G902), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n365), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n366), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n317), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n367), .A2(G902), .A3(new_n316), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT9), .B(G234), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT78), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n188), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G221), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(new_n188), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n254), .A2(G227), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT79), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G107), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n388), .A2(KEYINPUT3), .A3(G104), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT3), .B1(new_n388), .B2(G104), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n256), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(KEYINPUT81), .A3(G104), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n388), .B2(G104), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n386), .A2(G107), .ZN(new_n395));
  OAI211_X1 g209(.A(G101), .B(new_n392), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT82), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n264), .A2(KEYINPUT10), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n388), .A2(G104), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT3), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n386), .B2(G107), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(KEYINPUT3), .A3(G104), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n256), .B1(new_n395), .B2(KEYINPUT81), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n388), .A2(G104), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n387), .A2(new_n410), .A3(new_n393), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n408), .A2(new_n256), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n215), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT80), .A2(G101), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n408), .B2(new_n256), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n408), .A2(new_n416), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n403), .A2(new_n414), .B1(new_n422), .B2(new_n194), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n402), .A2(new_n423), .A3(new_n260), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n260), .B1(new_n402), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n385), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n412), .A2(new_n215), .A3(new_n216), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n214), .A2(new_n190), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n413), .B1(new_n429), .B2(new_n221), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n397), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n204), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT12), .B(new_n204), .C1(new_n428), .C2(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n384), .A3(new_n424), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n427), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n380), .B1(new_n438), .B2(new_n379), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n424), .A2(new_n384), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n426), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n424), .A2(KEYINPUT83), .A3(new_n384), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n384), .B1(new_n436), .B2(new_n424), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(G469), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n378), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n245), .A2(new_n422), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n270), .A2(KEYINPUT5), .A3(new_n271), .ZN(new_n452));
  INV_X1    g266(.A(G113), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n241), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n452), .A2(new_n455), .B1(new_n243), .B2(new_n244), .ZN(new_n456));
  INV_X1    g270(.A(new_n400), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n399), .B1(new_n391), .B2(new_n396), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(G110), .B(G122), .Z(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n451), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G125), .B1(new_n226), .B2(new_n227), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n191), .B(G125), .C1(new_n190), .C2(new_n192), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n254), .A2(G224), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n460), .A2(new_n472), .A3(new_n461), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n455), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n243), .A2(new_n244), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n478), .B2(new_n397), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n456), .A2(KEYINPUT84), .A3(new_n412), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n397), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n461), .B(KEYINPUT8), .Z(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT85), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT7), .B(new_n470), .C1(new_n466), .C2(new_n468), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n470), .A2(KEYINPUT7), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n469), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n464), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n482), .A2(new_n490), .A3(new_n483), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n474), .A2(new_n492), .A3(new_n188), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n474), .A2(new_n492), .A3(new_n188), .A4(new_n494), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n450), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n448), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G478), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n240), .A2(G122), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT14), .A3(G107), .ZN(new_n504));
  OAI21_X1  g318(.A(G122), .B1(new_n268), .B2(new_n269), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n505), .A2(new_n388), .A3(new_n503), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n388), .B1(new_n505), .B2(new_n503), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n209), .B2(G128), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n206), .A2(KEYINPUT90), .A3(G143), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n209), .A2(G128), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n512), .A2(G134), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G134), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n505), .A2(KEYINPUT14), .A3(G107), .A4(new_n503), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n196), .B1(KEYINPUT89), .B2(new_n521), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n506), .A2(new_n507), .ZN(new_n526));
  INV_X1    g340(.A(new_n524), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n514), .B2(new_n515), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n508), .A2(new_n516), .A3(KEYINPUT91), .A4(new_n517), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n520), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n374), .A2(new_n315), .A3(G953), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n520), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n188), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n501), .B1(new_n537), .B2(KEYINPUT92), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n539));
  INV_X1    g353(.A(new_n501), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n536), .A2(new_n539), .A3(new_n188), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(G234), .A2(G237), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n542), .A2(G952), .A3(new_n254), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n542), .A2(G902), .A3(G953), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT21), .B(G898), .Z(new_n547));
  OAI21_X1  g361(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n538), .A2(new_n541), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G475), .A2(G902), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n386), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n358), .B1(new_n342), .B2(new_n207), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n253), .A2(new_n254), .A3(G214), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n209), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n253), .A2(new_n254), .A3(G143), .A4(G214), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT18), .A3(G131), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT18), .A2(G131), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n355), .A2(new_n563), .A3(new_n343), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT88), .B1(new_n344), .B2(new_n349), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT17), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n558), .B2(G131), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT86), .B1(new_n558), .B2(G131), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n558), .A2(G131), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n556), .A2(new_n571), .A3(new_n231), .A4(new_n557), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n573), .B2(new_n567), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n553), .B(new_n562), .C1(new_n566), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT19), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n334), .A2(new_n338), .A3(new_n576), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n577), .A2(KEYINPUT87), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(KEYINPUT87), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(new_n579), .C1(new_n576), .C2(new_n342), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n355), .B(new_n573), .C1(G146), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n562), .ZN(new_n582));
  INV_X1    g396(.A(new_n553), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n551), .B1(new_n575), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT20), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(KEYINPUT20), .B(new_n551), .C1(new_n575), .C2(new_n584), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n562), .B1(new_n566), .B2(new_n574), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n583), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n590), .B2(new_n575), .ZN(new_n591));
  INV_X1    g405(.A(G475), .ZN(new_n592));
  OAI22_X1  g406(.A1(new_n587), .A2(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n549), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n499), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n314), .A2(new_n372), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  OR2_X1    g412(.A1(new_n370), .A2(new_n371), .ZN(new_n599));
  INV_X1    g413(.A(new_n548), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n499), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n279), .A2(new_n294), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n187), .B1(new_n602), .B2(new_n188), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n295), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n536), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n534), .A2(KEYINPUT33), .A3(new_n535), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(G478), .A3(new_n188), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n537), .A2(new_n500), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n593), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NOR2_X1   g432(.A1(new_n587), .A2(new_n588), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT95), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n587), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n538), .A2(new_n541), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n591), .A2(new_n592), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n605), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n388), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NAND2_X1  g445(.A1(new_n368), .A2(new_n369), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n316), .A2(G902), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n360), .B(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n632), .A2(new_n316), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n603), .A2(new_n295), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n596), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  OAI21_X1  g455(.A(new_n544), .B1(new_n546), .B2(G900), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n623), .A2(new_n626), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n499), .A2(new_n637), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n314), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  NAND2_X1  g461(.A1(new_n632), .A2(new_n316), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n636), .A2(new_n633), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n593), .A2(new_n624), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n651), .A3(new_n450), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT99), .Z(new_n653));
  INV_X1    g467(.A(new_n275), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n308), .A2(new_n286), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n654), .B1(new_n293), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n657), .B2(G902), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n297), .A2(new_n302), .A3(new_n313), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n496), .A2(new_n497), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n642), .B(KEYINPUT39), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n448), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT40), .Z(new_n665));
  NAND4_X1  g479(.A1(new_n653), .A2(new_n659), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NAND3_X1  g481(.A1(new_n593), .A2(new_n611), .A3(new_n642), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n314), .A2(new_n645), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT100), .B(G146), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G48));
  NAND2_X1  g486(.A1(new_n498), .A2(new_n548), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n438), .A2(new_n379), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n436), .A2(new_n384), .A3(new_n424), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n402), .A2(new_n423), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n204), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n384), .B1(new_n677), .B2(new_n424), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n379), .B(new_n188), .C1(new_n675), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n674), .A2(new_n377), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n673), .A2(new_n680), .A3(new_n612), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n314), .A2(new_n372), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT102), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n684), .B(new_n686), .ZN(G15));
  NOR4_X1   g501(.A1(new_n673), .A2(new_n623), .A3(new_n599), .A4(new_n626), .ZN(new_n688));
  INV_X1    g502(.A(new_n498), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n680), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n314), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR2_X1   g506(.A1(new_n595), .A2(new_n637), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n314), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  AOI21_X1  g509(.A(new_n259), .B1(new_n307), .B2(new_n309), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n187), .B(new_n188), .C1(new_n696), .C2(new_n300), .ZN(new_n697));
  AOI21_X1  g511(.A(G902), .B1(new_n279), .B2(new_n294), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n697), .B(new_n372), .C1(new_n698), .C2(new_n187), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n680), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n673), .A2(new_n651), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  OAI211_X1 g517(.A(new_n650), .B(new_n697), .C1(new_n698), .C2(new_n187), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n668), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n690), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n668), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n312), .A2(new_n313), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n372), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n714));
  INV_X1    g528(.A(new_n380), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n679), .A2(new_n715), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n379), .B(new_n445), .C1(new_n442), .C2(new_n443), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n377), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n496), .A2(new_n449), .A3(new_n497), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n496), .A2(new_n449), .A3(new_n497), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n448), .A2(new_n721), .A3(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n708), .B1(new_n713), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n311), .A2(G472), .B1(new_n295), .B2(KEYINPUT32), .ZN(new_n726));
  INV_X1    g540(.A(new_n712), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n599), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n723), .A4(new_n710), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n314), .A2(new_n723), .A3(new_n372), .A4(new_n669), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n709), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n731), .B2(new_n709), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  AND2_X1   g550(.A1(new_n314), .A2(new_n372), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n644), .A3(new_n723), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  INV_X1    g554(.A(new_n611), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n593), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT43), .ZN(new_n743));
  INV_X1    g557(.A(new_n604), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n650), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n740), .B1(new_n746), .B2(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n719), .B1(new_n746), .B2(KEYINPUT44), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(KEYINPUT107), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT108), .A4(new_n750), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n444), .A2(KEYINPUT45), .A3(new_n446), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(KEYINPUT106), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT106), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n444), .B2(new_n446), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n379), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n715), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n679), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT46), .B1(new_n760), .B2(new_n715), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n377), .B(new_n663), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n753), .A2(new_n754), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OAI21_X1  g581(.A(new_n377), .B1(new_n762), .B2(new_n763), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT47), .Z(new_n769));
  NOR4_X1   g583(.A1(new_n314), .A2(new_n372), .A3(new_n668), .A4(new_n719), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n314), .B(new_n690), .C1(new_n688), .C2(new_n693), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n700), .A2(new_n701), .B1(new_n596), .B2(new_n638), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n538), .A2(KEYINPUT110), .A3(new_n541), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT110), .B1(new_n538), .B2(new_n541), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(KEYINPUT111), .B(new_n612), .C1(new_n778), .C2(new_n593), .ZN(new_n779));
  INV_X1    g593(.A(new_n593), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n780), .B(new_n781), .C1(new_n776), .C2(new_n777), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n601), .A2(new_n779), .A3(new_n604), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n774), .A2(new_n775), .A3(new_n597), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n684), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n625), .A2(new_n642), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n637), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n778), .A3(new_n622), .A4(new_n620), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n448), .A2(new_n721), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n314), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n705), .A2(KEYINPUT112), .A3(new_n723), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT112), .B1(new_n705), .B2(new_n723), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n785), .A2(new_n735), .A3(new_n738), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n689), .A2(new_n651), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n718), .A2(new_n650), .A3(new_n643), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n659), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n646), .A2(new_n670), .A3(new_n799), .A4(new_n706), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT52), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n773), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(KEYINPUT113), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n796), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n802), .A2(new_n803), .B1(new_n809), .B2(KEYINPUT53), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n684), .A2(new_n784), .A3(new_n794), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n800), .B(new_n805), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n735), .A4(new_n738), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(KEYINPUT115), .A3(new_n773), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n814), .A2(new_n773), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT114), .B1(new_n809), .B2(KEYINPUT53), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n816), .B1(new_n821), .B2(new_n811), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n680), .A2(new_n719), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n372), .A3(new_n543), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n659), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n780), .A3(new_n741), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n743), .A2(new_n543), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n450), .B1(new_n828), .B2(KEYINPUT50), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n662), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n700), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(new_n828), .A3(KEYINPUT50), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n828), .B2(KEYINPUT50), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n823), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n704), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n699), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n721), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n674), .A2(new_n679), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n769), .B1(new_n378), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n826), .B(new_n836), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n827), .A2(new_n728), .A3(new_n823), .ZN(new_n849));
  XOR2_X1   g663(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n850));
  OR2_X1    g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n254), .A2(G952), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n838), .B2(new_n690), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n825), .A2(new_n613), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n850), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n847), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n822), .A2(new_n857), .B1(G952), .B2(G953), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n599), .A2(new_n450), .A3(new_n378), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n859), .B(new_n742), .C1(new_n860), .C2(new_n842), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n662), .B1(new_n860), .B2(new_n842), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n858), .B1(new_n659), .B2(new_n866), .ZN(G75));
  AOI21_X1  g681(.A(new_n188), .B1(new_n810), .B2(new_n815), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(G210), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n465), .A2(new_n473), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n471), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT55), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n869), .B2(new_n870), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n254), .A2(G952), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G51));
  NAND2_X1  g691(.A1(new_n802), .A2(new_n803), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n815), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n816), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n380), .B(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n678), .B2(new_n675), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n868), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n876), .B1(new_n885), .B2(new_n886), .ZN(G54));
  NAND3_X1  g701(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n575), .A2(new_n584), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n890), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(new_n892), .A3(new_n876), .ZN(G60));
  AND2_X1   g707(.A1(new_n607), .A2(new_n608), .ZN(new_n894));
  NAND2_X1  g708(.A1(G478), .A2(G902), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT59), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n822), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n882), .A2(new_n894), .A3(new_n896), .ZN(new_n898));
  INV_X1    g712(.A(new_n876), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(G63));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  INV_X1    g716(.A(new_n367), .ZN(new_n903));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n880), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n907), .B2(new_n876), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n810), .B2(new_n815), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT120), .B(new_n899), .C1(new_n909), .C2(new_n903), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n880), .A2(new_n636), .A3(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n899), .B1(new_n909), .B2(new_n903), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n880), .A2(new_n906), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n876), .B1(new_n919), .B2(new_n367), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n911), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n914), .A2(new_n922), .ZN(G66));
  AOI21_X1  g737(.A(new_n254), .B1(new_n547), .B2(G224), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n785), .B(KEYINPUT122), .Z(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n254), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n871), .B1(G898), .B2(new_n254), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n926), .B(new_n927), .Z(G69));
  AND3_X1   g742(.A1(new_n646), .A2(new_n670), .A3(new_n706), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n666), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n664), .A2(new_n719), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n737), .A2(new_n779), .A3(new_n782), .A4(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n766), .A2(new_n771), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n254), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n239), .A2(new_n251), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n580), .Z(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT123), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(G900), .B2(G953), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n735), .A2(new_n738), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n765), .A2(new_n728), .A3(new_n797), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(new_n929), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n766), .A2(new_n771), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n945), .B2(G953), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n254), .B1(G227), .B2(G900), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n940), .A2(new_n950), .A3(new_n946), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n949), .B1(new_n948), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(G72));
  XNOR2_X1  g768(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n945), .B2(new_n925), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n304), .A2(new_n259), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n876), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n305), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n961), .B2(new_n654), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n821), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n957), .B1(new_n935), .B2(new_n925), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n957), .C1(new_n935), .C2(new_n925), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(new_n259), .A3(new_n304), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(G57));
endmodule


