//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(G136), .B2(new_n470), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n471), .C1(new_n463), .C2(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(G126), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT67), .B1(new_n471), .B2(G114), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT68), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  AOI211_X1 g070(.A(new_n495), .B(new_n492), .C1(new_n487), .C2(new_n490), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n486), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n486), .B(new_n499), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n485), .B1(new_n498), .B2(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT70), .B(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n507), .A2(KEYINPUT72), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT73), .Z(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n507), .B2(KEYINPUT72), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(G651), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n517), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n506), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n513), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n512), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n519), .A2(new_n520), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  OR3_X1    g105(.A1(new_n529), .A2(KEYINPUT74), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT7), .Z(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n535), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n523), .A2(new_n542), .B1(new_n502), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n532), .B2(G52), .ZN(G171));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n523), .A2(new_n546), .B1(new_n502), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n532), .B2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n505), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n523), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n522), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n529), .A2(new_n530), .ZN(new_n566));
  INV_X1    g141(.A(new_n563), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(G53), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n560), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n529), .A2(new_n505), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G91), .B1(G651), .B2(new_n557), .ZN(new_n573));
  INV_X1    g148(.A(new_n568), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n567), .B1(new_n566), .B2(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  NAND2_X1  g155(.A1(new_n566), .A2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n572), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n566), .A2(G48), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n572), .A2(G86), .ZN(new_n586));
  INV_X1    g161(.A(new_n502), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n506), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT77), .Z(new_n590));
  OAI21_X1  g165(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(G305));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n523), .A2(new_n593), .B1(new_n502), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n532), .B2(G47), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(KEYINPUT78), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n523), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n572), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n505), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n603), .A2(new_n604), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n528), .A2(KEYINPUT79), .A3(new_n531), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G54), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT79), .B1(new_n528), .B2(new_n531), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n578), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n578), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n465), .A2(new_n472), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n470), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n478), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n471), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT81), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(G2072), .A2(G2078), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n442), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n658), .A2(KEYINPUT82), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(KEYINPUT82), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n664), .A3(new_n660), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n658), .B(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n656), .C1(new_n666), .C2(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n660), .A3(new_n655), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT83), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT84), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n681), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  OAI211_X1 g259(.A(new_n682), .B(new_n684), .C1(new_n681), .C2(new_n676), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  INV_X1    g267(.A(G34), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(KEYINPUT24), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(KEYINPUT24), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G160), .B2(new_n692), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT93), .B(G2084), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G2067), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n692), .A2(G26), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  AOI22_X1  g278(.A1(G128), .A2(new_n478), .B1(new_n470), .B2(G140), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n707));
  OAI221_X1 g282(.A(G2104), .B1(G116), .B2(new_n471), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(G29), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n470), .A2(G139), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT91), .Z(new_n713));
  NAND3_X1  g288(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT25), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n713), .B(new_n716), .C1(new_n471), .C2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G33), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n721), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n720), .A2(G2072), .B1(G1961), .B2(new_n723), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n478), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT26), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G32), .B(new_n729), .S(G29), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT94), .B(KEYINPUT31), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G11), .ZN(new_n734));
  INV_X1    g309(.A(G28), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(KEYINPUT95), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(KEYINPUT95), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n736), .A2(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n734), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n744), .B1(new_n692), .B2(new_n636), .C1(new_n710), .C2(new_n701), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n732), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G35), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G162), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AND4_X1   g326(.A1(new_n711), .A2(new_n724), .A3(new_n746), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n721), .A2(G20), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT23), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n721), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n549), .B2(new_n721), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT89), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1341), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n692), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n692), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n752), .A2(new_n756), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n613), .A2(new_n721), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G4), .B2(new_n721), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT88), .B(G1348), .Z(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n721), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n721), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n774), .B1(G1961), .B2(new_n723), .C1(new_n720), .C2(G2072), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n765), .A2(new_n769), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n692), .A2(G25), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT85), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n470), .A2(G131), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n478), .A2(G119), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n471), .A2(G107), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n780), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT86), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT86), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n779), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT35), .B(G1991), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n721), .A2(G24), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G290), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1986), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n721), .A2(G23), .ZN(new_n795));
  INV_X1    g370(.A(G288), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n721), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT33), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1976), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n721), .A2(G22), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT87), .Z(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G303), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(G6), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G305), .B2(new_n721), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT32), .B(G1981), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n808), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n802), .A2(new_n803), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n799), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OAI221_X1 g387(.A(new_n794), .B1(KEYINPUT34), .B2(new_n812), .C1(new_n793), .C2(new_n792), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(KEYINPUT34), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT36), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n777), .A2(new_n816), .ZN(G311));
  OR2_X1    g392(.A1(new_n777), .A2(new_n816), .ZN(G150));
  NAND2_X1  g393(.A1(new_n613), .A2(G559), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n523), .A2(new_n822), .B1(new_n502), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n532), .B2(G55), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n549), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n549), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n821), .B(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n825), .A2(new_n832), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n709), .B(KEYINPUT100), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n718), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n787), .B(new_n627), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n497), .B2(new_n485), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n471), .A2(KEYINPUT67), .A3(G114), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n493), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n495), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n491), .A2(KEYINPUT68), .A3(new_n493), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n483), .B(KEYINPUT4), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT99), .A4(new_n486), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n729), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n478), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n471), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G142), .B2(new_n470), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n841), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n474), .B(new_n636), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n860), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(G395));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n597), .A2(new_n796), .A3(new_n598), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n796), .B1(new_n597), .B2(new_n598), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(G290), .A2(G288), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n597), .A2(new_n796), .A3(new_n598), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(KEYINPUT105), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(G303), .B(G305), .Z(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n876), .A2(KEYINPUT105), .A3(new_n871), .A4(new_n872), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n875), .A2(KEYINPUT106), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT106), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n621), .B(new_n828), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n578), .A2(new_n612), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  INV_X1    g461(.A(new_n611), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(G54), .A3(new_n609), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n888), .A2(new_n571), .A3(new_n577), .A4(new_n608), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(G299), .A2(new_n613), .A3(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n885), .A2(new_n895), .A3(new_n889), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n578), .A2(KEYINPUT103), .A3(new_n612), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n890), .B2(new_n891), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n894), .B1(new_n884), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n875), .A2(new_n877), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n882), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n875), .A2(KEYINPUT106), .A3(new_n877), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  INV_X1    g487(.A(new_n905), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n825), .A2(G868), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G295));
  INV_X1    g493(.A(G868), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n903), .B1(new_n882), .B2(new_n905), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(new_n907), .A3(new_n913), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT107), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n915), .A2(new_n924), .A3(new_n917), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(G301), .A2(KEYINPUT108), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(G286), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(G168), .A2(new_n930), .A3(G171), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n828), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n829), .A2(new_n933), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n899), .B2(new_n901), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n937), .B(KEYINPUT109), .C1(new_n899), .C2(new_n901), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n934), .B2(new_n828), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n936), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n892), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n950), .B2(new_n911), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n940), .A2(new_n941), .B1(new_n948), .B2(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n880), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n928), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n952), .B2(new_n880), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n935), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n943), .A2(new_n947), .A3(new_n945), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n893), .B2(new_n900), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n960), .B2(new_n911), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n927), .B1(new_n954), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n927), .B1(new_n951), .B2(new_n955), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n953), .A2(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n964), .A2(KEYINPUT111), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT111), .B1(new_n964), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(G397));
  XNOR2_X1  g544(.A(new_n787), .B(new_n789), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT113), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n709), .B(new_n701), .ZN(new_n972));
  INV_X1    g547(.A(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n729), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n852), .A2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n468), .A2(G40), .A3(new_n473), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n981), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n985));
  OAI22_X1  g560(.A1(new_n976), .A2(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n984), .B2(new_n985), .ZN(new_n987));
  INV_X1    g562(.A(new_n981), .ZN(new_n988));
  INV_X1    g563(.A(new_n972), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n729), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n973), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(KEYINPUT46), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(KEYINPUT46), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  NAND3_X1  g570(.A1(new_n785), .A2(new_n789), .A3(new_n786), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n975), .A2(new_n996), .B1(G2067), .B2(new_n709), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n987), .B(new_n995), .C1(new_n988), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n847), .A2(new_n848), .B1(G126), .B2(new_n478), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n1000), .B2(new_n850), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n979), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n1002), .B2(G8), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n999), .A3(G8), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1005), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n585), .A2(new_n586), .A3(new_n1010), .A4(new_n591), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1009), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n1007), .A2(new_n1003), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n796), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1011), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1006), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n796), .A2(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1019), .B(new_n1020), .C1(new_n1007), .C2(new_n1003), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n1006), .B2(new_n1019), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G303), .A2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n468), .A2(G40), .A3(new_n473), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1001), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT115), .B1(new_n1034), .B2(G2090), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1030), .A2(new_n1036), .A3(new_n750), .A4(new_n1033), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n499), .B1(new_n849), .B2(new_n486), .ZN(new_n1039));
  INV_X1    g614(.A(new_n500), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n850), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n977), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1031), .B1(new_n1042), .B2(new_n980), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n843), .A2(new_n851), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n843), .A2(new_n851), .A3(new_n1047), .A4(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1971), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(new_n1029), .C1(new_n1038), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1018), .B1(new_n1026), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1051), .A2(new_n1025), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1043), .A2(new_n763), .A3(new_n1049), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  INV_X1    g630(.A(G1961), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1054), .A2(new_n1055), .B1(new_n1056), .B2(new_n1034), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n979), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n498), .A2(new_n500), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1384), .B1(new_n1059), .B2(new_n850), .ZN(new_n1060));
  INV_X1    g635(.A(new_n980), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1055), .A2(G2078), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(G171), .B(KEYINPUT54), .Z(new_n1066));
  NAND2_X1  g641(.A1(new_n979), .A2(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n978), .B2(new_n980), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(new_n1049), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1065), .A2(new_n1066), .B1(new_n1057), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1029), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n977), .B1(new_n497), .B2(new_n485), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1031), .B1(new_n1072), .B2(KEYINPUT50), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(G2090), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1050), .A2(new_n1075), .A3(KEYINPUT117), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1071), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1053), .A2(new_n1070), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1049), .A2(new_n973), .A3(new_n979), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1002), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1001), .A2(new_n979), .A3(KEYINPUT122), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT58), .B(G1341), .Z(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n549), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1091), .A3(new_n549), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1032), .B1(new_n1041), .B2(new_n977), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1033), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n768), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT122), .B1(new_n1001), .B2(new_n979), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1072), .A2(new_n1031), .A3(new_n1083), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n701), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1095), .A2(new_n613), .A3(KEYINPUT60), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  INV_X1    g675(.A(new_n768), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1102));
  AOI21_X1  g677(.A(G2067), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1098), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n612), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1090), .A2(new_n1092), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(KEYINPUT57), .C1(new_n569), .C2(KEYINPUT119), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT120), .B1(new_n576), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n576), .B2(KEYINPUT120), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1110), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1043), .A2(new_n1049), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1074), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT61), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(KEYINPUT121), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1117), .A2(new_n1115), .A3(new_n1119), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1120), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1108), .B(new_n1123), .C1(new_n1127), .C2(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n612), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1120), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1080), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G2084), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1033), .C1(new_n1060), .C2(new_n1032), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1062), .B2(G1966), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT51), .B(G8), .C1(new_n1135), .C2(G286), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G8), .ZN(new_n1139));
  NOR3_X1   g714(.A1(G164), .A2(G1384), .A3(new_n980), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n773), .B1(new_n1140), .B2(new_n1058), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1141), .B2(new_n1134), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G168), .A2(new_n1139), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(G168), .B2(new_n1139), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1135), .A2(G8), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1147), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(KEYINPUT124), .A3(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1138), .A2(new_n1144), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1135), .A2(new_n1143), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1152), .A2(KEYINPUT125), .A3(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1052), .B1(new_n1132), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1152), .A2(KEYINPUT125), .A3(new_n1153), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT125), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT62), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1156), .A2(new_n1163), .A3(new_n1157), .ZN(new_n1164));
  AND4_X1   g739(.A1(G171), .A2(new_n1053), .A3(new_n1079), .A4(new_n1065), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1149), .A2(G286), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1053), .A2(new_n1079), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT118), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1172), .A3(new_n1169), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1071), .B1(new_n1174), .B2(new_n1139), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1053), .A2(KEYINPUT63), .A3(new_n1167), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1171), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1159), .A2(new_n1166), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n1179));
  NAND2_X1  g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n976), .A2(new_n983), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n988), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1179), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n998), .B1(new_n1183), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g760(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1187), .A2(new_n864), .ZN(new_n1188));
  NOR2_X1   g762(.A1(new_n954), .A2(new_n962), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n1188), .A2(new_n1189), .ZN(G308));
  OR2_X1    g764(.A1(new_n1188), .A2(new_n1189), .ZN(G225));
endmodule


