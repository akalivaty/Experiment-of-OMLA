

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XOR2_X1 U321 ( .A(n393), .B(n392), .Z(n524) );
  XNOR2_X1 U322 ( .A(n392), .B(n349), .ZN(n350) );
  XOR2_X1 U323 ( .A(n439), .B(n438), .Z(n289) );
  INV_X1 U324 ( .A(n397), .ZN(n398) );
  INV_X1 U325 ( .A(KEYINPUT90), .ZN(n374) );
  XNOR2_X1 U326 ( .A(n375), .B(n374), .ZN(n394) );
  NAND2_X1 U327 ( .A1(n394), .A2(n524), .ZN(n408) );
  XNOR2_X1 U328 ( .A(n510), .B(KEYINPUT27), .ZN(n397) );
  INV_X1 U329 ( .A(KEYINPUT121), .ZN(n465) );
  XNOR2_X1 U330 ( .A(n440), .B(n289), .ZN(n441) );
  XNOR2_X1 U331 ( .A(n465), .B(KEYINPUT55), .ZN(n466) );
  XNOR2_X1 U332 ( .A(n348), .B(G204GAT), .ZN(n349) );
  XNOR2_X1 U333 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U334 ( .A(n467), .B(n466), .ZN(n468) );
  INV_X1 U335 ( .A(G50GAT), .ZN(n446) );
  XNOR2_X1 U336 ( .A(KEYINPUT38), .B(n445), .ZN(n490) );
  XNOR2_X1 U337 ( .A(n469), .B(G176GAT), .ZN(n470) );
  XNOR2_X1 U338 ( .A(n446), .B(KEYINPUT102), .ZN(n447) );
  XNOR2_X1 U339 ( .A(n471), .B(n470), .ZN(G1349GAT) );
  XNOR2_X1 U340 ( .A(n448), .B(n447), .ZN(G1331GAT) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G162GAT), .Z(n329) );
  XOR2_X1 U342 ( .A(G211GAT), .B(KEYINPUT82), .Z(n291) );
  XNOR2_X1 U343 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n344) );
  XNOR2_X1 U345 ( .A(n329), .B(n344), .ZN(n292) );
  XOR2_X1 U346 ( .A(G22GAT), .B(G155GAT), .Z(n309) );
  XNOR2_X1 U347 ( .A(n292), .B(n309), .ZN(n298) );
  XOR2_X1 U348 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n294) );
  XNOR2_X1 U349 ( .A(G141GAT), .B(KEYINPUT83), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n371) );
  XOR2_X1 U351 ( .A(n371), .B(KEYINPUT23), .Z(n296) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U354 ( .A(n298), .B(n297), .Z(n306) );
  XOR2_X1 U355 ( .A(G148GAT), .B(G106GAT), .Z(n300) );
  XNOR2_X1 U356 ( .A(G204GAT), .B(G78GAT), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U358 ( .A(KEYINPUT70), .B(n301), .ZN(n443) );
  XOR2_X1 U359 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n303) );
  XNOR2_X1 U360 ( .A(G218GAT), .B(KEYINPUT24), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U362 ( .A(n443), .B(n304), .Z(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n464) );
  XOR2_X1 U364 ( .A(n464), .B(KEYINPUT28), .Z(n523) );
  XOR2_X1 U365 ( .A(G211GAT), .B(G71GAT), .Z(n308) );
  XNOR2_X1 U366 ( .A(G183GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n322) );
  XOR2_X1 U368 ( .A(G57GAT), .B(KEYINPUT13), .Z(n436) );
  XOR2_X1 U369 ( .A(n436), .B(n309), .Z(n311) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U372 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n313) );
  XNOR2_X1 U373 ( .A(KEYINPUT15), .B(KEYINPUT73), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U375 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U376 ( .A(G15GAT), .B(G8GAT), .Z(n413) );
  XOR2_X1 U377 ( .A(KEYINPUT12), .B(G64GAT), .Z(n317) );
  XNOR2_X1 U378 ( .A(G1GAT), .B(G78GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n413), .B(n318), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n572) );
  INV_X1 U383 ( .A(n572), .ZN(n546) );
  XOR2_X1 U384 ( .A(G29GAT), .B(G43GAT), .Z(n324) );
  XNOR2_X1 U385 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n418) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n325), .B(G218GAT), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n418), .B(n340), .ZN(n338) );
  XOR2_X1 U390 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n327) );
  XNOR2_X1 U391 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U393 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n334) );
  XOR2_X1 U396 ( .A(KEYINPUT71), .B(G92GAT), .Z(n333) );
  XNOR2_X1 U397 ( .A(G99GAT), .B(G85GAT), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n433) );
  XOR2_X1 U399 ( .A(n334), .B(n433), .Z(n336) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U402 ( .A(n338), .B(n337), .Z(n558) );
  XNOR2_X1 U403 ( .A(KEYINPUT100), .B(KEYINPUT36), .ZN(n339) );
  XOR2_X1 U404 ( .A(n558), .B(n339), .Z(n578) );
  XOR2_X1 U405 ( .A(n340), .B(G8GAT), .Z(n342) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n351) );
  XOR2_X1 U409 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n346) );
  XNOR2_X1 U410 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U412 ( .A(G169GAT), .B(n347), .Z(n392) );
  XOR2_X1 U413 ( .A(G176GAT), .B(G64GAT), .Z(n437) );
  XOR2_X1 U414 ( .A(n437), .B(G92GAT), .Z(n348) );
  XOR2_X1 U415 ( .A(n351), .B(n350), .Z(n510) );
  XOR2_X1 U416 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n353) );
  XNOR2_X1 U417 ( .A(G148GAT), .B(G155GAT), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U419 ( .A(G57GAT), .B(KEYINPUT87), .Z(n355) );
  XNOR2_X1 U420 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U422 ( .A(n357), .B(n356), .Z(n368) );
  XOR2_X1 U423 ( .A(KEYINPUT85), .B(KEYINPUT1), .Z(n359) );
  XNOR2_X1 U424 ( .A(KEYINPUT86), .B(KEYINPUT6), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n366) );
  XOR2_X1 U426 ( .A(G113GAT), .B(G1GAT), .Z(n414) );
  XOR2_X1 U427 ( .A(G85GAT), .B(G162GAT), .Z(n361) );
  XNOR2_X1 U428 ( .A(G29GAT), .B(G120GAT), .ZN(n360) );
  XNOR2_X1 U429 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U430 ( .A(n414), .B(n362), .Z(n364) );
  NAND2_X1 U431 ( .A1(G225GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n373) );
  XOR2_X1 U435 ( .A(G127GAT), .B(KEYINPUT75), .Z(n370) );
  XNOR2_X1 U436 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n376) );
  XOR2_X1 U438 ( .A(n376), .B(n371), .Z(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n507) );
  NOR2_X1 U440 ( .A1(n397), .A2(n507), .ZN(n520) );
  NAND2_X1 U441 ( .A1(n520), .A2(n523), .ZN(n375) );
  XOR2_X1 U442 ( .A(G120GAT), .B(G71GAT), .Z(n432) );
  XOR2_X1 U443 ( .A(n432), .B(n376), .Z(n378) );
  XNOR2_X1 U444 ( .A(G99GAT), .B(G190GAT), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n380) );
  XNOR2_X1 U447 ( .A(G43GAT), .B(G113GAT), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U449 ( .A(KEYINPUT77), .B(G176GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U452 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U453 ( .A(KEYINPUT79), .B(KEYINPUT76), .Z(n386) );
  NAND2_X1 U454 ( .A1(G227GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U456 ( .A(KEYINPUT78), .B(n387), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n393) );
  NAND2_X1 U459 ( .A1(n524), .A2(n464), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n395), .B(KEYINPUT26), .ZN(n396) );
  XNOR2_X1 U461 ( .A(KEYINPUT91), .B(n396), .ZN(n562) );
  NAND2_X1 U462 ( .A1(n562), .A2(n398), .ZN(n405) );
  OR2_X1 U463 ( .A1(n524), .A2(n510), .ZN(n399) );
  XOR2_X1 U464 ( .A(KEYINPUT92), .B(n399), .Z(n400) );
  NOR2_X1 U465 ( .A1(n464), .A2(n400), .ZN(n403) );
  XOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n401) );
  XNOR2_X1 U467 ( .A(KEYINPUT25), .B(n401), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  NAND2_X1 U469 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n406), .A2(n507), .ZN(n407) );
  NAND2_X1 U471 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n409), .B(KEYINPUT95), .ZN(n474) );
  NOR2_X1 U473 ( .A1(n578), .A2(n474), .ZN(n410) );
  NAND2_X1 U474 ( .A1(n546), .A2(n410), .ZN(n411) );
  XNOR2_X1 U475 ( .A(KEYINPUT101), .B(n411), .ZN(n412) );
  XOR2_X1 U476 ( .A(KEYINPUT37), .B(n412), .Z(n506) );
  XOR2_X1 U477 ( .A(G36GAT), .B(G50GAT), .Z(n416) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U480 ( .A(n417), .B(G141GAT), .Z(n423) );
  XOR2_X1 U481 ( .A(n418), .B(KEYINPUT29), .Z(n420) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n431) );
  XOR2_X1 U486 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n425) );
  XNOR2_X1 U487 ( .A(G197GAT), .B(G22GAT), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U489 ( .A(KEYINPUT64), .B(KEYINPUT67), .Z(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT65), .B(KEYINPUT68), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U492 ( .A(n429), .B(n428), .Z(n430) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n540) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n435) );
  AND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n440) );
  XOR2_X1 U498 ( .A(KEYINPUT32), .B(KEYINPUT69), .Z(n439) );
  XNOR2_X1 U499 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n569) );
  NOR2_X1 U501 ( .A1(n540), .A2(n569), .ZN(n476) );
  NAND2_X1 U502 ( .A1(n506), .A2(n476), .ZN(n445) );
  NOR2_X1 U503 ( .A1(n523), .A2(n490), .ZN(n448) );
  XOR2_X1 U504 ( .A(n569), .B(KEYINPUT41), .Z(n528) );
  INV_X1 U505 ( .A(n528), .ZN(n542) );
  NOR2_X1 U506 ( .A1(n540), .A2(n542), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n449), .B(KEYINPUT46), .ZN(n450) );
  NOR2_X1 U508 ( .A1(n572), .A2(n450), .ZN(n451) );
  INV_X1 U509 ( .A(n558), .ZN(n550) );
  NAND2_X1 U510 ( .A1(n451), .A2(n550), .ZN(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT112), .B(KEYINPUT47), .Z(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n458) );
  NOR2_X1 U513 ( .A1(n578), .A2(n546), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT45), .B(n454), .Z(n455) );
  NOR2_X1 U515 ( .A1(n569), .A2(n455), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n456), .A2(n540), .ZN(n457) );
  NAND2_X1 U517 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT48), .ZN(n521) );
  INV_X1 U519 ( .A(n510), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n521), .A2(n460), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n463), .A2(n507), .ZN(n563) );
  NOR2_X1 U524 ( .A1(n464), .A2(n563), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n524), .A2(n468), .ZN(n559) );
  NAND2_X1 U526 ( .A1(n559), .A2(n528), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n469) );
  NOR2_X1 U528 ( .A1(n546), .A2(n558), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  NOR2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT96), .B(n475), .ZN(n493) );
  NAND2_X1 U532 ( .A1(n476), .A2(n493), .ZN(n483) );
  NOR2_X1 U533 ( .A1(n507), .A2(n483), .ZN(n477) );
  XOR2_X1 U534 ( .A(n477), .B(KEYINPUT34), .Z(n478) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NOR2_X1 U536 ( .A1(n510), .A2(n483), .ZN(n479) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n524), .A2(n483), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT97), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U541 ( .A(G15GAT), .B(n482), .Z(G1326GAT) );
  NOR2_X1 U542 ( .A1(n523), .A2(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  NOR2_X1 U546 ( .A1(n490), .A2(n507), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n490), .A2(n510), .ZN(n489) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n489), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n490), .A2(n524), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(n491), .Z(n492) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n492), .ZN(G1330GAT) );
  INV_X1 U554 ( .A(n540), .ZN(n565) );
  NOR2_X1 U555 ( .A1(n565), .A2(n542), .ZN(n505) );
  AND2_X1 U556 ( .A1(n493), .A2(n505), .ZN(n494) );
  XOR2_X1 U557 ( .A(KEYINPUT104), .B(n494), .Z(n502) );
  NOR2_X1 U558 ( .A1(n502), .A2(n507), .ZN(n496) );
  XNOR2_X1 U559 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n497), .ZN(G1332GAT) );
  NOR2_X1 U562 ( .A1(n502), .A2(n510), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(G1333GAT) );
  NOR2_X1 U565 ( .A1(n502), .A2(n524), .ZN(n500) );
  XOR2_X1 U566 ( .A(KEYINPUT106), .B(n500), .Z(n501) );
  XNOR2_X1 U567 ( .A(G71GAT), .B(n501), .ZN(G1334GAT) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n504) );
  NOR2_X1 U569 ( .A1(n523), .A2(n502), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NAND2_X1 U571 ( .A1(n506), .A2(n505), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n507), .A2(n517), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U575 ( .A1(n510), .A2(n517), .ZN(n511) );
  XOR2_X1 U576 ( .A(G92GAT), .B(n511), .Z(G1337GAT) );
  NOR2_X1 U577 ( .A1(n524), .A2(n517), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(n514), .ZN(G1338GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n516) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n519) );
  NOR2_X1 U584 ( .A1(n523), .A2(n517), .ZN(n518) );
  XOR2_X1 U585 ( .A(n519), .B(n518), .Z(G1339GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT113), .ZN(n539) );
  NAND2_X1 U588 ( .A1(n523), .A2(n539), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT114), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n535), .A2(n565), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U594 ( .A1(n528), .A2(n535), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n531), .Z(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n533) );
  NAND2_X1 U598 ( .A1(n535), .A2(n572), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U602 ( .A1(n535), .A2(n558), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n538), .Z(G1343GAT) );
  NAND2_X1 U605 ( .A1(n539), .A2(n562), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n540), .A2(n549), .ZN(n541) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n549), .ZN(n544) );
  XNOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n549), .ZN(n547) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(n547), .Z(n548) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n559), .A2(n565), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U621 ( .A1(n572), .A2(n559), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT123), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(n557), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  INV_X1 U629 ( .A(n562), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U635 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n576), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n580) );
  INV_X1 U642 ( .A(n576), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1355GAT) );
endmodule

