//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1227,
    new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n448), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(G137), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n468), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT68), .B1(new_n468), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G101), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n467), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n468), .B1(new_n481), .B2(new_n483), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n465), .B2(new_n466), .ZN(new_n493));
  AND2_X1   g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n468), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n465), .B2(new_n466), .ZN(new_n497));
  AND2_X1   g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n468), .C1(new_n474), .C2(new_n475), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT70), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(G88), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n507), .A2(new_n509), .A3(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n515), .B2(new_n516), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n528), .B(G62), .C1(new_n511), .C2(new_n512), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(G651), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G62), .B1(new_n511), .B2(new_n512), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n506), .B1(new_n536), .B2(new_n530), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n524), .A2(new_n534), .A3(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND2_X1  g115(.A1(new_n514), .A2(new_n519), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n521), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n518), .A2(KEYINPUT73), .A3(G543), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G51), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n551));
  AND2_X1   g126(.A1(G63), .A2(G651), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n517), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n543), .A2(new_n548), .A3(new_n553), .ZN(G168));
  AOI22_X1  g129(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n506), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n514), .A2(G90), .A3(new_n519), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT74), .B(G52), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n545), .A2(new_n546), .A3(new_n558), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n557), .A2(KEYINPUT75), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT75), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G171));
  NAND2_X1  g138(.A1(new_n547), .A2(G43), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n514), .A2(G81), .A3(new_n519), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n506), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT77), .Z(G188));
  NAND3_X1  g151(.A1(new_n514), .A2(G91), .A3(new_n519), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(KEYINPUT9), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n522), .B(new_n580), .C1(new_n579), .C2(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n513), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n586));
  OAI211_X1 g161(.A(KEYINPUT78), .B(new_n586), .C1(new_n521), .C2(new_n578), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n577), .A2(new_n581), .A3(new_n585), .A4(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n590), .B(new_n556), .C1(new_n560), .C2(new_n561), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G301));
  NAND3_X1  g168(.A1(new_n543), .A2(new_n548), .A3(new_n553), .ZN(G286));
  INV_X1    g169(.A(G74), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n506), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(G49), .B2(new_n522), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n514), .A2(G87), .A3(new_n519), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n513), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n522), .B2(G48), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n514), .A2(G86), .A3(new_n519), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n547), .A2(G47), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI221_X1 g184(.A(new_n607), .B1(new_n608), .B2(new_n541), .C1(new_n506), .C2(new_n609), .ZN(G290));
  NAND3_X1  g185(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n541), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT80), .B(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n513), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n547), .A2(G54), .B1(G651), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  MUX2_X1   g201(.A(G301), .B(new_n625), .S(new_n626), .Z(G284));
  MUX2_X1   g202(.A(G301), .B(new_n625), .S(new_n626), .Z(G321));
  NAND2_X1  g203(.A1(G299), .A2(new_n626), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G168), .B2(new_n626), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(G168), .B2(new_n626), .ZN(G280));
  INV_X1    g206(.A(new_n625), .ZN(new_n632));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n636), .A2(KEYINPUT82), .B1(new_n626), .B2(new_n568), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(KEYINPUT82), .B2(new_n636), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g214(.A1(new_n470), .A2(new_n471), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(new_n467), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n484), .A2(G135), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n486), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n663), .B(KEYINPUT85), .Z(new_n672));
  INV_X1    g247(.A(new_n665), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n669), .B1(new_n674), .B2(new_n666), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n657), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n670), .B1(new_n667), .B2(new_n668), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n669), .A3(new_n666), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n656), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(G14), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2084), .B(G2090), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(KEYINPUT17), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2072), .B(G2078), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n685), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G2096), .B(G2100), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1956), .B(G2474), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1961), .B(G1966), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT20), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  INV_X1    g282(.A(new_n704), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(new_n710), .B(new_n709), .S(new_n701), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n706), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n697), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(new_n697), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n716), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1991), .B(G1996), .ZN(new_n719));
  INV_X1    g294(.A(G1981), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n715), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n715), .B2(new_n718), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(G229));
  INV_X1    g299(.A(G28), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n725), .B2(KEYINPUT30), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n726), .A2(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n732), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n730), .B1(new_n731), .B2(new_n651), .C1(new_n734), .C2(G1966), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(G1966), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT97), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n732), .A2(G5), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G171), .B2(new_n732), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT98), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n735), .B(new_n737), .C1(new_n740), .C2(G1961), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT99), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n732), .A2(G4), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n632), .B2(new_n732), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1348), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n732), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n569), .B2(new_n732), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1341), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n731), .A2(G27), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT100), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n731), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G2078), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(G2078), .ZN(new_n754));
  AND2_X1   g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n731), .B1(KEYINPUT24), .B2(G34), .ZN(new_n756));
  OAI22_X1  g331(.A1(G160), .A2(new_n731), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2084), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n749), .A2(new_n753), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n731), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n486), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n640), .B2(G105), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n640), .A2(new_n766), .A3(G105), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n768), .A2(new_n769), .B1(G141), .B2(new_n484), .ZN(new_n770));
  AOI21_X1  g345(.A(KEYINPUT95), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n484), .A2(G141), .ZN(new_n772));
  INV_X1    g347(.A(new_n769), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n767), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n774), .A2(new_n764), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n760), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n731), .A2(G33), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(new_n468), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT25), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n484), .B2(G139), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(KEYINPUT93), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n783), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n781), .B1(new_n791), .B2(new_n731), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n778), .A2(new_n780), .B1(G2072), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n731), .A2(G26), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT28), .Z(new_n795));
  OR2_X1    g370(.A1(G104), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT92), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G128), .B2(new_n486), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n484), .A2(G140), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n732), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT23), .ZN(new_n805));
  INV_X1    g380(.A(G299), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n732), .ZN(new_n807));
  INV_X1    g382(.A(G1956), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n759), .A2(new_n793), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n746), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n740), .A2(G1961), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n731), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n731), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2090), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT101), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n815), .A2(G2090), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n792), .A2(G2072), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n778), .A2(new_n780), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n743), .A2(new_n811), .A3(new_n812), .A4(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n732), .A2(G23), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n599), .B2(new_n732), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT33), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1976), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT91), .ZN(new_n830));
  MUX2_X1   g405(.A(G6), .B(G305), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT32), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n720), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n732), .A2(G22), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G166), .B2(new_n732), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(G1971), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(G1971), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n825), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  MUX2_X1   g414(.A(G24), .B(G290), .S(G16), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1986), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n731), .A2(G25), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n484), .A2(G131), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n486), .A2(G119), .ZN(new_n844));
  OR2_X1    g419(.A1(G95), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n842), .B1(new_n848), .B2(new_n731), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G1991), .Z(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n841), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n839), .A2(new_n852), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n830), .A2(new_n825), .A3(new_n838), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n823), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n823), .A3(new_n854), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n822), .B1(new_n856), .B2(new_n857), .ZN(G311));
  AND3_X1   g433(.A1(new_n821), .A2(new_n811), .A3(new_n812), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n743), .B(new_n859), .C1(new_n860), .C2(new_n855), .ZN(G150));
  NAND2_X1  g436(.A1(new_n632), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n547), .A2(G55), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n514), .A2(G93), .A3(new_n519), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n867), .A2(new_n506), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n569), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n568), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n864), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  AOI21_X1  g450(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G145));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n882));
  INV_X1    g457(.A(G106), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n468), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n484), .B2(G142), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n486), .A2(KEYINPUT103), .A3(G130), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT103), .B1(new_n486), .B2(G130), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n642), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n642), .B(new_n885), .C1(new_n888), .C2(new_n887), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n848), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n848), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT104), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n791), .B1(new_n771), .B2(new_n776), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n774), .A2(new_n764), .ZN(new_n901));
  INV_X1    g476(.A(new_n790), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n786), .A2(KEYINPUT93), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n904), .B2(new_n783), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n801), .A2(G164), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n799), .A2(new_n503), .A3(new_n800), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n900), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n900), .B2(new_n905), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n896), .B(new_n899), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n898), .B1(new_n897), .B2(new_n893), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n900), .A2(new_n905), .ZN(new_n913));
  INV_X1    g488(.A(new_n908), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n900), .A2(new_n905), .A3(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n651), .B(G160), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G162), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n911), .B2(new_n917), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n881), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n911), .A2(new_n917), .ZN(new_n925));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(KEYINPUT105), .A3(new_n921), .A4(new_n920), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g505(.A(new_n873), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n635), .B(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n615), .A2(G299), .A3(new_n619), .ZN(new_n934));
  AOI21_X1  g509(.A(G299), .B1(new_n615), .B2(new_n619), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n620), .A2(new_n806), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n615), .A2(G299), .A3(new_n619), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n934), .A2(new_n935), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n932), .ZN(new_n944));
  XOR2_X1   g519(.A(G290), .B(G303), .Z(new_n945));
  XOR2_X1   g520(.A(new_n599), .B(G305), .Z(new_n946));
  XNOR2_X1  g521(.A(new_n945), .B(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n944), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n869), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n869), .ZN(G331));
  AND2_X1   g528(.A1(new_n562), .A2(G286), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n592), .B2(G168), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT106), .B1(new_n955), .B2(new_n931), .ZN(new_n956));
  AOI21_X1  g531(.A(G286), .B1(new_n589), .B2(new_n591), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  NOR4_X1   g533(.A1(new_n957), .A2(new_n873), .A3(new_n954), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n592), .A2(G168), .ZN(new_n961));
  INV_X1    g536(.A(new_n954), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n931), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n943), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n931), .A3(new_n962), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n873), .B1(new_n957), .B2(new_n954), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n960), .A2(new_n964), .B1(new_n941), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n947), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n965), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n956), .A2(new_n959), .A3(new_n963), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(new_n940), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n947), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n965), .A2(new_n958), .ZN(new_n978));
  INV_X1    g553(.A(new_n943), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n955), .A2(KEYINPUT106), .A3(new_n931), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n966), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n967), .A2(new_n941), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n969), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n970), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT44), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n970), .A2(new_n974), .A3(new_n976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n969), .A3(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n921), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n989), .B2(new_n983), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n986), .B1(new_n992), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n503), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G125), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n465), .B2(new_n466), .ZN(new_n999));
  INV_X1    g574(.A(new_n477), .ZN(new_n1000));
  OAI21_X1  g575(.A(G2105), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(G40), .A3(new_n472), .A4(new_n469), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1003), .B(G1996), .C1(new_n764), .C2(new_n774), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT108), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n801), .A2(G2067), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n801), .A2(G2067), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1007), .B(new_n1008), .C1(new_n777), .C2(G1996), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n850), .A3(new_n848), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1004), .B1(new_n1011), .B2(new_n1008), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n1004), .B2(G1996), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT125), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n1008), .A2(new_n1007), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n901), .B1(new_n1013), .B2(G1996), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1003), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  XNOR2_X1  g595(.A(new_n847), .B(new_n850), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1004), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1010), .A2(new_n1024), .ZN(new_n1025));
  OR3_X1    g600(.A1(new_n1004), .A2(G1986), .A3(G290), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT48), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n1012), .B(new_n1020), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n806), .A2(KEYINPUT116), .A3(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(KEYINPUT116), .ZN(new_n1034));
  NAND3_X1  g609(.A1(G299), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n996), .A2(G1384), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1002), .B1(new_n503), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT56), .B(G2072), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n997), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n503), .A2(new_n1044), .A3(new_n994), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n503), .B2(new_n994), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1002), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT115), .B1(new_n1047), .B2(G1956), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1002), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n503), .A2(new_n1044), .A3(new_n994), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n808), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1348), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n995), .A2(G2067), .A3(new_n1002), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1056), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1058), .B(new_n1059), .C1(new_n1047), .C2(G1348), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g636(.A1(new_n1038), .A2(new_n1054), .B1(new_n1061), .B2(new_n620), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1036), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1042), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1030), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1030), .A3(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1054), .A2(new_n1064), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1043), .B(new_n1036), .C1(new_n1048), .C2(new_n1053), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n503), .A2(new_n1039), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1002), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n503), .B2(new_n994), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(G1996), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n995), .A2(new_n1002), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT58), .B(G1341), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n569), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT59), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1065), .B(KEYINPUT61), .C1(new_n1054), .C2(new_n1038), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1072), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1061), .A2(KEYINPUT60), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n620), .B1(new_n1061), .B2(KEYINPUT60), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1061), .A2(KEYINPUT60), .A3(new_n620), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1067), .B(new_n1068), .C1(new_n1084), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n520), .B(new_n523), .C1(new_n537), .C2(KEYINPUT72), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n532), .A2(new_n533), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1093), .B(G8), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(G303), .B2(G8), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G8), .ZN(new_n1100));
  INV_X1    g675(.A(G1971), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n1103));
  INV_X1    g678(.A(G2090), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1074), .A4(new_n1050), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1092), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1096), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1110), .B(KEYINPUT113), .C1(new_n1111), .C2(new_n1100), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1102), .A2(KEYINPUT110), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1105), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1102), .A2(KEYINPUT110), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1099), .B(G8), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n597), .A2(new_n598), .A3(G1976), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1118), .B(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(G1976), .B1(new_n597), .B2(new_n598), .ZN(new_n1121));
  OR3_X1    g696(.A1(new_n1121), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n995), .B2(new_n1002), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT112), .B1(new_n1121), .B2(KEYINPUT52), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1120), .A2(new_n1122), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1118), .B(KEYINPUT111), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT52), .B1(new_n1127), .B2(new_n1123), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n720), .B1(new_n604), .B2(new_n605), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n604), .A2(new_n605), .A3(new_n720), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(KEYINPUT49), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT49), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1131), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1129), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1124), .A3(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1126), .A2(new_n1128), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1117), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1091), .B1(new_n1113), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1140), .A2(KEYINPUT123), .A3(new_n1117), .A4(new_n1137), .ZN(new_n1141));
  INV_X1    g716(.A(G1966), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(KEYINPUT114), .B(new_n1142), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1146));
  INV_X1    g721(.A(G2084), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1103), .A2(new_n1147), .A3(new_n1074), .A4(new_n1050), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1145), .A2(G168), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G8), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(G1966), .B1(new_n997), .B2(new_n1040), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1148), .B1(new_n1153), .B2(KEYINPUT114), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1146), .ZN(new_n1155));
  OAI21_X1  g730(.A(G286), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1151), .A2(new_n1100), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT120), .B(G1961), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1051), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(G2078), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1073), .A2(KEYINPUT53), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(new_n1074), .A3(new_n997), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n997), .A2(new_n1040), .A3(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1162), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n592), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n997), .A2(KEYINPUT122), .A3(new_n1074), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1076), .B2(new_n1002), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1164), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n1162), .A3(new_n1168), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1170), .B1(new_n592), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1169), .A2(new_n592), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1175), .B2(G171), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1176), .A2(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND4_X1   g755(.A1(new_n1139), .A2(new_n1141), .A3(new_n1160), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1090), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1170), .B1(new_n1159), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1152), .A2(KEYINPUT62), .A3(new_n1158), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1184), .A2(new_n1139), .A3(new_n1141), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(G288), .A2(G1976), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1136), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1124), .B1(new_n1188), .B2(new_n1134), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1137), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n1117), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1192), .A2(new_n1100), .A3(G286), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1140), .A2(new_n1193), .A3(new_n1117), .A4(new_n1137), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1117), .A2(new_n1137), .ZN(new_n1197));
  OAI21_X1  g772(.A(G8), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1110), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1197), .A2(KEYINPUT63), .A3(new_n1193), .A4(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1191), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1182), .A2(new_n1186), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1003), .A2(G1986), .A3(G290), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1026), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT107), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1025), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1029), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1139), .A2(new_n1160), .A3(new_n1180), .A4(new_n1141), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1088), .ZN(new_n1209));
  OAI22_X1  g784(.A1(new_n1209), .A2(new_n1086), .B1(KEYINPUT60), .B2(new_n1061), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1210), .A2(new_n1083), .A3(new_n1082), .A4(new_n1072), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1068), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1212), .A2(new_n1066), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1208), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1201), .A2(new_n1186), .ZN(new_n1215));
  OAI211_X1 g790(.A(new_n1029), .B(new_n1206), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1028), .B1(new_n1207), .B2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n1220));
  NOR2_X1   g794(.A1(G227), .A2(new_n461), .ZN(new_n1221));
  OAI211_X1 g795(.A(new_n680), .B(new_n1221), .C1(new_n722), .C2(new_n723), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n924), .B2(new_n928), .ZN(new_n1223));
  AND3_X1   g797(.A1(new_n991), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1220), .B1(new_n991), .B2(new_n1223), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n1224), .A2(new_n1225), .ZN(G308));
  NAND2_X1  g800(.A1(new_n991), .A2(new_n1223), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n1227), .A2(KEYINPUT126), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n991), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1229), .ZN(G225));
endmodule


