//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  NAND2_X1  g0006(.A1(G97), .A2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n210), .B(new_n212), .C1(G77), .C2(G244), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(new_n203), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n206), .B(new_n219), .C1(new_n222), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(G250), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  INV_X1    g0038(.A(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n220), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n221), .B1(new_n223), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n221), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT67), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI211_X1 g0064(.A(new_n258), .B(new_n260), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n250), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n253), .B1(G50), .B2(new_n254), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT74), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G223), .A2(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n281), .C1(G77), .C2(new_n274), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n251), .B(G274), .C1(G41), .C2(G45), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n267), .A2(new_n268), .ZN(new_n290));
  INV_X1    g0090(.A(new_n288), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(G190), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n271), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n229), .A2(G1698), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n274), .B(new_n295), .C1(G226), .C2(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n280), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n287), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n284), .A2(new_n209), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR4_X1   g0103(.A1(new_n298), .A2(KEYINPUT13), .A3(new_n299), .A4(new_n300), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n305), .A2(KEYINPUT14), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(G179), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT14), .B1(new_n305), .B2(new_n306), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n262), .A2(G77), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n208), .A2(G20), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n311), .B(new_n312), .C1(new_n259), .C2(new_n256), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(new_n250), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n315));
  OR2_X1    g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n251), .A2(G13), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(G68), .B2(new_n252), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n313), .A2(new_n250), .A3(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n305), .B2(G190), .ZN(new_n324));
  OAI21_X1  g0124(.A(G200), .B1(new_n303), .B2(new_n304), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n288), .A2(KEYINPUT68), .A3(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n288), .A2(new_n306), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT68), .B1(new_n288), .B2(G179), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n328), .A2(new_n267), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n252), .A2(G77), .ZN(new_n332));
  INV_X1    g0132(.A(new_n254), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G20), .A2(G77), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n337), .B1(new_n263), .B2(new_n256), .C1(new_n261), .C2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT70), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n250), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n339), .B2(new_n250), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n332), .B(new_n336), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n250), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n341), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n332), .A4(new_n336), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G238), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n274), .B(new_n351), .C1(new_n229), .C2(G1698), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT69), .B(G107), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(new_n281), .C1(new_n274), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G244), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n354), .B(new_n287), .C1(new_n355), .C2(new_n284), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n345), .A2(new_n350), .B1(new_n306), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(G179), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n294), .A2(new_n327), .A3(new_n331), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n263), .A2(new_n254), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n252), .B2(new_n263), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G58), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n208), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n255), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT76), .ZN(new_n370));
  AND2_X1   g0170(.A1(KEYINPUT3), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n371), .A2(new_n372), .A3(G20), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n370), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n272), .A2(new_n221), .A3(new_n273), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(KEYINPUT76), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n273), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT77), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n371), .A2(new_n372), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT7), .A4(new_n221), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n374), .A2(new_n377), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n369), .B1(new_n383), .B2(G68), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n266), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n375), .A2(new_n376), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT78), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n378), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n373), .A2(KEYINPUT78), .A3(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G68), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n369), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n364), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n280), .A2(G232), .A3(new_n283), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n287), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT80), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT80), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n399), .A3(new_n287), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(G1698), .C1(new_n371), .C2(new_n372), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n274), .A2(KEYINPUT79), .A3(G226), .A4(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n274), .A2(G223), .A3(new_n275), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n281), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n401), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n398), .A2(new_n400), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n281), .B2(new_n408), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n413), .B2(G200), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT17), .B1(new_n395), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n383), .A2(G68), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n394), .A3(new_n250), .ZN(new_n418));
  AND4_X1   g0218(.A1(KEYINPUT17), .A2(new_n418), .A3(new_n363), .A4(new_n414), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n401), .A2(new_n409), .A3(G179), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n413), .B2(new_n306), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n421), .B1(new_n395), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n418), .A2(new_n363), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n356), .A2(G200), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n356), .A2(new_n410), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n345), .A2(new_n350), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n420), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n361), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT5), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G41), .ZN(new_n435));
  INV_X1    g0235(.A(new_n220), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n279), .ZN(new_n437));
  INV_X1    g0237(.A(G41), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n251), .B(G45), .C1(new_n438), .C2(KEYINPUT5), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n434), .A2(G41), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT82), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(G274), .B(new_n437), .C1(new_n441), .C2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT83), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(new_n440), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(KEYINPUT82), .A3(new_n444), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(KEYINPUT83), .A3(new_n437), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G294), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n274), .B1(G257), .B2(new_n275), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G250), .A2(G1698), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n439), .A2(new_n435), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n281), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n458), .A2(new_n281), .B1(new_n460), .B2(G264), .ZN(new_n461));
  INV_X1    g0261(.A(G179), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n454), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n454), .A2(new_n461), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n306), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT92), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT23), .B1(new_n239), .B2(G20), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n239), .A2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G107), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n467), .B1(new_n472), .B2(G20), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT91), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n474), .B(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n466), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n474), .B(KEYINPUT91), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n353), .A2(new_n468), .A3(new_n221), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(KEYINPUT92), .C1(new_n479), .C2(new_n467), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n274), .A2(new_n221), .A3(G87), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n482), .B(KEYINPUT22), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT24), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n481), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n266), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n333), .A2(new_n239), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT25), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n251), .A2(G33), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n254), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n266), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(G107), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n463), .B(new_n465), .C1(new_n488), .C2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n275), .A2(G257), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G264), .A2(G1698), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n274), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n281), .C1(G303), .C2(new_n274), .ZN(new_n502));
  OAI211_X1 g0302(.A(G270), .B(new_n280), .C1(new_n439), .C2(new_n435), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n454), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n241), .A2(G20), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n317), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n507), .B(new_n221), .C1(G33), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n250), .A3(new_n505), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT20), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT89), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n493), .B2(new_n241), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n492), .A2(KEYINPUT89), .A3(new_n266), .A4(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(G169), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n498), .B1(new_n504), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n514), .A2(new_n518), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n504), .A2(G179), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n454), .A2(new_n502), .A3(new_n503), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT21), .A4(G169), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n481), .A2(new_n486), .A3(new_n483), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n486), .B1(new_n481), .B2(new_n483), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n250), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n464), .A2(G200), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n454), .A2(new_n461), .A3(G190), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n495), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n514), .A2(new_n518), .ZN(new_n532));
  INV_X1    g0332(.A(G200), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT90), .B(new_n532), .C1(new_n504), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT90), .ZN(new_n535));
  INV_X1    g0335(.A(new_n503), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n448), .B2(new_n453), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n533), .B1(new_n537), .B2(new_n502), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(new_n521), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n504), .A2(G190), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n497), .A2(new_n525), .A3(new_n531), .A4(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n280), .B(G250), .C1(G1), .C2(new_n442), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n355), .A2(G1698), .ZN(new_n545));
  OAI221_X1 g0345(.A(new_n545), .B1(G238), .B2(G1698), .C1(new_n371), .C2(new_n372), .ZN(new_n546));
  INV_X1    g0346(.A(G33), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n241), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n548), .B2(new_n281), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n443), .A2(G274), .ZN(new_n550));
  XOR2_X1   g0350(.A(new_n550), .B(KEYINPUT86), .Z(new_n551));
  AND2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT87), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(G190), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n551), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT87), .B1(new_n555), .B2(new_n410), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT88), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n554), .B2(new_n556), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n552), .A2(new_n533), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n297), .A2(new_n221), .ZN(new_n562));
  INV_X1    g0362(.A(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n508), .ZN(new_n564));
  OAI211_X1 g0364(.A(KEYINPUT19), .B(new_n562), .C1(new_n353), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n274), .A2(new_n221), .A3(G68), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n297), .A2(G20), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n566), .C1(KEYINPUT19), .C2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n250), .B1(new_n333), .B2(new_n338), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n563), .B2(new_n493), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n558), .A2(new_n560), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n542), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT81), .ZN(new_n574));
  AND2_X1   g0374(.A1(G250), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n274), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n371), .C2(new_n372), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n507), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(new_n275), .C1(new_n371), .C2(new_n372), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n281), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(new_n280), .C1(new_n439), .C2(new_n435), .ZN(new_n586));
  AND4_X1   g0386(.A1(KEYINPUT85), .A2(new_n454), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n586), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n448), .B2(new_n453), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT85), .B1(new_n589), .B2(new_n585), .ZN(new_n590));
  OAI21_X1  g0390(.A(G190), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n493), .A2(new_n508), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n254), .A2(G97), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n388), .A2(new_n353), .A3(new_n389), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n239), .A2(KEYINPUT6), .A3(G97), .ZN(new_n595));
  XOR2_X1   g0395(.A(G97), .B(G107), .Z(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(KEYINPUT6), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI211_X1 g0399(.A(new_n592), .B(new_n593), .C1(new_n599), .C2(new_n250), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n454), .A2(new_n585), .A3(new_n586), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G200), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT84), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n604), .A3(G200), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n591), .A2(new_n600), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n600), .ZN(new_n608));
  INV_X1    g0408(.A(new_n601), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n462), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n589), .A2(KEYINPUT85), .A3(new_n585), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n608), .B(new_n610), .C1(new_n614), .C2(G169), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n493), .A2(new_n338), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n569), .A2(new_n618), .B1(new_n555), .B2(new_n306), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n552), .A2(new_n462), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n433), .A2(new_n573), .A3(new_n617), .A4(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n572), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(KEYINPUT26), .A3(new_n616), .ZN(new_n624));
  INV_X1    g0424(.A(new_n571), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n557), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n465), .A2(new_n463), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n528), .B2(new_n495), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n606), .B(new_n531), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n631), .B2(new_n615), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n624), .B1(new_n632), .B2(KEYINPUT26), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n621), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n433), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT93), .ZN(new_n636));
  INV_X1    g0436(.A(new_n331), .ZN(new_n637));
  INV_X1    g0437(.A(new_n360), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n326), .A2(new_n638), .B1(new_n322), .B2(new_n310), .ZN(new_n639));
  INV_X1    g0439(.A(new_n420), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n428), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n637), .B1(new_n641), .B2(new_n294), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n636), .A2(new_n642), .ZN(G369));
  NAND3_X1  g0443(.A1(new_n251), .A2(new_n221), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G343), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT94), .Z(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n532), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT95), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n525), .A3(new_n541), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n525), .B2(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n497), .A2(new_n531), .ZN(new_n656));
  INV_X1    g0456(.A(new_n649), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n488), .B2(new_n496), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n497), .B2(new_n649), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n531), .B1(new_n629), .B2(new_n630), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(new_n657), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n204), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n353), .A2(G116), .A3(new_n564), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n225), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n634), .A2(new_n649), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT29), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n572), .A2(KEYINPUT26), .A3(new_n615), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n627), .A2(KEYINPUT26), .B1(new_n620), .B2(new_n619), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n615), .B1(new_n662), .B2(new_n607), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT26), .B1(new_n677), .B2(new_n626), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n675), .B(new_n676), .C1(new_n678), .C2(new_n616), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n649), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n674), .B1(new_n673), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n587), .A2(new_n590), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n504), .A2(G179), .A3(new_n461), .A4(new_n552), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n461), .A2(new_n549), .A3(new_n551), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n523), .A2(new_n686), .A3(new_n462), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n614), .A2(new_n687), .A3(KEYINPUT30), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n523), .A2(new_n464), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n462), .A3(new_n555), .A4(new_n601), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT31), .B1(new_n691), .B2(new_n657), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT96), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n657), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT96), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n573), .A2(new_n617), .A3(new_n621), .A4(new_n649), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n702), .A2(KEYINPUT97), .A3(G330), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT97), .B1(new_n702), .B2(G330), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n671), .B1(new_n707), .B2(G1), .ZN(G364));
  NOR2_X1   g0508(.A1(G13), .A2(G33), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n653), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n226), .A2(new_n442), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n665), .A2(new_n274), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n714), .B(new_n715), .C1(new_n247), .C2(new_n442), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n665), .A2(new_n380), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT99), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G355), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n716), .B(new_n719), .C1(G116), .C2(new_n204), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT100), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n220), .B1(G20), .B2(new_n306), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G13), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(new_n442), .A3(G20), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n666), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n533), .A2(G179), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(G20), .A3(G190), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n274), .B1(new_n732), .B2(new_n563), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT101), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n508), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n221), .A2(new_n462), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n410), .A3(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n739), .B1(G58), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n741), .A2(new_n533), .A3(G190), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G68), .A2(new_n744), .B1(new_n745), .B2(G77), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n221), .A2(G190), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n735), .ZN(new_n748));
  INV_X1    g0548(.A(G159), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT32), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G50), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n743), .A2(new_n746), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n731), .A2(new_n747), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n734), .B(new_n755), .C1(G107), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n752), .B(KEYINPUT102), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT103), .B(G326), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n737), .A2(G294), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n732), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G303), .ZN(new_n766));
  INV_X1    g0566(.A(new_n748), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n274), .B1(new_n767), .B2(G329), .ZN(new_n768));
  AND4_X1   g0568(.A1(new_n762), .A2(new_n764), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(G283), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G311), .A2(new_n745), .B1(new_n742), .B2(G322), .ZN(new_n771));
  AND4_X1   g0571(.A1(new_n761), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n722), .B1(new_n758), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n713), .A2(new_n724), .A3(new_n730), .A4(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n653), .A2(G330), .ZN(new_n775));
  INV_X1    g0575(.A(new_n730), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(new_n654), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n777), .ZN(G396));
  NAND2_X1  g0578(.A1(new_n638), .A2(new_n649), .ZN(new_n779));
  INV_X1    g0579(.A(new_n431), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n649), .B1(new_n345), .B2(new_n350), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n360), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n705), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n783), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n703), .B2(new_n704), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n672), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n657), .B1(new_n633), .B2(new_n621), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n784), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(new_n776), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G132), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n274), .B1(new_n748), .B2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G143), .A2(new_n742), .B1(new_n745), .B2(G159), .ZN(new_n794));
  INV_X1    g0594(.A(G137), .ZN(new_n795));
  INV_X1    g0595(.A(new_n744), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n752), .C1(new_n257), .C2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G50), .B2(new_n765), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n757), .A2(G68), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n793), .B(new_n801), .C1(G58), .C2(new_n737), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n745), .A2(G116), .B1(G87), .B2(new_n757), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n239), .B2(new_n732), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G303), .B2(new_n753), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n274), .B(new_n739), .C1(G311), .C2(new_n767), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  INV_X1    g0607(.A(new_n742), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G283), .B2(new_n744), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n722), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n722), .A2(new_n709), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n334), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n783), .A2(new_n709), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n811), .A2(new_n730), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n791), .A2(new_n815), .ZN(G384));
  AOI21_X1  g0616(.A(new_n241), .B1(new_n597), .B2(KEYINPUT35), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n222), .C1(KEYINPUT35), .C2(new_n597), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT36), .ZN(new_n819));
  OAI21_X1  g0619(.A(G77), .B1(new_n365), .B2(new_n208), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n225), .A2(new_n820), .B1(G50), .B2(new_n208), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n821), .A2(G1), .A3(new_n725), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n692), .A2(new_n693), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n701), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n322), .A2(new_n657), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n323), .A2(new_n326), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n310), .A2(new_n825), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n783), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n824), .A2(KEYINPUT40), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT105), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n415), .B2(new_n419), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n418), .A2(new_n414), .A3(new_n363), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT17), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n395), .A2(KEYINPUT17), .A3(new_n414), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT105), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n832), .A2(new_n428), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n647), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n395), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n426), .B1(new_n423), .B2(new_n647), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n833), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n833), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT37), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n838), .A2(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT106), .B1(new_n846), .B2(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n837), .A2(new_n428), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT105), .B1(new_n835), .B2(new_n836), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n845), .A2(new_n843), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT106), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n384), .A2(KEYINPUT16), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n364), .B1(new_n858), .B2(new_n385), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n859), .B2(new_n839), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n417), .A2(new_n250), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n363), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(KEYINPUT104), .A3(new_n647), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n423), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n860), .A2(new_n863), .A3(new_n833), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n843), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n420), .A2(new_n428), .B1(new_n860), .B2(new_n863), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n847), .A2(new_n855), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n830), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n841), .A2(new_n842), .A3(new_n833), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n854), .B1(new_n875), .B2(new_n868), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n606), .A2(new_n615), .A3(new_n621), .ZN(new_n878));
  NOR4_X1   g0678(.A1(new_n542), .A2(new_n878), .A3(new_n572), .A4(new_n657), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n697), .A2(new_n699), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n829), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n873), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n872), .A2(new_n882), .A3(G330), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n433), .A2(G330), .A3(new_n824), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT107), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n872), .A2(new_n882), .A3(new_n433), .A4(new_n824), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n428), .A2(new_n647), .ZN(new_n889));
  INV_X1    g0689(.A(new_n827), .ZN(new_n890));
  INV_X1    g0690(.A(new_n828), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n634), .A2(new_n649), .A3(new_n782), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n779), .ZN(new_n894));
  INV_X1    g0694(.A(new_n877), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n870), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n871), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n323), .A2(new_n657), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n888), .B(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n674), .B(new_n433), .C1(new_n673), .C2(new_n680), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n642), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n251), .B1(G13), .B2(new_n221), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n819), .B(new_n822), .C1(new_n906), .C2(new_n907), .ZN(G367));
  AOI22_X1  g0708(.A1(new_n767), .A2(G317), .B1(new_n737), .B2(new_n353), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n910));
  INV_X1    g0710(.A(G303), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n909), .B(new_n910), .C1(new_n808), .C2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT46), .B1(new_n765), .B2(G116), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n796), .A2(new_n807), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n745), .A2(G283), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n757), .A2(G97), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n915), .A2(new_n380), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(G311), .B2(new_n759), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT111), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n767), .A2(G137), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n738), .A2(new_n208), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n759), .B2(G143), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n257), .B2(new_n808), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n274), .B1(new_n732), .B2(new_n365), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n757), .A2(G77), .ZN(new_n926));
  INV_X1    g0726(.A(new_n745), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n926), .B1(new_n927), .B2(new_n259), .C1(new_n749), .C2(new_n796), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n920), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT47), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n722), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n657), .A2(new_n570), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n621), .B1(new_n627), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n621), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n711), .ZN(new_n937));
  INV_X1    g0737(.A(new_n715), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n723), .B1(new_n204), .B2(new_n338), .C1(new_n236), .C2(new_n938), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n932), .A2(new_n730), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n525), .A2(new_n657), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n656), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n606), .B(new_n615), .C1(new_n600), .C2(new_n649), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT42), .Z(new_n945));
  OR2_X1    g0745(.A1(new_n943), .A2(new_n497), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n657), .B1(new_n946), .B2(new_n615), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT43), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n945), .A2(new_n947), .B1(new_n948), .B2(new_n936), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n936), .A2(new_n948), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n661), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n943), .B1(new_n615), .B2(new_n649), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n951), .B(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n663), .A2(new_n617), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT44), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(KEYINPUT110), .A3(new_n958), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n956), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n953), .A2(new_n663), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n952), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n959), .A2(new_n661), .A3(new_n960), .A4(new_n963), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n942), .B1(new_n660), .B2(new_n941), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n654), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n707), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n666), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n729), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n940), .B1(new_n955), .B2(new_n973), .ZN(G387));
  INV_X1    g0774(.A(new_n969), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n707), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n706), .A2(new_n969), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n666), .B(KEYINPUT116), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n975), .A2(new_n729), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT112), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n927), .A2(new_n208), .B1(new_n732), .B2(new_n334), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n380), .B(new_n983), .C1(G150), .C2(new_n767), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n744), .A2(new_n264), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n808), .A2(new_n259), .B1(new_n749), .B2(new_n752), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n738), .A2(new_n338), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n917), .A3(new_n985), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n759), .A2(G322), .B1(G311), .B2(new_n744), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT115), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G303), .A2(new_n745), .B1(new_n742), .B2(G317), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  INV_X1    g0794(.A(G283), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n994), .B1(new_n995), .B2(new_n738), .C1(new_n807), .C2(new_n732), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT49), .Z(new_n997));
  INV_X1    g0797(.A(new_n760), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n380), .B1(new_n756), .B2(new_n241), .C1(new_n998), .C2(new_n748), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n989), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n722), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n938), .B1(new_n232), .B2(G45), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n208), .A2(new_n334), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n263), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT50), .B1(new_n263), .B2(G50), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1004), .A2(new_n442), .A3(new_n668), .A4(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n668), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n718), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1007), .B(new_n1009), .C1(G107), .C2(new_n204), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT113), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n723), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n730), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1001), .B(new_n1016), .C1(new_n660), .C2(new_n712), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n980), .A2(new_n982), .A3(new_n1017), .ZN(G393));
  NAND3_X1  g0818(.A1(new_n965), .A2(new_n729), .A3(new_n966), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n953), .A2(new_n712), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n742), .A2(G311), .B1(new_n753), .B2(G317), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n274), .B(new_n1022), .C1(G294), .C2(new_n745), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n911), .B2(new_n796), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n767), .A2(G322), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n732), .A2(new_n995), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n738), .A2(new_n241), .B1(new_n756), .B2(new_n239), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n742), .A2(G159), .B1(new_n753), .B2(G150), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT117), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n745), .A2(new_n264), .B1(G68), .B2(new_n765), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n334), .B2(new_n738), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n380), .B1(new_n767), .B2(G143), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n563), .B2(new_n756), .C1(new_n796), .C2(new_n259), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n722), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n723), .B1(new_n508), .B2(new_n204), .C1(new_n243), .C2(new_n938), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1020), .A2(new_n730), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n976), .A2(new_n967), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n979), .B1(new_n976), .B2(new_n967), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1019), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(G390));
  INV_X1    g0842(.A(new_n892), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n785), .B(new_n1043), .C1(new_n703), .C2(new_n704), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n679), .A2(new_n649), .A3(new_n782), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n779), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(G330), .B(new_n785), .C1(new_n880), .C2(new_n879), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT118), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n892), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n892), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT118), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1044), .A2(new_n1047), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n824), .A2(G330), .A3(new_n829), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n786), .B2(new_n892), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n779), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n789), .B2(new_n782), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n904), .A2(new_n642), .A3(new_n884), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n782), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n657), .B(new_n1063), .C1(new_n633), .C2(new_n621), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1043), .B1(new_n1064), .B2(new_n1057), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n900), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n871), .A2(new_n898), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n897), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1065), .A2(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n871), .A2(new_n1066), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1055), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1066), .B1(new_n1058), .B2(new_n892), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1046), .A2(new_n1043), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1070), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1075), .A2(new_n1078), .A3(new_n1044), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1062), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT119), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1059), .A2(new_n1079), .A3(new_n1072), .A4(new_n1061), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT119), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1062), .A2(new_n1084), .A3(new_n1080), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n979), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n800), .B1(new_n563), .B2(new_n732), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n744), .A2(new_n353), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n808), .B2(new_n241), .C1(new_n508), .C2(new_n927), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(G77), .C2(new_n737), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n274), .B1(new_n767), .B2(G294), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n995), .C2(new_n752), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g0893(.A(G128), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n752), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n738), .A2(new_n749), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  AOI21_X1  g0897(.A(new_n380), .B1(new_n745), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n259), .B2(new_n756), .C1(new_n792), .C2(new_n808), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(G137), .C2(new_n744), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n732), .A2(new_n257), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n767), .A2(G125), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1093), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n776), .B1(new_n1105), .B2(new_n722), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n812), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n264), .B2(new_n1107), .C1(new_n899), .C2(new_n710), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT121), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1072), .A2(new_n1079), .A3(new_n729), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1086), .A2(new_n1109), .A3(new_n1110), .ZN(G378));
  NAND2_X1  g0911(.A1(new_n294), .A2(new_n331), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n267), .A2(new_n647), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n709), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n259), .B1(new_n371), .B2(G41), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1097), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n732), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n927), .A2(new_n795), .B1(new_n808), .B2(new_n1094), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(G125), .C2(new_n753), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n792), .B2(new_n796), .C1(new_n257), .C2(new_n738), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n757), .A2(G159), .ZN(new_n1125));
  AOI21_X1  g0925(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n547), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1123), .A2(KEYINPUT59), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1118), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n922), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n334), .B2(new_n732), .C1(new_n338), .C2(new_n927), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n380), .B1(new_n796), .B2(new_n508), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n438), .B1(new_n752), .B2(new_n241), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n756), .A2(new_n365), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n239), .B2(new_n808), .C1(new_n995), .C2(new_n748), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT58), .Z(new_n1137));
  OAI21_X1  g0937(.A(new_n722), .B1(new_n1129), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n812), .A2(new_n259), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1117), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n730), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1114), .B(new_n1115), .Z(new_n1142));
  INV_X1    g0942(.A(new_n883), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(KEYINPUT122), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n872), .A2(new_n882), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n896), .A2(new_n1145), .A3(new_n901), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n896), .B2(new_n901), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1065), .A2(new_n877), .B1(new_n428), .B2(new_n647), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1066), .B(new_n897), .C1(new_n871), .C2(new_n898), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1143), .B(KEYINPUT122), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n896), .A2(new_n901), .A3(new_n1145), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT122), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1116), .B1(new_n883), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n729), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1141), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n702), .A2(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT97), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n702), .A2(KEYINPUT97), .A3(G330), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n783), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1054), .B1(new_n1164), .B2(new_n1043), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1058), .ZN(new_n1166));
  AND4_X1   g0966(.A1(new_n779), .A2(new_n1052), .A3(new_n1045), .A4(new_n1050), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1165), .A2(new_n1166), .B1(new_n1167), .B2(new_n1044), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1061), .B1(new_n1080), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1169), .A2(KEYINPUT57), .A3(new_n1155), .A4(new_n1148), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n979), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1169), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1159), .B1(new_n1171), .B2(new_n1173), .ZN(G375));
  NAND2_X1  g0974(.A1(new_n892), .A2(new_n709), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n745), .A2(new_n353), .B1(G97), .B2(new_n765), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1176), .A2(new_n926), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n241), .B2(new_n796), .C1(new_n995), .C2(new_n808), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n752), .A2(new_n807), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n380), .B1(new_n748), .B2(new_n911), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1178), .A2(new_n987), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n753), .A2(G132), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT124), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n1094), .B2(new_n748), .C1(new_n795), .C2(new_n808), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n732), .A2(new_n749), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n927), .A2(new_n257), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n380), .B(new_n1134), .C1(G50), .C2(new_n737), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n796), .B2(new_n1119), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n722), .B1(new_n1181), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n730), .B1(G68), .B2(new_n1107), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT123), .Z(new_n1192));
  NAND3_X1  g0992(.A1(new_n1175), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1168), .B2(new_n1157), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1053), .B(new_n1060), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1062), .A2(new_n972), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(G381));
  NOR2_X1   g0998(.A1(G375), .A2(G378), .ZN(new_n1199));
  INV_X1    g0999(.A(G384), .ZN(new_n1200));
  INV_X1    g1000(.A(G381), .ZN(new_n1201));
  INV_X1    g1001(.A(G396), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n980), .A2(new_n1202), .A3(new_n982), .A4(new_n1017), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(G387), .A2(G390), .A3(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1204), .ZN(G407));
  INV_X1    g1005(.A(new_n1199), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G407), .B(G213), .C1(G343), .C2(new_n1206), .ZN(G409));
  INV_X1    g1007(.A(KEYINPUT126), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(G387), .B2(G390), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1203), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1211), .A3(new_n1203), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1210), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1216), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1215), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1213), .A2(new_n1218), .B1(new_n1219), .B2(new_n1209), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(G213), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(G343), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G375), .B2(G378), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n979), .B1(new_n1196), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n1196), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1200), .B1(new_n1229), .B2(new_n1194), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1060), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1226), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1196), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n979), .B(new_n1231), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(G384), .A3(new_n1195), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1156), .B1(new_n1061), .B2(new_n1083), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1158), .B1(new_n1238), .B2(new_n972), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1239), .A2(new_n1109), .A3(new_n1110), .A4(new_n1086), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1224), .A2(new_n1225), .A3(new_n1237), .A4(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G375), .A2(G378), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1223), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1244), .A2(new_n1240), .A3(new_n1237), .A4(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1240), .A3(new_n1245), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1223), .A2(G2897), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1230), .A2(new_n1235), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1246), .A2(KEYINPUT62), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1221), .B1(new_n1243), .B2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1224), .A2(KEYINPUT63), .A3(new_n1237), .A4(new_n1240), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT61), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT63), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1258), .B2(new_n1246), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1261), .A2(new_n1257), .A3(new_n1242), .A4(new_n1241), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1221), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1246), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1255), .B(new_n1254), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n1265), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1260), .A2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(new_n1206), .A2(new_n1244), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(new_n1237), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(new_n1221), .ZN(G402));
endmodule


