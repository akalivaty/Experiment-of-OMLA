

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n432), .B(n431), .ZN(n433) );
  AND2_X1 U324 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U325 ( .A(G29GAT), .B(G43GAT), .Z(n292) );
  XOR2_X1 U326 ( .A(KEYINPUT120), .B(n558), .Z(n293) );
  XOR2_X1 U327 ( .A(KEYINPUT118), .B(n552), .Z(n294) );
  XNOR2_X1 U328 ( .A(n502), .B(KEYINPUT45), .ZN(n503) );
  NOR2_X1 U329 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U330 ( .A(n430), .B(n291), .ZN(n431) );
  XNOR2_X1 U331 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n546) );
  XNOR2_X1 U332 ( .A(n547), .B(n546), .ZN(n566) );
  XNOR2_X1 U333 ( .A(n442), .B(n441), .ZN(n562) );
  XNOR2_X1 U334 ( .A(KEYINPUT82), .B(KEYINPUT0), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n295), .B(KEYINPUT81), .ZN(n358) );
  XNOR2_X1 U336 ( .A(n358), .B(KEYINPUT91), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n296), .B(KEYINPUT4), .ZN(n316) );
  XOR2_X1 U338 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n298) );
  XNOR2_X1 U339 ( .A(G141GAT), .B(G57GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U341 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n300) );
  XNOR2_X1 U342 ( .A(KEYINPUT88), .B(KEYINPUT5), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(n302), .B(n301), .Z(n314) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT75), .Z(n425) );
  XNOR2_X1 U346 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n303), .B(KEYINPUT2), .ZN(n386) );
  XOR2_X1 U348 ( .A(n425), .B(n386), .Z(n305) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n312) );
  XOR2_X1 U351 ( .A(G148GAT), .B(G162GAT), .Z(n307) );
  XNOR2_X1 U352 ( .A(G127GAT), .B(G120GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U354 ( .A(n308), .B(G85GAT), .Z(n310) );
  XOR2_X1 U355 ( .A(G113GAT), .B(G1GAT), .Z(n328) );
  XNOR2_X1 U356 ( .A(n328), .B(G29GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U360 ( .A(n316), .B(n315), .Z(n565) );
  XNOR2_X1 U361 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n317) );
  XNOR2_X1 U362 ( .A(n292), .B(n317), .ZN(n432) );
  XOR2_X1 U363 ( .A(G141GAT), .B(G22GAT), .Z(n391) );
  XNOR2_X1 U364 ( .A(n432), .B(n391), .ZN(n318) );
  XOR2_X1 U365 ( .A(G169GAT), .B(G8GAT), .Z(n367) );
  XNOR2_X1 U366 ( .A(n318), .B(n367), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n320) );
  NAND2_X1 U368 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U370 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n324) );
  XNOR2_X1 U372 ( .A(G15GAT), .B(G197GAT), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n325), .B(KEYINPUT30), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U376 ( .A(n329), .B(n328), .Z(n331) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G50GAT), .ZN(n330) );
  XOR2_X1 U378 ( .A(n331), .B(n330), .Z(n475) );
  INV_X1 U379 ( .A(n475), .ZN(n569) );
  XOR2_X1 U380 ( .A(G120GAT), .B(G71GAT), .Z(n348) );
  XOR2_X1 U381 ( .A(G78GAT), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n379) );
  XOR2_X1 U384 ( .A(G64GAT), .B(G92GAT), .Z(n335) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n370) );
  XNOR2_X1 U387 ( .A(n379), .B(n370), .ZN(n340) );
  XOR2_X1 U388 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n337) );
  NAND2_X1 U389 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n338), .B(KEYINPUT71), .Z(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U393 ( .A(KEYINPUT33), .B(n341), .Z(n343) );
  XOR2_X1 U394 ( .A(KEYINPUT13), .B(G57GAT), .Z(n410) );
  XNOR2_X1 U395 ( .A(n410), .B(KEYINPUT72), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n348), .B(n344), .ZN(n345) );
  XOR2_X1 U398 ( .A(G99GAT), .B(G85GAT), .Z(n426) );
  XNOR2_X1 U399 ( .A(n345), .B(n426), .ZN(n573) );
  INV_X1 U400 ( .A(n573), .ZN(n505) );
  NOR2_X1 U401 ( .A1(n569), .A2(n505), .ZN(n460) );
  XOR2_X1 U402 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n347) );
  XNOR2_X1 U403 ( .A(KEYINPUT65), .B(KEYINPUT83), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n366) );
  XOR2_X1 U405 ( .A(G190GAT), .B(n348), .Z(n350) );
  XOR2_X1 U406 ( .A(G15GAT), .B(G127GAT), .Z(n418) );
  XNOR2_X1 U407 ( .A(G43GAT), .B(n418), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n362) );
  XOR2_X1 U409 ( .A(G176GAT), .B(G99GAT), .Z(n352) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(G134GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U412 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n354) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U415 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n357), .B(KEYINPUT18), .ZN(n374) );
  XNOR2_X1 U418 ( .A(n358), .B(n374), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U421 ( .A1(G227GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n492) );
  XOR2_X1 U424 ( .A(G36GAT), .B(G190GAT), .Z(n430) );
  XNOR2_X1 U425 ( .A(n367), .B(n430), .ZN(n378) );
  XOR2_X1 U426 ( .A(G183GAT), .B(KEYINPUT77), .Z(n411) );
  XOR2_X1 U427 ( .A(KEYINPUT92), .B(n411), .Z(n369) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U431 ( .A(G211GAT), .B(KEYINPUT21), .Z(n373) );
  XNOR2_X1 U432 ( .A(G197GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n374), .B(n387), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U436 ( .A(n378), .B(n377), .Z(n543) );
  XNOR2_X1 U437 ( .A(n543), .B(KEYINPUT27), .ZN(n512) );
  XOR2_X1 U438 ( .A(n379), .B(G204GAT), .Z(n381) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U441 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n383) );
  XNOR2_X1 U442 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U444 ( .A(n385), .B(n384), .Z(n389) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U448 ( .A(G50GAT), .B(G162GAT), .ZN(n438) );
  XNOR2_X1 U449 ( .A(n392), .B(n438), .ZN(n542) );
  XNOR2_X1 U450 ( .A(KEYINPUT28), .B(n542), .ZN(n514) );
  INV_X1 U451 ( .A(n514), .ZN(n471) );
  NOR2_X1 U452 ( .A1(n512), .A2(n471), .ZN(n393) );
  NAND2_X1 U453 ( .A1(n492), .A2(n393), .ZN(n394) );
  INV_X1 U454 ( .A(n565), .ZN(n510) );
  NAND2_X1 U455 ( .A1(n394), .A2(n510), .ZN(n403) );
  INV_X1 U456 ( .A(n492), .ZN(n550) );
  INV_X1 U457 ( .A(n543), .ZN(n466) );
  NAND2_X1 U458 ( .A1(n550), .A2(n466), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n542), .A2(n395), .ZN(n396) );
  XOR2_X1 U460 ( .A(KEYINPUT25), .B(n396), .Z(n401) );
  NOR2_X1 U461 ( .A1(n550), .A2(n542), .ZN(n397) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(n397), .Z(n398) );
  XOR2_X1 U463 ( .A(KEYINPUT26), .B(n398), .Z(n528) );
  NOR2_X1 U464 ( .A1(n528), .A2(n512), .ZN(n399) );
  NOR2_X1 U465 ( .A1(n510), .A2(n399), .ZN(n400) );
  NAND2_X1 U466 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U467 ( .A1(n403), .A2(n402), .ZN(n457) );
  XOR2_X1 U468 ( .A(G155GAT), .B(G211GAT), .Z(n405) );
  XNOR2_X1 U469 ( .A(G22GAT), .B(G8GAT), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U471 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n407) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G64GAT), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n422) );
  XOR2_X1 U475 ( .A(n411), .B(n410), .Z(n413) );
  XNOR2_X1 U476 ( .A(G71GAT), .B(G78GAT), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U478 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n415) );
  NAND2_X1 U479 ( .A1(G231GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U481 ( .A(n417), .B(n416), .Z(n420) );
  XNOR2_X1 U482 ( .A(n418), .B(KEYINPUT12), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n578) );
  XOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n424) );
  XNOR2_X1 U486 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n423) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n442) );
  XOR2_X1 U488 ( .A(KEYINPUT74), .B(n425), .Z(n429) );
  INV_X1 U489 ( .A(n426), .ZN(n427) );
  XOR2_X1 U490 ( .A(G218GAT), .B(n427), .Z(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U492 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n436) );
  XNOR2_X1 U494 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U496 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n441) );
  INV_X1 U498 ( .A(n562), .ZN(n443) );
  NOR2_X1 U499 ( .A1(n578), .A2(n443), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT80), .B(n444), .Z(n445) );
  XNOR2_X1 U501 ( .A(n445), .B(KEYINPUT16), .ZN(n446) );
  NOR2_X1 U502 ( .A1(n457), .A2(n446), .ZN(n477) );
  NAND2_X1 U503 ( .A1(n460), .A2(n477), .ZN(n454) );
  NOR2_X1 U504 ( .A1(n565), .A2(n454), .ZN(n448) );
  XNOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U507 ( .A(G1GAT), .B(n449), .Z(G1324GAT) );
  NOR2_X1 U508 ( .A1(n543), .A2(n454), .ZN(n451) );
  XNOR2_X1 U509 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(G1325GAT) );
  NOR2_X1 U511 ( .A1(n492), .A2(n454), .ZN(n453) );
  XNOR2_X1 U512 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(G1326GAT) );
  NOR2_X1 U514 ( .A1(n514), .A2(n454), .ZN(n455) );
  XOR2_X1 U515 ( .A(G22GAT), .B(n455), .Z(G1327GAT) );
  XNOR2_X1 U516 ( .A(KEYINPUT36), .B(KEYINPUT97), .ZN(n456) );
  XOR2_X1 U517 ( .A(n456), .B(n562), .Z(n584) );
  NOR2_X1 U518 ( .A1(n584), .A2(n457), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n578), .A2(n458), .ZN(n459) );
  XNOR2_X1 U520 ( .A(KEYINPUT37), .B(n459), .ZN(n488) );
  NAND2_X1 U521 ( .A1(n488), .A2(n460), .ZN(n461) );
  XOR2_X1 U522 ( .A(KEYINPUT38), .B(n461), .Z(n472) );
  NAND2_X1 U523 ( .A1(n472), .A2(n510), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n463) );
  XNOR2_X1 U525 ( .A(G29GAT), .B(KEYINPUT98), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(G1328GAT) );
  NAND2_X1 U528 ( .A1(n472), .A2(n466), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n467), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n469) );
  NAND2_X1 U531 ( .A1(n550), .A2(n472), .ZN(n468) );
  XNOR2_X1 U532 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U533 ( .A(G43GAT), .B(n470), .ZN(G1330GAT) );
  NAND2_X1 U534 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n473), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U536 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n474) );
  XOR2_X1 U537 ( .A(n474), .B(n573), .Z(n553) );
  NOR2_X1 U538 ( .A1(n553), .A2(n475), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(KEYINPUT100), .ZN(n487) );
  NAND2_X1 U540 ( .A1(n477), .A2(n487), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n565), .A2(n483), .ZN(n478) );
  XOR2_X1 U542 ( .A(G57GAT), .B(n478), .Z(n479) );
  XNOR2_X1 U543 ( .A(KEYINPUT42), .B(n479), .ZN(G1332GAT) );
  NOR2_X1 U544 ( .A1(n543), .A2(n483), .ZN(n481) );
  XNOR2_X1 U545 ( .A(G64GAT), .B(KEYINPUT101), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(G1333GAT) );
  NOR2_X1 U547 ( .A1(n492), .A2(n483), .ZN(n482) );
  XOR2_X1 U548 ( .A(G71GAT), .B(n482), .Z(G1334GAT) );
  NOR2_X1 U549 ( .A1(n514), .A2(n483), .ZN(n485) );
  XNOR2_X1 U550 ( .A(KEYINPUT43), .B(KEYINPUT102), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U552 ( .A(G78GAT), .B(n486), .ZN(G1335GAT) );
  NAND2_X1 U553 ( .A1(n488), .A2(n487), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n565), .A2(n494), .ZN(n489) );
  XOR2_X1 U555 ( .A(G85GAT), .B(n489), .Z(G1336GAT) );
  NOR2_X1 U556 ( .A1(n543), .A2(n494), .ZN(n491) );
  XNOR2_X1 U557 ( .A(G92GAT), .B(KEYINPUT103), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n491), .B(n490), .ZN(G1337GAT) );
  NOR2_X1 U559 ( .A1(n492), .A2(n494), .ZN(n493) );
  XOR2_X1 U560 ( .A(G99GAT), .B(n493), .Z(G1338GAT) );
  NOR2_X1 U561 ( .A1(n514), .A2(n494), .ZN(n496) );
  XNOR2_X1 U562 ( .A(KEYINPUT44), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U564 ( .A(G106GAT), .B(n497), .Z(G1339GAT) );
  NAND2_X1 U565 ( .A1(n562), .A2(n578), .ZN(n500) );
  NOR2_X1 U566 ( .A1(n569), .A2(n553), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n498), .B(KEYINPUT46), .ZN(n499) );
  NOR2_X1 U568 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n501), .B(KEYINPUT47), .ZN(n508) );
  NOR2_X1 U570 ( .A1(n578), .A2(n584), .ZN(n502) );
  NAND2_X1 U571 ( .A1(n503), .A2(n569), .ZN(n504) );
  XNOR2_X1 U572 ( .A(KEYINPUT105), .B(n506), .ZN(n507) );
  NAND2_X1 U573 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(KEYINPUT48), .ZN(n544) );
  NAND2_X1 U575 ( .A1(n544), .A2(n510), .ZN(n511) );
  NOR2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT106), .B(n513), .ZN(n529) );
  AND2_X1 U578 ( .A1(n529), .A2(n514), .ZN(n515) );
  NAND2_X1 U579 ( .A1(n550), .A2(n515), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n569), .A2(n523), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G113GAT), .B(KEYINPUT107), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1340GAT) );
  NOR2_X1 U583 ( .A1(n553), .A2(n523), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT49), .B(KEYINPUT108), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G120GAT), .B(n520), .ZN(G1341GAT) );
  NOR2_X1 U587 ( .A1(n578), .A2(n523), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT50), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G127GAT), .B(n522), .ZN(G1342GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n562), .ZN(n527) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(KEYINPUT51), .Z(n525) );
  XNOR2_X1 U592 ( .A(G134GAT), .B(KEYINPUT109), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1343GAT) );
  INV_X1 U595 ( .A(n528), .ZN(n567) );
  NAND2_X1 U596 ( .A1(n567), .A2(n529), .ZN(n540) );
  NOR2_X1 U597 ( .A1(n569), .A2(n540), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G141GAT), .B(KEYINPUT111), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1344GAT) );
  NOR2_X1 U600 ( .A1(n553), .A2(n540), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n533) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n532) );
  XNOR2_X1 U603 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U604 ( .A(KEYINPUT53), .B(n534), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(G1345GAT) );
  NOR2_X1 U606 ( .A1(n578), .A2(n540), .ZN(n538) );
  XNOR2_X1 U607 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U609 ( .A(G155GAT), .B(n539), .ZN(G1346GAT) );
  NOR2_X1 U610 ( .A1(n562), .A2(n540), .ZN(n541) );
  XOR2_X1 U611 ( .A(G162GAT), .B(n541), .Z(G1347GAT) );
  AND2_X1 U612 ( .A1(n542), .A2(n565), .ZN(n548) );
  XOR2_X1 U613 ( .A(KEYINPUT116), .B(n543), .Z(n545) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n548), .A2(n566), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT55), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n569), .A2(n561), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n294), .ZN(G1348GAT) );
  NOR2_X1 U620 ( .A1(n561), .A2(n553), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT119), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n578), .A2(n561), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n293), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n560) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U631 ( .A(n564), .B(n563), .Z(G1351GAT) );
  AND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n583) );
  NOR2_X1 U634 ( .A1(n569), .A2(n583), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n583), .A2(n573), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

