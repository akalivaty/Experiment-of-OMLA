//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n187), .B2(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT73), .B1(new_n187), .B2(G128), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G110), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  AOI211_X1 g018(.A(new_n201), .B(new_n203), .C1(KEYINPUT16), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(new_n203), .ZN(new_n207));
  AOI21_X1  g021(.A(G146), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n195), .B(new_n200), .C1(new_n205), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n191), .A2(new_n192), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT74), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n191), .A2(new_n192), .A3(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n211), .B(new_n213), .C1(new_n199), .C2(G110), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n215));
  INV_X1    g029(.A(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n202), .A2(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n214), .B2(KEYINPUT75), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n209), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XOR2_X1   g040(.A(new_n224), .B(new_n226), .Z(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n209), .B(new_n227), .C1(new_n215), .C2(new_n222), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n230), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(G234), .B2(new_n230), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n229), .A2(new_n231), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT30), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT11), .A2(G134), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G137), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n251), .A2(new_n256), .A3(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n248), .A2(new_n250), .A3(new_n253), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n247), .A2(G134), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n245), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G131), .ZN(new_n265));
  INV_X1    g079(.A(new_n246), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n249), .A2(G137), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT11), .B1(new_n247), .B2(G134), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n247), .A2(G134), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n258), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n265), .A2(new_n273), .A3(KEYINPUT66), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT1), .B1(new_n275), .B2(G146), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n201), .A2(G143), .ZN(new_n278));
  OAI211_X1 g092(.A(G128), .B(new_n276), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n201), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(G146), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n280), .B(new_n281), .C1(KEYINPUT1), .C2(new_n189), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n262), .A2(new_n263), .A3(new_n274), .A4(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n251), .B2(new_n256), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n273), .A3(KEYINPUT65), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n288), .B(G131), .C1(new_n251), .C2(new_n256), .ZN(new_n289));
  XNOR2_X1  g103(.A(G143), .B(G146), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT0), .A3(G128), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT0), .B(G128), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n287), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n285), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n265), .A2(new_n273), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n283), .B1(new_n297), .B2(new_n245), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n263), .B1(new_n298), .B2(new_n274), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n244), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(KEYINPUT69), .A2(G116), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT69), .A2(G116), .ZN(new_n302));
  OAI21_X1  g116(.A(G119), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G116), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G119), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT2), .A2(G113), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT68), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT2), .A3(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n309), .A2(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n306), .A3(new_n303), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n284), .A2(new_n273), .A3(new_n265), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n295), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(new_n244), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n300), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n322), .A2(new_n320), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n328));
  NOR2_X1   g142(.A1(G237), .A2(G953), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G210), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G101), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n325), .A2(new_n327), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT31), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n262), .A2(new_n274), .A3(new_n284), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT67), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n295), .A3(new_n285), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n320), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n333), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n325), .A2(new_n346), .A3(new_n327), .A4(new_n334), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n348), .B2(new_n349), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G472), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n337), .A2(new_n343), .A3(new_n338), .A4(new_n334), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n323), .B1(new_n342), .B2(new_n244), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n326), .B1(new_n357), .B2(new_n320), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n355), .B(new_n356), .C1(new_n358), .C2(new_n334), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n322), .A2(new_n320), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n333), .A2(new_n355), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n337), .A2(new_n338), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(new_n230), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n354), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n243), .B1(new_n353), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT93), .B1(new_n205), .B2(new_n208), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n207), .B1(new_n219), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n201), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n206), .A2(G146), .A3(new_n207), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G237), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n225), .A3(G214), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n275), .ZN(new_n377));
  AOI21_X1  g191(.A(G143), .B1(new_n329), .B2(G214), .ZN(new_n378));
  OAI21_X1  g192(.A(G131), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n275), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n329), .A2(G143), .A3(G214), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT88), .A3(G131), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n387));
  INV_X1    g201(.A(new_n384), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n258), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n381), .A3(new_n390), .A4(new_n385), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n374), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n388), .B1(new_n396), .B2(new_n258), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n384), .A2(KEYINPUT18), .A3(G131), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n204), .B(new_n201), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n392), .A2(KEYINPUT94), .A3(new_n395), .A4(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n217), .A2(new_n218), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT19), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n217), .A2(new_n218), .A3(new_n406), .A4(KEYINPUT19), .ZN(new_n410));
  AOI21_X1  g224(.A(G146), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n371), .B1(new_n411), .B2(KEYINPUT90), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n413), .B(G146), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT91), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n389), .A2(new_n381), .A3(new_n385), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT19), .B1(new_n204), .B2(new_n406), .ZN(new_n417));
  INV_X1    g231(.A(new_n410), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n201), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n413), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT90), .B(new_n201), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n371), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n400), .ZN(new_n425));
  INV_X1    g239(.A(new_n395), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT92), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n428), .B(new_n395), .C1(new_n424), .C2(new_n400), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n405), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n431));
  NOR2_X1   g245(.A1(G475), .A2(G902), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n432), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(KEYINPUT95), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT95), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(new_n405), .C1(new_n427), .C2(new_n429), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n434), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n433), .B1(new_n438), .B2(new_n431), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n392), .A2(new_n400), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n405), .B1(new_n395), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n230), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  XOR2_X1   g257(.A(KEYINPUT9), .B(G234), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n445), .A2(new_n237), .A3(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n275), .A2(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n189), .A2(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(G134), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n304), .A2(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT69), .B(G116), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(G122), .ZN(new_n454));
  OAI211_X1 g268(.A(KEYINPUT14), .B(G107), .C1(new_n304), .C2(G122), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n454), .B(G107), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n451), .B(new_n457), .C1(new_n458), .C2(new_n456), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT13), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n253), .B1(new_n449), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n450), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n447), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n459), .A3(new_n446), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n230), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n469), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n439), .A2(new_n443), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(G952), .A3(new_n225), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT21), .B(G898), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n290), .A2(new_n292), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n202), .B1(new_n492), .B2(new_n291), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n283), .A2(new_n202), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G224), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G953), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n496), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n502));
  INV_X1    g316(.A(G107), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(G104), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n394), .A2(G107), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G101), .ZN(new_n508));
  INV_X1    g322(.A(G101), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G101), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(new_n504), .C1(new_n506), .C2(new_n505), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n514), .A3(KEYINPUT4), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n516), .A3(G101), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n320), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n303), .A2(KEYINPUT5), .A3(new_n306), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT5), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n314), .B1(new_n305), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n305), .B1(new_n453), .B2(G119), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n519), .A2(new_n521), .B1(new_n522), .B2(new_n318), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n503), .A2(G104), .ZN(new_n524));
  OAI21_X1  g338(.A(G101), .B1(new_n506), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n510), .A2(new_n512), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n507), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(G110), .B(G122), .Z(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n518), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(KEYINPUT81), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n518), .A2(new_n529), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT80), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(new_n529), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n532), .B1(new_n539), .B2(KEYINPUT6), .ZN(new_n540));
  INV_X1    g354(.A(new_n538), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n518), .B2(new_n529), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT6), .B(new_n533), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n501), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G210), .B1(G237), .B2(G902), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n499), .A4(new_n495), .ZN(new_n548));
  INV_X1    g362(.A(new_n495), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n550));
  OAI22_X1  g364(.A1(new_n549), .A2(new_n493), .B1(new_n550), .B2(new_n498), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n532), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n307), .A2(new_n316), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n527), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n519), .A2(KEYINPUT82), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n303), .A2(new_n556), .A3(KEYINPUT5), .A4(new_n306), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n521), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT83), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n558), .A3(KEYINPUT83), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT84), .B1(new_n523), .B2(new_n528), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT84), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n519), .A2(new_n521), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n564), .B(new_n527), .C1(new_n565), .C2(new_n553), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n530), .B(KEYINPUT8), .Z(new_n568));
  AOI21_X1  g382(.A(new_n552), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n547), .B1(new_n569), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n568), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n566), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT83), .B1(new_n554), .B2(new_n558), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n574), .B2(new_n562), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT85), .B(new_n230), .C1(new_n575), .C2(new_n552), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n545), .A2(new_n546), .A3(new_n570), .A4(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n576), .A2(new_n570), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n546), .A4(new_n545), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n546), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n576), .A2(new_n570), .ZN(new_n585));
  INV_X1    g399(.A(new_n532), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n533), .B1(new_n541), .B2(new_n542), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT6), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n500), .B1(new_n589), .B2(new_n543), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n584), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(KEYINPUT86), .B(new_n584), .C1(new_n585), .C2(new_n590), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n491), .B1(new_n583), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G469), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n507), .A2(new_n516), .A3(G101), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n516), .B1(new_n507), .B2(G101), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n514), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT77), .B1(new_n527), .B2(new_n283), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n600), .A2(new_n294), .B1(new_n601), .B2(KEYINPUT10), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n287), .A2(new_n289), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT77), .B(new_n605), .C1(new_n527), .C2(new_n283), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n601), .A2(KEYINPUT10), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n294), .A2(new_n515), .A3(new_n517), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n604), .A3(new_n609), .A4(new_n606), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(G110), .B(G140), .ZN(new_n613));
  INV_X1    g427(.A(G227), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(G953), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n613), .B(new_n615), .Z(new_n616));
  INV_X1    g430(.A(new_n604), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n527), .B(new_n283), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT12), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT12), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n612), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n608), .A2(new_n606), .A3(new_n609), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n608), .A2(KEYINPUT79), .A3(new_n609), .A4(new_n606), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n616), .B1(new_n612), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n597), .B(new_n230), .C1(new_n624), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(G469), .A2(G902), .ZN(new_n632));
  INV_X1    g446(.A(new_n616), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n607), .B2(new_n611), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n629), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n607), .A2(new_n611), .B1(new_n621), .B2(new_n622), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n635), .B(G469), .C1(new_n616), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n631), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G221), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n444), .B2(new_n230), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n366), .A2(new_n479), .A3(new_n596), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT97), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n526), .ZN(G3));
  NAND2_X1  g460(.A1(new_n348), .A2(new_n230), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(G472), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n348), .A2(new_n349), .ZN(new_n649));
  INV_X1    g463(.A(new_n243), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n643), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n439), .A2(new_n443), .ZN(new_n653));
  AOI21_X1  g467(.A(G478), .B1(new_n468), .B2(new_n230), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  INV_X1    g469(.A(new_n467), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n446), .B1(new_n466), .B2(new_n459), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT33), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n468), .A2(KEYINPUT99), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n660), .B1(new_n663), .B2(KEYINPUT33), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n470), .A2(G902), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n489), .B(new_n487), .C1(new_n591), .C2(new_n577), .ZN(new_n668));
  AND4_X1   g482(.A1(KEYINPUT100), .A2(new_n653), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n666), .B1(new_n439), .B2(new_n443), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT100), .B1(new_n670), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n652), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(new_n487), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n443), .A2(new_n476), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n435), .A2(new_n437), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n431), .B1(new_n678), .B2(new_n432), .ZN(new_n679));
  AOI211_X1 g493(.A(KEYINPUT20), .B(new_n434), .C1(new_n435), .C2(new_n437), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n675), .B(new_n677), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n400), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n389), .A2(new_n381), .A3(new_n385), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n420), .A2(new_n371), .A3(new_n422), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(KEYINPUT91), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n684), .B1(new_n687), .B2(new_n423), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n428), .B1(new_n688), .B2(new_n395), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n425), .A2(KEYINPUT92), .A3(new_n426), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n436), .B1(new_n691), .B2(new_n405), .ZN(new_n692));
  INV_X1    g506(.A(new_n437), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n432), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT20), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n438), .A2(new_n431), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(KEYINPUT101), .A3(new_n675), .A4(new_n677), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n489), .B1(new_n591), .B2(new_n577), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n652), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT35), .B(G107), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  AND2_X1   g518(.A1(new_n348), .A2(new_n349), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n354), .B1(new_n348), .B2(new_n230), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n228), .A2(KEYINPUT36), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n223), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n223), .A2(new_n707), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n708), .A2(new_n241), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n236), .B2(new_n238), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n705), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n479), .A2(new_n596), .A3(new_n643), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT37), .B(G110), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G12));
  AOI21_X1  g529(.A(new_n642), .B1(new_n353), .B2(new_n365), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n481), .B1(new_n485), .B2(G900), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT102), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n676), .B(new_n718), .C1(new_n695), .C2(new_n696), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n489), .B(new_n711), .C1(new_n591), .C2(new_n577), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G128), .ZN(G30));
  XOR2_X1   g536(.A(new_n718), .B(KEYINPUT39), .Z(new_n723));
  NAND2_X1  g537(.A1(new_n643), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT40), .Z(new_n725));
  NAND2_X1  g539(.A1(new_n583), .A2(new_n595), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT38), .ZN(new_n727));
  INV_X1    g541(.A(new_n711), .ZN(new_n728));
  INV_X1    g542(.A(new_n360), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n333), .B1(new_n729), .B2(new_n326), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT103), .ZN(new_n731));
  INV_X1    g545(.A(new_n335), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n230), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G472), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n489), .B(new_n728), .C1(new_n353), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n477), .B1(new_n439), .B2(new_n443), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n725), .A2(new_n727), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G143), .ZN(G45));
  AOI211_X1 g552(.A(new_n718), .B(new_n666), .C1(new_n439), .C2(new_n443), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n716), .A3(new_n740), .A4(new_n720), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n742), .B(new_n365), .C1(new_n705), .C2(new_n351), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n720), .A3(new_n643), .ZN(new_n744));
  INV_X1    g558(.A(new_n718), .ZN(new_n745));
  INV_X1    g559(.A(new_n433), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n694), .B2(KEYINPUT20), .ZN(new_n747));
  INV_X1    g561(.A(G475), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n441), .B2(new_n230), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n667), .B(new_n745), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT104), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n741), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  NAND2_X1  g567(.A1(new_n612), .A2(new_n629), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n754), .A2(new_n633), .B1(new_n634), .B2(new_n623), .ZN(new_n755));
  OAI21_X1  g569(.A(G469), .B1(new_n755), .B2(G902), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n756), .A2(new_n641), .A3(new_n631), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n743), .A2(new_n650), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n669), .B2(new_n671), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NAND2_X1  g576(.A1(new_n701), .A2(new_n757), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n743), .A3(new_n650), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n683), .A3(new_n698), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G116), .ZN(G18));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n711), .A2(new_n487), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n701), .A2(new_n757), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n743), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n769), .B1(new_n772), .B2(new_n478), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n350), .A2(new_n352), .A3(new_n364), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n701), .A2(new_n757), .A3(new_n770), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT105), .A3(new_n479), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G119), .ZN(G21));
  INV_X1    g593(.A(new_n757), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n487), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n333), .B1(new_n339), .B2(new_n729), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n336), .A2(new_n347), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n349), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n706), .A3(new_n243), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n736), .A2(new_n781), .A3(new_n785), .A4(new_n701), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  NOR3_X1   g601(.A1(new_n784), .A2(new_n706), .A3(new_n711), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n750), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT106), .B1(new_n670), .B2(new_n745), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n764), .B(new_n788), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G125), .ZN(G27));
  NAND2_X1  g607(.A1(new_n750), .A2(new_n789), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n670), .A2(KEYINPUT106), .A3(new_n745), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n705), .A2(KEYINPUT32), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n365), .A2(new_n742), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n650), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n632), .B(KEYINPUT107), .Z(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n631), .A2(new_n637), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n641), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n583), .A2(new_n595), .A3(new_n804), .A4(new_n488), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n743), .A2(new_n650), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n805), .A3(KEYINPUT42), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n807), .A2(KEYINPUT42), .B1(new_n796), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G131), .ZN(G33));
  INV_X1    g625(.A(new_n594), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n545), .A2(new_n570), .A3(new_n576), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT86), .B1(new_n813), .B2(new_n584), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n815), .A2(new_n582), .A3(new_n803), .A4(new_n489), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n366), .A3(new_n719), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G134), .ZN(G36));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n747), .A2(new_n749), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n667), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT43), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(KEYINPUT43), .A3(new_n667), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(KEYINPUT108), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n711), .B1(new_n648), .B2(new_n649), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT108), .B1(new_n823), .B2(new_n824), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n819), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n828), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT44), .A3(new_n825), .A4(new_n826), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n583), .A2(new_n595), .A3(new_n488), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n635), .B1(new_n616), .B2(new_n636), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT45), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n597), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(KEYINPUT46), .A3(new_n801), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n631), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT46), .B1(new_n837), .B2(new_n801), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n641), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n723), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n829), .A2(new_n831), .A3(new_n833), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G137), .ZN(G39));
  OR2_X1    g661(.A1(new_n842), .A2(KEYINPUT47), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n842), .A2(KEYINPUT47), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n750), .A2(new_n832), .A3(new_n743), .A4(new_n650), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(new_n216), .ZN(G42));
  AOI21_X1  g666(.A(new_n481), .B1(new_n823), .B2(new_n824), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n785), .ZN(new_n854));
  INV_X1    g668(.A(new_n727), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n757), .A2(new_n489), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT114), .Z(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT50), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(new_n833), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n756), .A2(new_n631), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n848), .A2(new_n849), .B1(new_n640), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n832), .A2(new_n780), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n853), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n866), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n353), .A2(new_n734), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n868), .A2(new_n243), .A3(new_n481), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n653), .A2(new_n667), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n867), .A2(new_n788), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n860), .A2(new_n864), .A3(new_n865), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n864), .A2(new_n872), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n874), .B2(new_n859), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n788), .B(new_n816), .C1(new_n790), .C2(new_n791), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT112), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n796), .A2(new_n880), .A3(new_n788), .A4(new_n816), .ZN(new_n881));
  NOR4_X1   g695(.A1(new_n711), .A2(new_n476), .A3(new_n749), .A4(new_n718), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n833), .A2(new_n716), .A3(new_n697), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n796), .A2(new_n809), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n805), .B(new_n799), .C1(new_n794), .C2(new_n795), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT42), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n885), .B(new_n817), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n778), .A2(new_n760), .A3(new_n767), .A4(new_n786), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n786), .B1(new_n699), .B2(new_n765), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(KEYINPUT110), .A3(new_n760), .A4(new_n778), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n652), .A2(new_n596), .A3(new_n670), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n644), .A2(new_n897), .A3(new_n713), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n490), .B1(new_n815), .B2(new_n582), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n439), .A2(new_n677), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT111), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n747), .A2(new_n676), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT111), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n596), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n651), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n889), .A2(new_n896), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n803), .A2(new_n728), .A3(new_n718), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n869), .A2(new_n736), .A3(new_n701), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n792), .A2(new_n752), .A3(new_n721), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT52), .ZN(new_n911));
  INV_X1    g725(.A(new_n744), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n741), .A2(new_n751), .B1(new_n912), .B2(new_n719), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT52), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n792), .A4(new_n909), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n877), .B1(new_n907), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n911), .A2(new_n915), .ZN(new_n918));
  INV_X1    g732(.A(new_n906), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n892), .B2(new_n895), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT53), .A4(new_n889), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT113), .ZN(new_n925));
  INV_X1    g739(.A(new_n884), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT105), .B1(new_n776), .B2(new_n479), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n478), .A2(new_n774), .A3(new_n775), .A4(new_n769), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n653), .A2(new_n667), .A3(new_n668), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT100), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n670), .A2(KEYINPUT100), .A3(new_n668), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n758), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n929), .A2(new_n893), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n898), .A2(new_n905), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n926), .A2(new_n810), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n925), .B1(new_n938), .B2(new_n916), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n935), .A2(new_n937), .A3(new_n810), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n884), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(KEYINPUT113), .A3(new_n918), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n917), .A2(new_n924), .A3(new_n939), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT48), .ZN(new_n944));
  OAI221_X1 g758(.A(new_n650), .B1(KEYINPUT115), .B2(new_n944), .C1(new_n797), .C2(new_n798), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n867), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(KEYINPUT115), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n854), .A2(new_n764), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n225), .A2(G952), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n870), .B2(new_n670), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(KEYINPUT115), .B2(new_n944), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n876), .A2(new_n923), .A3(new_n943), .A4(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(G952), .B2(G953), .ZN(new_n956));
  OR4_X1    g770(.A1(new_n243), .A2(new_n821), .A3(new_n489), .A4(new_n640), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT109), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n862), .B(KEYINPUT49), .Z(new_n961));
  NOR3_X1   g775(.A1(new_n727), .A2(new_n869), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n956), .B1(new_n959), .B2(new_n963), .ZN(G75));
  NAND3_X1  g778(.A1(new_n917), .A2(new_n939), .A3(new_n942), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(G210), .A3(G902), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n540), .A2(new_n544), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n500), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n545), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(KEYINPUT116), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT56), .B1(new_n970), .B2(KEYINPUT116), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n966), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n225), .A2(G952), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(G51));
  XNOR2_X1  g790(.A(new_n800), .B(KEYINPUT57), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n918), .A2(new_n920), .A3(new_n889), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n916), .A2(new_n940), .A3(new_n884), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n877), .A2(new_n978), .B1(new_n979), .B2(KEYINPUT113), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n924), .B1(new_n980), .B2(new_n939), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n924), .A2(new_n917), .A3(new_n939), .A4(new_n942), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n755), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n230), .B1(new_n980), .B2(new_n939), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n837), .B(KEYINPUT117), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n975), .B1(new_n985), .B2(new_n988), .ZN(G54));
  NAND2_X1  g803(.A1(new_n965), .A2(G902), .ZN(new_n990));
  NAND2_X1  g804(.A1(KEYINPUT58), .A2(G475), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n435), .B(new_n437), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n975), .ZN(new_n993));
  INV_X1    g807(.A(new_n991), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n965), .A2(G902), .A3(new_n678), .A4(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n992), .A2(KEYINPUT118), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT118), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n678), .B1(new_n986), .B2(new_n994), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n993), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(G60));
  XNOR2_X1  g815(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n470), .A2(new_n230), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n664), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n981), .B2(new_n982), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n993), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1004), .B1(new_n923), .B2(new_n943), .ZN(new_n1010));
  OAI21_X1  g824(.A(KEYINPUT120), .B1(new_n1010), .B2(new_n664), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n924), .B1(new_n917), .B2(new_n921), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1005), .B1(new_n982), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT120), .ZN(new_n1014));
  INV_X1    g828(.A(new_n664), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1009), .B1(new_n1011), .B2(new_n1016), .ZN(G63));
  NAND2_X1  g831(.A1(G217), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT60), .Z(new_n1019));
  NAND2_X1  g833(.A1(new_n965), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n240), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n965), .A2(new_n708), .A3(new_n709), .A4(new_n1019), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1022), .A2(new_n993), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g838(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1022), .A2(new_n993), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(G66));
  OAI21_X1  g843(.A(G953), .B1(new_n484), .B2(new_n497), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n920), .B2(G953), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT123), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n967), .B1(G898), .B2(new_n225), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT124), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT122), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1032), .B(new_n1035), .ZN(G69));
  NOR2_X1   g850(.A1(new_n417), .A2(new_n418), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n357), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n851), .ZN(new_n1039));
  INV_X1    g853(.A(new_n888), .ZN(new_n1040));
  AND2_X1   g854(.A1(new_n913), .A2(new_n792), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n829), .A2(new_n831), .A3(new_n833), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n736), .A2(new_n701), .ZN(new_n1044));
  OR2_X1    g858(.A1(new_n1044), .A2(new_n799), .ZN(new_n1045));
  AND2_X1   g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1042), .B(KEYINPUT125), .C1(new_n1046), .C2(new_n844), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT125), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n844), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g865(.A(G953), .B(new_n1038), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(G900), .ZN(new_n1053));
  OAI21_X1  g867(.A(G953), .B1(new_n1038), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n900), .B1(new_n820), .B2(new_n666), .ZN(new_n1055));
  NOR3_X1   g869(.A1(new_n808), .A2(new_n832), .A3(new_n724), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n851), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1041), .A2(KEYINPUT62), .A3(new_n737), .ZN(new_n1058));
  AOI21_X1  g872(.A(KEYINPUT62), .B1(new_n1041), .B2(new_n737), .ZN(new_n1059));
  OAI211_X1 g873(.A(new_n1057), .B(new_n846), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1038), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1054), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g876(.A(G953), .B1(new_n614), .B2(new_n1053), .C1(new_n1038), .C2(KEYINPUT126), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1063), .ZN(new_n1064));
  OR3_X1    g878(.A1(new_n1052), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1064), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1065), .A2(new_n1066), .ZN(G72));
  INV_X1    g881(.A(KEYINPUT127), .ZN(new_n1068));
  NAND2_X1  g882(.A1(G472), .A2(G902), .ZN(new_n1069));
  XOR2_X1   g883(.A(new_n1069), .B(KEYINPUT63), .Z(new_n1070));
  INV_X1    g884(.A(new_n920), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n1070), .B1(new_n1060), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g886(.A1(new_n358), .A2(new_n333), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n975), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g888(.A(new_n922), .ZN(new_n1075));
  NOR2_X1   g889(.A1(new_n358), .A2(new_n334), .ZN(new_n1076));
  OAI21_X1  g890(.A(new_n1070), .B1(new_n1076), .B2(new_n732), .ZN(new_n1077));
  OAI21_X1  g891(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g892(.A(new_n358), .ZN(new_n1079));
  NOR2_X1   g893(.A1(new_n1079), .A2(new_n334), .ZN(new_n1080));
  INV_X1    g894(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g895(.A1(new_n1047), .A2(new_n920), .A3(new_n1051), .ZN(new_n1082));
  AOI21_X1  g896(.A(new_n1081), .B1(new_n1082), .B2(new_n1070), .ZN(new_n1083));
  OAI21_X1  g897(.A(new_n1068), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g898(.A1(new_n1082), .A2(new_n1070), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1085), .A2(new_n1080), .ZN(new_n1086));
  OR2_X1    g900(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1087));
  NAND4_X1  g901(.A1(new_n1086), .A2(KEYINPUT127), .A3(new_n1087), .A4(new_n1074), .ZN(new_n1088));
  NAND2_X1  g902(.A1(new_n1084), .A2(new_n1088), .ZN(G57));
endmodule


