

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n538), .A2(G2104), .ZN(n889) );
  INV_X1 U552 ( .A(n731), .ZN(n726) );
  INV_X1 U553 ( .A(KEYINPUT17), .ZN(n526) );
  AND2_X1 U554 ( .A1(n707), .A2(n532), .ZN(n711) );
  NAND2_X1 U555 ( .A1(n693), .A2(n781), .ZN(n731) );
  XNOR2_X1 U556 ( .A(n544), .B(n543), .ZN(G164) );
  NOR2_X2 U557 ( .A1(n563), .A2(n562), .ZN(G160) );
  NOR2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  NAND2_X1 U559 ( .A1(n522), .A2(n737), .ZN(n521) );
  XNOR2_X1 U560 ( .A(n735), .B(n734), .ZN(n522) );
  NAND2_X1 U561 ( .A1(G160), .A2(G40), .ZN(n780) );
  NOR2_X2 U562 ( .A1(G2104), .A2(n538), .ZN(n893) );
  AND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  XNOR2_X1 U564 ( .A(n525), .B(n524), .ZN(n523) );
  INV_X1 U565 ( .A(KEYINPUT65), .ZN(n524) );
  NAND2_X1 U566 ( .A1(n888), .A2(G137), .ZN(n525) );
  INV_X1 U567 ( .A(KEYINPUT27), .ZN(n714) );
  NOR2_X1 U568 ( .A1(n751), .A2(n530), .ZN(n529) );
  XNOR2_X1 U569 ( .A(n521), .B(n520), .ZN(n739) );
  XNOR2_X1 U570 ( .A(n738), .B(KEYINPUT93), .ZN(n520) );
  AND2_X1 U571 ( .A1(n731), .A2(n527), .ZN(n751) );
  AND2_X1 U572 ( .A1(n528), .A2(G8), .ZN(n527) );
  INV_X1 U573 ( .A(G1966), .ZN(n528) );
  INV_X1 U574 ( .A(n780), .ZN(n693) );
  AND2_X1 U575 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U576 ( .A1(n731), .A2(G8), .ZN(n776) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n781) );
  NAND2_X1 U578 ( .A1(n559), .A2(n523), .ZN(n563) );
  XNOR2_X1 U579 ( .A(n746), .B(n745), .ZN(n771) );
  AND2_X1 U580 ( .A1(n779), .A2(n778), .ZN(n519) );
  XNOR2_X2 U581 ( .A(n535), .B(n526), .ZN(n888) );
  INV_X1 U582 ( .A(n749), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n531), .A2(n529), .ZN(n732) );
  INV_X1 U584 ( .A(G8), .ZN(n530) );
  XNOR2_X1 U585 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U586 ( .A1(n726), .A2(G2072), .ZN(n715) );
  AND2_X1 U587 ( .A1(n706), .A2(n705), .ZN(n532) );
  XOR2_X1 U588 ( .A(n722), .B(KEYINPUT28), .Z(n533) );
  XOR2_X1 U589 ( .A(n603), .B(KEYINPUT71), .Z(n534) );
  INV_X1 U590 ( .A(KEYINPUT92), .ZN(n734) );
  INV_X1 U591 ( .A(KEYINPUT29), .ZN(n724) );
  XNOR2_X1 U592 ( .A(n725), .B(n724), .ZN(n730) );
  NAND2_X1 U593 ( .A1(n819), .A2(n815), .ZN(n807) );
  NOR2_X1 U594 ( .A1(G651), .A2(n647), .ZN(n659) );
  INV_X1 U595 ( .A(KEYINPUT87), .ZN(n544) );
  INV_X1 U596 ( .A(G2105), .ZN(n538) );
  NAND2_X1 U597 ( .A1(G126), .A2(n893), .ZN(n537) );
  NAND2_X1 U598 ( .A1(G138), .A2(n888), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G114), .A2(n894), .ZN(n540) );
  NAND2_X1 U601 ( .A1(G102), .A2(n889), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U604 ( .A1(G543), .A2(G651), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n545), .B(KEYINPUT64), .ZN(n655) );
  NAND2_X1 U606 ( .A1(G89), .A2(n655), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT0), .B(G543), .Z(n647) );
  INV_X1 U609 ( .A(G651), .ZN(n550) );
  NOR2_X1 U610 ( .A1(n647), .A2(n550), .ZN(n658) );
  NAND2_X1 U611 ( .A1(G76), .A2(n658), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(KEYINPUT5), .ZN(n556) );
  NOR2_X1 U614 ( .A1(G543), .A2(n550), .ZN(n551) );
  XOR2_X1 U615 ( .A(KEYINPUT1), .B(n551), .Z(n600) );
  BUF_X1 U616 ( .A(n600), .Z(n654) );
  NAND2_X1 U617 ( .A1(G63), .A2(n654), .ZN(n553) );
  NAND2_X1 U618 ( .A1(G51), .A2(n659), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n554), .Z(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(G101), .A2(n889), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT23), .B(n558), .Z(n559) );
  NAND2_X1 U626 ( .A1(G125), .A2(n893), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G113), .A2(n894), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n658), .A2(G72), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G85), .A2(n655), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G60), .A2(n654), .ZN(n567) );
  NAND2_X1 U633 ( .A1(G47), .A2(n659), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  OR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(G290) );
  AND2_X1 U636 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U637 ( .A(G57), .ZN(G237) );
  INV_X1 U638 ( .A(G132), .ZN(G219) );
  INV_X1 U639 ( .A(G82), .ZN(G220) );
  NAND2_X1 U640 ( .A1(n658), .A2(G75), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G88), .A2(n655), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT80), .B(n572), .Z(n576) );
  NAND2_X1 U644 ( .A1(G62), .A2(n654), .ZN(n574) );
  NAND2_X1 U645 ( .A1(G50), .A2(n659), .ZN(n573) );
  AND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(G303) );
  NAND2_X1 U648 ( .A1(G90), .A2(n655), .ZN(n577) );
  XOR2_X1 U649 ( .A(KEYINPUT67), .B(n577), .Z(n579) );
  NAND2_X1 U650 ( .A1(n658), .A2(G77), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U652 ( .A(n580), .B(KEYINPUT9), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G64), .A2(n654), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n659), .A2(G52), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT66), .B(n583), .Z(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G171) );
  NAND2_X1 U658 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U660 ( .A(G223), .ZN(n828) );
  NAND2_X1 U661 ( .A1(n828), .A2(G567), .ZN(n587) );
  XOR2_X1 U662 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U663 ( .A1(G56), .A2(n654), .ZN(n588) );
  XOR2_X1 U664 ( .A(KEYINPUT14), .B(n588), .Z(n594) );
  NAND2_X1 U665 ( .A1(G81), .A2(n655), .ZN(n589) );
  XNOR2_X1 U666 ( .A(n589), .B(KEYINPUT12), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G68), .A2(n658), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U669 ( .A(KEYINPUT13), .B(n592), .Z(n593) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n659), .A2(G43), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n995) );
  INV_X1 U673 ( .A(G860), .ZN(n620) );
  OR2_X1 U674 ( .A1(n995), .A2(n620), .ZN(n597) );
  XNOR2_X1 U675 ( .A(KEYINPUT70), .B(n597), .ZN(G153) );
  INV_X1 U676 ( .A(G171), .ZN(G301) );
  NAND2_X1 U677 ( .A1(G79), .A2(n658), .ZN(n599) );
  NAND2_X1 U678 ( .A1(G54), .A2(n659), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G66), .A2(n600), .ZN(n602) );
  NAND2_X1 U681 ( .A1(G92), .A2(n655), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n534), .ZN(n605) );
  XOR2_X1 U684 ( .A(KEYINPUT15), .B(n605), .Z(n606) );
  XNOR2_X2 U685 ( .A(KEYINPUT72), .B(n606), .ZN(n987) );
  NOR2_X1 U686 ( .A1(G868), .A2(n987), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT73), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U690 ( .A1(n658), .A2(G78), .ZN(n611) );
  NAND2_X1 U691 ( .A1(G91), .A2(n655), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT68), .B(n612), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G65), .A2(n654), .ZN(n613) );
  XNOR2_X1 U695 ( .A(KEYINPUT69), .B(n613), .ZN(n614) );
  NOR2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n659), .A2(G53), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(G299) );
  INV_X1 U699 ( .A(G868), .ZN(n624) );
  NOR2_X1 U700 ( .A1(G286), .A2(n624), .ZN(n619) );
  NOR2_X1 U701 ( .A1(G868), .A2(G299), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U703 ( .A1(n620), .A2(G559), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n621), .A2(n987), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n622), .B(KEYINPUT74), .ZN(n623) );
  XNOR2_X1 U706 ( .A(KEYINPUT16), .B(n623), .ZN(G148) );
  NOR2_X1 U707 ( .A1(G559), .A2(n624), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n625), .A2(n987), .ZN(n626) );
  XNOR2_X1 U709 ( .A(n626), .B(KEYINPUT75), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n995), .A2(G868), .ZN(n627) );
  NOR2_X1 U711 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U712 ( .A1(G123), .A2(n893), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n629), .B(KEYINPUT18), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT76), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G111), .A2(n894), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G135), .A2(n888), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G99), .A2(n889), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n936) );
  XNOR2_X1 U721 ( .A(n936), .B(G2096), .ZN(n638) );
  INV_X1 U722 ( .A(G2100), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(G156) );
  NAND2_X1 U724 ( .A1(G61), .A2(n654), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G86), .A2(n655), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n658), .A2(G73), .ZN(n641) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n659), .A2(G48), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n646) );
  XNOR2_X1 U733 ( .A(n646), .B(KEYINPUT78), .ZN(n652) );
  NAND2_X1 U734 ( .A1(G49), .A2(n659), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G87), .A2(n647), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U737 ( .A1(n654), .A2(n650), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U739 ( .A(KEYINPUT79), .B(n653), .Z(G288) );
  INV_X1 U740 ( .A(G299), .ZN(n983) );
  XNOR2_X1 U741 ( .A(n983), .B(G303), .ZN(n670) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n666) );
  NAND2_X1 U743 ( .A1(G67), .A2(n654), .ZN(n657) );
  NAND2_X1 U744 ( .A1(G93), .A2(n655), .ZN(n656) );
  NAND2_X1 U745 ( .A1(n657), .A2(n656), .ZN(n663) );
  NAND2_X1 U746 ( .A1(G80), .A2(n658), .ZN(n661) );
  NAND2_X1 U747 ( .A1(G55), .A2(n659), .ZN(n660) );
  NAND2_X1 U748 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U749 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U750 ( .A(KEYINPUT77), .B(n664), .Z(n837) );
  XNOR2_X1 U751 ( .A(G290), .B(n837), .ZN(n665) );
  XNOR2_X1 U752 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U753 ( .A(n667), .B(G288), .Z(n668) );
  XNOR2_X1 U754 ( .A(G305), .B(n668), .ZN(n669) );
  XNOR2_X1 U755 ( .A(n670), .B(n669), .ZN(n915) );
  NAND2_X1 U756 ( .A1(n987), .A2(G559), .ZN(n671) );
  XNOR2_X1 U757 ( .A(n995), .B(n671), .ZN(n836) );
  XOR2_X1 U758 ( .A(n915), .B(n836), .Z(n672) );
  NAND2_X1 U759 ( .A1(n672), .A2(G868), .ZN(n673) );
  XOR2_X1 U760 ( .A(KEYINPUT82), .B(n673), .Z(n675) );
  NOR2_X1 U761 ( .A1(n837), .A2(G868), .ZN(n674) );
  NOR2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U763 ( .A(KEYINPUT83), .B(n676), .ZN(G295) );
  NAND2_X1 U764 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XOR2_X1 U765 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n677) );
  XNOR2_X1 U766 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U767 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U768 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U769 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U770 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U774 ( .A1(G218), .A2(n683), .ZN(n684) );
  XOR2_X1 U775 ( .A(KEYINPUT85), .B(n684), .Z(n685) );
  NAND2_X1 U776 ( .A1(G96), .A2(n685), .ZN(n834) );
  NAND2_X1 U777 ( .A1(n834), .A2(G2106), .ZN(n689) );
  NAND2_X1 U778 ( .A1(G108), .A2(G120), .ZN(n686) );
  NOR2_X1 U779 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U780 ( .A1(G69), .A2(n687), .ZN(n835) );
  NAND2_X1 U781 ( .A1(n835), .A2(G567), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n926) );
  NOR2_X1 U783 ( .A1(n690), .A2(n926), .ZN(n691) );
  XNOR2_X1 U784 ( .A(n691), .B(KEYINPUT86), .ZN(n833) );
  NAND2_X1 U785 ( .A1(G36), .A2(n833), .ZN(G176) );
  XOR2_X1 U786 ( .A(KEYINPUT99), .B(G1981), .Z(n692) );
  XNOR2_X1 U787 ( .A(G305), .B(n692), .ZN(n997) );
  INV_X1 U788 ( .A(n776), .ZN(n694) );
  NOR2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NAND2_X1 U790 ( .A1(n694), .A2(n760), .ZN(n695) );
  NAND2_X1 U791 ( .A1(KEYINPUT33), .A2(n695), .ZN(n696) );
  NOR2_X1 U792 ( .A1(n997), .A2(n696), .ZN(n770) );
  NOR2_X1 U793 ( .A1(G1971), .A2(n776), .ZN(n698) );
  NOR2_X1 U794 ( .A1(G2090), .A2(n731), .ZN(n697) );
  NOR2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U796 ( .A(KEYINPUT95), .B(n699), .Z(n700) );
  NAND2_X1 U797 ( .A1(n700), .A2(G303), .ZN(n742) );
  AND2_X1 U798 ( .A1(n726), .A2(G2067), .ZN(n701) );
  XOR2_X1 U799 ( .A(n701), .B(KEYINPUT90), .Z(n703) );
  NAND2_X1 U800 ( .A1(n731), .A2(G1348), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n726), .A2(G1996), .ZN(n704) );
  XNOR2_X1 U803 ( .A(n704), .B(KEYINPUT26), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n731), .A2(G1341), .ZN(n706) );
  INV_X1 U805 ( .A(n995), .ZN(n705) );
  NAND2_X1 U806 ( .A1(n711), .A2(n987), .ZN(n708) );
  NAND2_X1 U807 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U808 ( .A(KEYINPUT91), .B(n710), .Z(n713) );
  OR2_X1 U809 ( .A1(n987), .A2(n711), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n731), .A2(G1956), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U813 ( .A(n718), .B(KEYINPUT89), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n983), .A2(n721), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U816 ( .A1(n983), .A2(n721), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n533), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G1961), .A2(n731), .ZN(n728) );
  XOR2_X1 U819 ( .A(G2078), .B(KEYINPUT25), .Z(n958) );
  NAND2_X1 U820 ( .A1(n726), .A2(n958), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n736) );
  OR2_X1 U822 ( .A1(G301), .A2(n736), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n740) );
  INV_X1 U824 ( .A(KEYINPUT31), .ZN(n738) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n731), .ZN(n749) );
  XNOR2_X1 U826 ( .A(n732), .B(KEYINPUT30), .ZN(n733) );
  NOR2_X1 U827 ( .A1(G168), .A2(n733), .ZN(n735) );
  NAND2_X1 U828 ( .A1(G301), .A2(n736), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n748) );
  NAND2_X1 U830 ( .A1(n748), .A2(G286), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U832 ( .A(n743), .B(KEYINPUT96), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n744), .A2(G8), .ZN(n746) );
  XOR2_X1 U834 ( .A(KEYINPUT97), .B(KEYINPUT32), .Z(n745) );
  INV_X1 U835 ( .A(KEYINPUT94), .ZN(n747) );
  XNOR2_X1 U836 ( .A(n748), .B(n747), .ZN(n753) );
  AND2_X1 U837 ( .A1(G8), .A2(n749), .ZN(n750) );
  OR2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n772) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n997), .ZN(n758) );
  AND2_X1 U841 ( .A1(n772), .A2(n758), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G288), .A2(G1976), .ZN(n754) );
  XOR2_X1 U843 ( .A(KEYINPUT98), .B(n754), .Z(n981) );
  INV_X1 U844 ( .A(n981), .ZN(n755) );
  AND2_X1 U845 ( .A1(n771), .A2(n757), .ZN(n767) );
  INV_X1 U846 ( .A(n758), .ZN(n761) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n979) );
  OR2_X1 U849 ( .A1(n761), .A2(n979), .ZN(n762) );
  OR2_X1 U850 ( .A1(n981), .A2(n762), .ZN(n765) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U852 ( .A(KEYINPUT24), .B(n763), .Z(n764) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n768), .A2(n776), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n779) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n775) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U862 ( .A1(n781), .A2(n780), .ZN(n822) );
  XNOR2_X1 U863 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NAND2_X1 U864 ( .A1(G140), .A2(n888), .ZN(n783) );
  NAND2_X1 U865 ( .A1(G104), .A2(n889), .ZN(n782) );
  NAND2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n784), .ZN(n789) );
  NAND2_X1 U868 ( .A1(G128), .A2(n893), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G116), .A2(n894), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U871 ( .A(KEYINPUT35), .B(n787), .Z(n788) );
  NOR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n790), .ZN(n912) );
  NOR2_X1 U874 ( .A1(n811), .A2(n912), .ZN(n927) );
  NAND2_X1 U875 ( .A1(n822), .A2(n927), .ZN(n819) );
  NAND2_X1 U876 ( .A1(G119), .A2(n893), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G131), .A2(n888), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G107), .A2(n894), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G95), .A2(n889), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n903) );
  NAND2_X1 U883 ( .A1(G1991), .A2(n903), .ZN(n806) );
  NAND2_X1 U884 ( .A1(G129), .A2(n893), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G117), .A2(n894), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n889), .A2(G105), .ZN(n799) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U890 ( .A(n802), .B(KEYINPUT88), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G141), .A2(n888), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n886) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n886), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n935) );
  NAND2_X1 U895 ( .A1(n822), .A2(n935), .ZN(n815) );
  NOR2_X1 U896 ( .A1(n519), .A2(n807), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(KEYINPUT100), .ZN(n810) );
  XNOR2_X1 U898 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U899 ( .A1(n993), .A2(n822), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n825) );
  NAND2_X1 U901 ( .A1(n811), .A2(n912), .ZN(n929) );
  NOR2_X1 U902 ( .A1(n886), .A2(G1996), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n812), .B(KEYINPUT101), .ZN(n941) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n903), .ZN(n937) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n937), .A2(n813), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT102), .B(n814), .Z(n816) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n941), .A2(n817), .ZN(n818) );
  XOR2_X1 U910 ( .A(KEYINPUT39), .B(n818), .Z(n820) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n929), .A2(n821), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n826) );
  XNOR2_X1 U916 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n828), .ZN(G217) );
  NAND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n829) );
  XNOR2_X1 U919 ( .A(KEYINPUT107), .B(n829), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n830), .A2(G661), .ZN(n831) );
  XNOR2_X1 U921 ( .A(KEYINPUT108), .B(n831), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U926 ( .A(G108), .ZN(G238) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  NOR2_X1 U930 ( .A1(n836), .A2(G860), .ZN(n838) );
  XNOR2_X1 U931 ( .A(n838), .B(n837), .ZN(G145) );
  XNOR2_X1 U932 ( .A(G2427), .B(G2451), .ZN(n848) );
  XOR2_X1 U933 ( .A(G2430), .B(G2443), .Z(n840) );
  XNOR2_X1 U934 ( .A(KEYINPUT105), .B(G2435), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U936 ( .A(G2438), .B(G2454), .Z(n842) );
  XNOR2_X1 U937 ( .A(G1341), .B(G1348), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U940 ( .A(KEYINPUT104), .B(G2446), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n849) );
  NAND2_X1 U943 ( .A1(n849), .A2(G14), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT106), .B(n850), .Z(G401) );
  XOR2_X1 U945 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n852) );
  XNOR2_X1 U946 ( .A(G2678), .B(KEYINPUT43), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n854) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U951 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U952 ( .A(G2096), .B(G2100), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U954 ( .A(G2084), .B(G2078), .Z(n859) );
  XNOR2_X1 U955 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U957 ( .A(G1961), .B(G1956), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U959 ( .A(n863), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(G2474), .B(G1981), .Z(n867) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1966), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G112), .A2(n894), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G100), .A2(n889), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U969 ( .A1(G136), .A2(n888), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n872), .B(KEYINPUT112), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G124), .A2(n893), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G130), .A2(n893), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G118), .A2(n894), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U978 ( .A1(n889), .A2(G106), .ZN(n880) );
  XOR2_X1 U979 ( .A(KEYINPUT113), .B(n880), .Z(n882) );
  NAND2_X1 U980 ( .A1(n888), .A2(G142), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n907) );
  XOR2_X1 U985 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n901) );
  NAND2_X1 U986 ( .A1(G139), .A2(n888), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT115), .B(n892), .Z(n899) );
  NAND2_X1 U990 ( .A1(G127), .A2(n893), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n930) );
  XNOR2_X1 U995 ( .A(n930), .B(KEYINPUT48), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U997 ( .A(KEYINPUT46), .B(n902), .ZN(n905) );
  XNOR2_X1 U998 ( .A(n903), .B(KEYINPUT114), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1001 ( .A(n936), .B(G162), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G164), .B(G160), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1005 ( .A(n913), .B(n912), .Z(n914) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n914), .ZN(G395) );
  XOR2_X1 U1007 ( .A(KEYINPUT118), .B(n915), .Z(n917) );
  XOR2_X1 U1008 ( .A(n987), .B(G286), .Z(n916) );
  XNOR2_X1 U1009 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1010 ( .A(n995), .B(G171), .ZN(n918) );
  XNOR2_X1 U1011 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n920), .ZN(G397) );
  OR2_X1 U1013 ( .A1(n926), .A2(G401), .ZN(n923) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G303), .ZN(G166) );
  INV_X1 U1021 ( .A(n926), .ZN(G319) );
  INV_X1 U1022 ( .A(G69), .ZN(G235) );
  INV_X1 U1023 ( .A(n927), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n950) );
  XOR2_X1 U1025 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(KEYINPUT50), .B(n933), .ZN(n948) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n940) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1032 ( .A(KEYINPUT119), .B(n938), .Z(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G162), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n943), .B(KEYINPUT120), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n944), .Z(n945) );
  NOR2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1040 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n973) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n973), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(n953), .A2(G29), .ZN(n1033) );
  XOR2_X1 U1045 ( .A(KEYINPUT122), .B(G34), .Z(n955) );
  XNOR2_X1 U1046 ( .A(G2084), .B(KEYINPUT54), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n955), .B(n954), .ZN(n971) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n969) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G32), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G2072), .B(G33), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G27), .B(n958), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n966) );
  XOR2_X1 U1056 ( .A(G1991), .B(G25), .Z(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(G28), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT121), .B(n964), .Z(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(n967), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n973), .B(n972), .ZN(n975) );
  INV_X1 U1064 ( .A(G29), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n976), .ZN(n1031) );
  INV_X1 U1067 ( .A(G16), .ZN(n1027) );
  XNOR2_X1 U1068 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n1027), .B(n977), .ZN(n1004) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(n982), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n983), .B(G1956), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n986), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(G301), .B(G1961), .ZN(n989) );
  XOR2_X1 U1078 ( .A(n987), .B(G1348), .Z(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n994), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(n995), .B(G1341), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(G1966), .B(G168), .Z(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT57), .B(n998), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1029) );
  XOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(G4), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1956), .B(G20), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1012), .B(KEYINPUT127), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1013), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G21), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G5), .B(G1961), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1024) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G23), .B(G1976), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(G1986), .B(G24), .Z(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT58), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

