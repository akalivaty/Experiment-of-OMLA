

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845;

  OR2_X1 U371 ( .A1(n740), .A2(G902), .ZN(n591) );
  XNOR2_X1 U372 ( .A(n573), .B(n446), .ZN(n445) );
  INV_X1 U373 ( .A(G902), .ZN(n460) );
  XNOR2_X1 U374 ( .A(n350), .B(KEYINPUT77), .ZN(n428) );
  NAND2_X1 U375 ( .A1(n415), .A2(n416), .ZN(n350) );
  OR2_X2 U376 ( .A1(n756), .A2(n459), .ZN(n458) );
  AND2_X1 U377 ( .A1(n645), .A2(n363), .ZN(n653) );
  XNOR2_X1 U378 ( .A(n639), .B(n638), .ZN(n645) );
  XNOR2_X2 U379 ( .A(n575), .B(n563), .ZN(n775) );
  XNOR2_X1 U380 ( .A(G101), .B(KEYINPUT79), .ZN(n492) );
  BUF_X1 U381 ( .A(n732), .Z(n735) );
  NAND2_X2 U382 ( .A1(n468), .A2(n466), .ZN(n696) );
  AND2_X2 U383 ( .A1(n379), .A2(n380), .ZN(n468) );
  OR2_X2 U384 ( .A1(n470), .A2(n469), .ZN(n380) );
  XNOR2_X2 U385 ( .A(G116), .B(G113), .ZN(n465) );
  XNOR2_X2 U386 ( .A(n635), .B(KEYINPUT1), .ZN(n676) );
  INV_X1 U387 ( .A(n695), .ZN(n799) );
  NOR2_X1 U388 ( .A1(n659), .A2(n834), .ZN(n386) );
  INV_X1 U389 ( .A(n816), .ZN(n413) );
  AND2_X1 U390 ( .A1(n434), .A2(n432), .ZN(n431) );
  AND2_X1 U391 ( .A1(n358), .A2(n357), .ZN(n356) );
  XNOR2_X1 U392 ( .A(n500), .B(n460), .ZN(n737) );
  INV_X1 U393 ( .A(KEYINPUT109), .ZN(n362) );
  NAND2_X1 U394 ( .A1(n359), .A2(n356), .ZN(n355) );
  OR2_X1 U395 ( .A1(n762), .A2(n360), .ZN(n359) );
  NOR2_X1 U396 ( .A1(n736), .A2(n377), .ZN(n388) );
  NAND2_X1 U397 ( .A1(n365), .A2(n407), .ZN(n405) );
  NOR2_X1 U398 ( .A1(n396), .A2(n395), .ZN(n398) );
  AND2_X1 U399 ( .A1(n425), .A2(n712), .ZN(n713) );
  AND2_X1 U400 ( .A1(n451), .A2(n384), .ZN(n415) );
  NAND2_X1 U401 ( .A1(n394), .A2(n390), .ZN(n397) );
  NAND2_X1 U402 ( .A1(n413), .A2(n419), .ZN(n394) );
  XNOR2_X1 U403 ( .A(n386), .B(n385), .ZN(n730) );
  XNOR2_X1 U404 ( .A(n652), .B(n362), .ZN(n416) );
  NAND2_X1 U405 ( .A1(n431), .A2(n430), .ZN(n626) );
  NAND2_X1 U406 ( .A1(n429), .A2(n611), .ZN(n623) );
  NAND2_X1 U407 ( .A1(n778), .A2(n361), .ZN(n358) );
  INV_X1 U408 ( .A(n634), .ZN(n429) );
  NAND2_X1 U409 ( .A1(n461), .A2(n458), .ZN(n695) );
  INV_X1 U410 ( .A(n807), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n492), .B(G110), .ZN(n444) );
  INV_X1 U412 ( .A(n737), .ZN(n352) );
  INV_X4 U413 ( .A(G953), .ZN(n532) );
  XNOR2_X1 U414 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n500) );
  NAND2_X2 U415 ( .A1(n655), .A2(n556), .ZN(n557) );
  XNOR2_X2 U416 ( .A(n353), .B(n525), .ZN(n655) );
  NAND2_X2 U417 ( .A1(n435), .A2(n524), .ZN(n353) );
  NAND2_X2 U418 ( .A1(n383), .A2(n410), .ZN(n435) );
  NOR2_X1 U419 ( .A1(n355), .A2(n354), .ZN(G54) );
  AND2_X1 U420 ( .A1(n762), .A2(n778), .ZN(n354) );
  INV_X1 U421 ( .A(n779), .ZN(n357) );
  OR2_X1 U422 ( .A1(n778), .A2(n361), .ZN(n360) );
  INV_X1 U423 ( .A(G469), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n416), .B(G143), .ZN(G45) );
  AND2_X1 U425 ( .A1(n645), .A2(n644), .ZN(n651) );
  AND2_X1 U426 ( .A1(n644), .A2(n351), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n590), .ZN(n367) );
  NOR2_X1 U428 ( .A1(n586), .A2(n739), .ZN(n364) );
  XNOR2_X2 U429 ( .A(n411), .B(n489), .ZN(n683) );
  XNOR2_X2 U430 ( .A(n683), .B(G146), .ZN(n575) );
  XNOR2_X2 U431 ( .A(n441), .B(n692), .ZN(n748) );
  XNOR2_X2 U432 ( .A(n445), .B(n562), .ZN(n692) );
  OR2_X1 U433 ( .A1(n713), .A2(KEYINPUT89), .ZN(n475) );
  INV_X1 U434 ( .A(KEYINPUT28), .ZN(n457) );
  NAND2_X1 U435 ( .A1(G472), .A2(n460), .ZN(n459) );
  AND2_X1 U436 ( .A1(n463), .A2(n462), .ZN(n461) );
  NAND2_X1 U437 ( .A1(n478), .A2(n714), .ZN(n477) );
  INV_X1 U438 ( .A(KEYINPUT89), .ZN(n478) );
  NAND2_X1 U439 ( .A1(n426), .A2(n711), .ZN(n425) );
  NAND2_X1 U440 ( .A1(n710), .A2(n838), .ZN(n426) );
  INV_X1 U441 ( .A(KEYINPUT46), .ZN(n661) );
  NAND2_X1 U442 ( .A1(n504), .A2(G210), .ZN(n507) );
  XNOR2_X1 U443 ( .A(G134), .B(G131), .ZN(n558) );
  NOR2_X1 U444 ( .A1(G953), .A2(G237), .ZN(n566) );
  XNOR2_X1 U445 ( .A(KEYINPUT10), .B(G140), .ZN(n544) );
  OR2_X1 U446 ( .A1(n807), .A2(n640), .ZN(n621) );
  NAND2_X1 U447 ( .A1(n703), .A2(n704), .ZN(n420) );
  NOR2_X1 U448 ( .A1(n461), .A2(n457), .ZN(n454) );
  NAND2_X1 U449 ( .A1(n455), .A2(n461), .ZN(n434) );
  NOR2_X1 U450 ( .A1(n456), .A2(n623), .ZN(n455) );
  INV_X1 U451 ( .A(KEYINPUT0), .ZN(n525) );
  XNOR2_X1 U452 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n534) );
  XNOR2_X1 U453 ( .A(n577), .B(KEYINPUT23), .ZN(n579) );
  XNOR2_X1 U454 ( .A(G110), .B(KEYINPUT24), .ZN(n577) );
  AND2_X1 U455 ( .A1(n709), .A2(KEYINPUT34), .ZN(n419) );
  INV_X1 U456 ( .A(KEYINPUT67), .ZN(n437) );
  XNOR2_X1 U457 ( .A(n490), .B(G122), .ZN(n446) );
  XNOR2_X1 U458 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n490) );
  NAND2_X1 U459 ( .A1(n672), .A2(n671), .ZN(n384) );
  NAND2_X1 U460 ( .A1(G953), .A2(G902), .ZN(n603) );
  AND2_X1 U461 ( .A1(n479), .A2(n474), .ZN(n473) );
  NAND2_X1 U462 ( .A1(n472), .A2(n373), .ZN(n471) );
  INV_X1 U463 ( .A(G237), .ZN(n501) );
  NAND2_X1 U464 ( .A1(n458), .A2(n457), .ZN(n456) );
  INV_X1 U465 ( .A(KEYINPUT103), .ZN(n469) );
  XNOR2_X1 U466 ( .A(G113), .B(G104), .ZN(n540) );
  XOR2_X1 U467 ( .A(KEYINPUT12), .B(G122), .Z(n541) );
  XNOR2_X1 U468 ( .A(G137), .B(KEYINPUT71), .ZN(n582) );
  INV_X1 U469 ( .A(KEYINPUT4), .ZN(n499) );
  INV_X1 U470 ( .A(KEYINPUT80), .ZN(n638) );
  XNOR2_X1 U471 ( .A(n507), .B(KEYINPUT93), .ZN(n617) );
  AND2_X1 U472 ( .A1(n695), .A2(KEYINPUT67), .ZN(n440) );
  OR2_X1 U473 ( .A1(n695), .A2(KEYINPUT67), .ZN(n438) );
  XNOR2_X1 U474 ( .A(G101), .B(KEYINPUT78), .ZN(n569) );
  XOR2_X1 U475 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n568) );
  XNOR2_X1 U476 ( .A(G107), .B(G104), .ZN(n491) );
  XNOR2_X1 U477 ( .A(G116), .B(G134), .ZN(n526) );
  XNOR2_X1 U478 ( .A(G107), .B(G122), .ZN(n527) );
  XOR2_X1 U479 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n528) );
  NAND2_X1 U480 ( .A1(G237), .A2(G234), .ZN(n520) );
  NAND2_X1 U481 ( .A1(n452), .A2(KEYINPUT2), .ZN(n783) );
  XNOR2_X1 U482 ( .A(n622), .B(KEYINPUT41), .ZN(n805) );
  NAND2_X1 U483 ( .A1(n506), .A2(n352), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n648), .A2(n427), .ZN(n400) );
  NOR2_X1 U485 ( .A1(n412), .A2(n399), .ZN(n395) );
  AND2_X1 U486 ( .A1(n412), .A2(n372), .ZN(n390) );
  NAND2_X1 U487 ( .A1(n424), .A2(n799), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n626), .B(n625), .ZN(n628) );
  NAND2_X1 U489 ( .A1(n408), .A2(n375), .ZN(n402) );
  XNOR2_X1 U490 ( .A(n585), .B(n684), .ZN(n740) );
  XNOR2_X1 U491 ( .A(n579), .B(n578), .ZN(n580) );
  BUF_X1 U492 ( .A(n774), .Z(n762) );
  XNOR2_X1 U493 ( .A(n767), .B(KEYINPUT59), .ZN(n768) );
  NOR2_X1 U494 ( .A1(n774), .A2(n745), .ZN(n422) );
  NAND2_X1 U495 ( .A1(n742), .A2(G953), .ZN(n770) );
  INV_X1 U496 ( .A(KEYINPUT40), .ZN(n385) );
  XNOR2_X1 U497 ( .A(n656), .B(KEYINPUT31), .ZN(n710) );
  NOR2_X1 U498 ( .A1(n703), .A2(n423), .ZN(n656) );
  AND2_X1 U499 ( .A1(n439), .A2(n374), .ZN(n365) );
  AND2_X1 U500 ( .A1(n438), .A2(n429), .ZN(n366) );
  AND2_X1 U501 ( .A1(n467), .A2(n470), .ZN(n368) );
  AND2_X1 U502 ( .A1(n518), .A2(KEYINPUT19), .ZN(n369) );
  AND2_X1 U503 ( .A1(n419), .A2(n401), .ZN(n370) );
  AND2_X1 U504 ( .A1(n470), .A2(n469), .ZN(n371) );
  AND2_X1 U505 ( .A1(n420), .A2(n427), .ZN(n372) );
  AND2_X1 U506 ( .A1(n705), .A2(KEYINPUT35), .ZN(n401) );
  AND2_X1 U507 ( .A1(n713), .A2(n478), .ZN(n373) );
  AND2_X1 U508 ( .A1(n366), .A2(n436), .ZN(n374) );
  AND2_X1 U509 ( .A1(n437), .A2(KEYINPUT104), .ZN(n375) );
  INV_X1 U510 ( .A(KEYINPUT35), .ZN(n427) );
  XOR2_X1 U511 ( .A(n748), .B(n747), .Z(n376) );
  AND2_X1 U512 ( .A1(n738), .A2(n781), .ZN(n377) );
  AND2_X1 U513 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n378) );
  NAND2_X1 U514 ( .A1(n476), .A2(n475), .ZN(n474) );
  NAND2_X1 U515 ( .A1(n398), .A2(n397), .ZN(n715) );
  INV_X1 U516 ( .A(n698), .ZN(n424) );
  NAND2_X1 U517 ( .A1(n595), .A2(KEYINPUT103), .ZN(n379) );
  NAND2_X1 U518 ( .A1(n676), .A2(n654), .ZN(n698) );
  XNOR2_X1 U519 ( .A(n493), .B(n545), .ZN(n443) );
  INV_X1 U520 ( .A(n413), .ZN(n381) );
  INV_X1 U521 ( .A(n470), .ZN(n382) );
  XNOR2_X1 U522 ( .A(n702), .B(n701), .ZN(n816) );
  INV_X1 U523 ( .A(n736), .ZN(n452) );
  BUF_X1 U524 ( .A(n733), .Z(n736) );
  NOR2_X1 U525 ( .A1(n454), .A2(n624), .ZN(n430) );
  NAND2_X1 U526 ( .A1(n651), .A2(n650), .ZN(n652) );
  OR2_X1 U527 ( .A1(n748), .A2(n737), .ZN(n616) );
  NAND2_X1 U528 ( .A1(n417), .A2(n697), .ZN(n717) );
  NAND2_X1 U529 ( .A1(n409), .A2(n519), .ZN(n383) );
  OR2_X2 U530 ( .A1(n748), .A2(n418), .ZN(n518) );
  NAND2_X1 U531 ( .A1(n634), .A2(n633), .ZN(n792) );
  XNOR2_X2 U532 ( .A(n367), .B(n591), .ZN(n634) );
  XNOR2_X1 U533 ( .A(n496), .B(n443), .ZN(n442) );
  XNOR2_X1 U534 ( .A(n387), .B(n679), .ZN(n447) );
  NAND2_X1 U535 ( .A1(n449), .A2(n448), .ZN(n387) );
  AND2_X2 U536 ( .A1(n516), .A2(n515), .ZN(n517) );
  NAND2_X1 U537 ( .A1(n735), .A2(n388), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n389), .A2(n401), .ZN(n393) );
  INV_X1 U539 ( .A(n420), .ZN(n389) );
  NAND2_X1 U540 ( .A1(n392), .A2(n391), .ZN(n396) );
  NAND2_X1 U541 ( .A1(n370), .A2(n413), .ZN(n391) );
  AND2_X1 U542 ( .A1(n393), .A2(n400), .ZN(n392) );
  INV_X1 U543 ( .A(n401), .ZN(n399) );
  AND2_X2 U544 ( .A1(n403), .A2(n402), .ZN(n406) );
  NAND2_X1 U545 ( .A1(n404), .A2(KEYINPUT104), .ZN(n403) );
  NAND2_X1 U546 ( .A1(n439), .A2(n366), .ZN(n404) );
  NAND2_X2 U547 ( .A1(n406), .A2(n405), .ZN(n417) );
  NAND2_X1 U548 ( .A1(n408), .A2(n437), .ZN(n407) );
  INV_X1 U549 ( .A(n696), .ZN(n408) );
  NAND2_X1 U550 ( .A1(n517), .A2(n518), .ZN(n409) );
  NAND2_X1 U551 ( .A1(n369), .A2(n517), .ZN(n410) );
  NAND2_X1 U552 ( .A1(n517), .A2(n518), .ZN(n673) );
  XNOR2_X1 U553 ( .A(n411), .B(n442), .ZN(n441) );
  XNOR2_X2 U554 ( .A(n531), .B(n499), .ZN(n411) );
  NAND2_X1 U555 ( .A1(n816), .A2(n704), .ZN(n412) );
  XNOR2_X1 U556 ( .A(n417), .B(G110), .ZN(G12) );
  XNOR2_X1 U557 ( .A(n422), .B(n376), .ZN(n749) );
  XNOR2_X1 U558 ( .A(n421), .B(n744), .ZN(G66) );
  NAND2_X1 U559 ( .A1(n743), .A2(n770), .ZN(n421) );
  AND2_X1 U560 ( .A1(n789), .A2(n737), .ZN(n487) );
  NAND2_X1 U561 ( .A1(n484), .A2(n483), .ZN(n482) );
  XNOR2_X1 U562 ( .A(n662), .B(n661), .ZN(n448) );
  NAND2_X1 U563 ( .A1(n803), .A2(n423), .ZN(n804) );
  INV_X1 U564 ( .A(n715), .ZN(n753) );
  NAND2_X1 U565 ( .A1(n428), .A2(n843), .ZN(n678) );
  OR2_X1 U566 ( .A1(n634), .A2(n633), .ZN(n797) );
  AND2_X1 U567 ( .A1(n676), .A2(n429), .ZN(n593) );
  NAND2_X1 U568 ( .A1(n433), .A2(KEYINPUT28), .ZN(n432) );
  NAND2_X1 U569 ( .A1(n453), .A2(n458), .ZN(n433) );
  NAND2_X1 U570 ( .A1(n628), .A2(n435), .ZN(n668) );
  INV_X1 U571 ( .A(KEYINPUT104), .ZN(n436) );
  NAND2_X1 U572 ( .A1(n696), .A2(n440), .ZN(n439) );
  XNOR2_X2 U573 ( .A(n498), .B(n497), .ZN(n531) );
  XNOR2_X2 U574 ( .A(n444), .B(n491), .ZN(n562) );
  XNOR2_X2 U575 ( .A(n465), .B(n464), .ZN(n573) );
  NAND2_X1 U576 ( .A1(n447), .A2(n682), .ZN(n733) );
  XNOR2_X1 U577 ( .A(n678), .B(KEYINPUT73), .ZN(n449) );
  NAND2_X1 U578 ( .A1(n450), .A2(n667), .ZN(n451) );
  NAND2_X1 U579 ( .A1(n665), .A2(n664), .ZN(n450) );
  INV_X1 U580 ( .A(n623), .ZN(n453) );
  NAND2_X1 U581 ( .A1(n754), .A2(G902), .ZN(n462) );
  NAND2_X1 U582 ( .A1(n756), .A2(n754), .ZN(n463) );
  XNOR2_X2 U583 ( .A(n557), .B(KEYINPUT22), .ZN(n595) );
  XNOR2_X2 U584 ( .A(KEYINPUT3), .B(G119), .ZN(n464) );
  NAND2_X1 U585 ( .A1(n467), .A2(n371), .ZN(n466) );
  INV_X1 U586 ( .A(n595), .ZN(n467) );
  INV_X1 U587 ( .A(n676), .ZN(n470) );
  NAND2_X1 U588 ( .A1(n473), .A2(n471), .ZN(n721) );
  INV_X1 U589 ( .A(n480), .ZN(n472) );
  NAND2_X1 U590 ( .A1(n713), .A2(n477), .ZN(n476) );
  NAND2_X1 U591 ( .A1(n480), .A2(n378), .ZN(n479) );
  NAND2_X1 U592 ( .A1(n706), .A2(n715), .ZN(n480) );
  INV_X1 U593 ( .A(n735), .ZN(n780) );
  XNOR2_X2 U594 ( .A(n482), .B(n481), .ZN(n774) );
  INV_X1 U595 ( .A(KEYINPUT65), .ZN(n481) );
  NAND2_X1 U596 ( .A1(n486), .A2(n485), .ZN(n484) );
  INV_X1 U597 ( .A(KEYINPUT87), .ZN(n485) );
  NAND2_X1 U598 ( .A1(n488), .A2(n487), .ZN(n486) );
  INV_X1 U599 ( .A(n734), .ZN(n488) );
  XOR2_X1 U600 ( .A(n558), .B(KEYINPUT72), .Z(n489) );
  INV_X1 U601 ( .A(n792), .ZN(n654) );
  XNOR2_X1 U602 ( .A(n722), .B(KEYINPUT45), .ZN(n732) );
  XNOR2_X2 U603 ( .A(G146), .B(G125), .ZN(n545) );
  XNOR2_X1 U604 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n493) );
  XNOR2_X1 U605 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n495) );
  NAND2_X1 U606 ( .A1(n532), .A2(G224), .ZN(n494) );
  XNOR2_X1 U607 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X2 U608 ( .A(G143), .B(KEYINPUT64), .ZN(n498) );
  INV_X1 U609 ( .A(G128), .ZN(n497) );
  NAND2_X1 U610 ( .A1(n460), .A2(n501), .ZN(n504) );
  INV_X1 U611 ( .A(KEYINPUT90), .ZN(n502) );
  XNOR2_X1 U612 ( .A(n502), .B(KEYINPUT93), .ZN(n503) );
  XNOR2_X1 U613 ( .A(n507), .B(n503), .ZN(n505) );
  AND2_X1 U614 ( .A1(n504), .A2(G214), .ZN(n640) );
  INV_X1 U615 ( .A(n640), .ZN(n808) );
  AND2_X1 U616 ( .A1(n505), .A2(n808), .ZN(n506) );
  OR2_X1 U617 ( .A1(n617), .A2(KEYINPUT90), .ZN(n511) );
  INV_X1 U618 ( .A(n617), .ZN(n509) );
  NAND2_X1 U619 ( .A1(n808), .A2(KEYINPUT90), .ZN(n508) );
  OR2_X1 U620 ( .A1(n509), .A2(n508), .ZN(n510) );
  NAND2_X1 U621 ( .A1(n511), .A2(n510), .ZN(n512) );
  NAND2_X1 U622 ( .A1(n748), .A2(n512), .ZN(n516) );
  NAND2_X1 U623 ( .A1(n512), .A2(n737), .ZN(n514) );
  OR2_X1 U624 ( .A1(n808), .A2(KEYINPUT90), .ZN(n513) );
  AND2_X1 U625 ( .A1(n514), .A2(n513), .ZN(n515) );
  INV_X1 U626 ( .A(KEYINPUT19), .ZN(n519) );
  XNOR2_X1 U627 ( .A(n520), .B(KEYINPUT14), .ZN(n822) );
  NAND2_X1 U628 ( .A1(n532), .A2(G952), .ZN(n607) );
  INV_X1 U629 ( .A(G898), .ZN(n693) );
  INV_X1 U630 ( .A(n603), .ZN(n521) );
  NAND2_X1 U631 ( .A1(n693), .A2(n521), .ZN(n522) );
  NAND2_X1 U632 ( .A1(n607), .A2(n522), .ZN(n523) );
  AND2_X1 U633 ( .A1(n822), .A2(n523), .ZN(n524) );
  XNOR2_X1 U634 ( .A(n526), .B(KEYINPUT100), .ZN(n530) );
  XNOR2_X1 U635 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U636 ( .A(n530), .B(n529), .Z(n537) );
  AND2_X1 U637 ( .A1(n532), .A2(G234), .ZN(n533) );
  XNOR2_X1 U638 ( .A(n534), .B(n533), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n576), .A2(G217), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n531), .B(n535), .ZN(n536) );
  XNOR2_X1 U641 ( .A(n537), .B(n536), .ZN(n763) );
  NAND2_X1 U642 ( .A1(n763), .A2(n460), .ZN(n538) );
  INV_X1 U643 ( .A(G478), .ZN(n761) );
  XNOR2_X1 U644 ( .A(n538), .B(n761), .ZN(n646) );
  XNOR2_X1 U645 ( .A(G143), .B(G131), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n539), .B(KEYINPUT11), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U648 ( .A(n543), .B(n542), .Z(n548) );
  XNOR2_X1 U649 ( .A(n545), .B(n544), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n566), .A2(G214), .ZN(n546) );
  XNOR2_X1 U651 ( .A(n584), .B(n546), .ZN(n547) );
  XNOR2_X1 U652 ( .A(n548), .B(n547), .ZN(n767) );
  NAND2_X1 U653 ( .A1(n767), .A2(n460), .ZN(n551) );
  XNOR2_X1 U654 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n549) );
  INV_X1 U655 ( .A(G475), .ZN(n766) );
  XNOR2_X1 U656 ( .A(n549), .B(n766), .ZN(n550) );
  XNOR2_X1 U657 ( .A(n551), .B(n550), .ZN(n647) );
  NAND2_X1 U658 ( .A1(n646), .A2(n647), .ZN(n811) );
  NAND2_X1 U659 ( .A1(n352), .A2(G234), .ZN(n553) );
  XNOR2_X1 U660 ( .A(KEYINPUT95), .B(KEYINPUT20), .ZN(n552) );
  XNOR2_X1 U661 ( .A(n553), .B(n552), .ZN(n586) );
  INV_X1 U662 ( .A(G221), .ZN(n554) );
  OR2_X1 U663 ( .A1(n586), .A2(n554), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n555), .B(KEYINPUT21), .ZN(n796) );
  NOR2_X1 U665 ( .A1(n811), .A2(n796), .ZN(n556) );
  NAND2_X1 U666 ( .A1(n532), .A2(G227), .ZN(n559) );
  XNOR2_X1 U667 ( .A(n559), .B(G140), .ZN(n560) );
  XNOR2_X1 U668 ( .A(n560), .B(n582), .ZN(n561) );
  XNOR2_X1 U669 ( .A(n562), .B(n561), .ZN(n563) );
  OR2_X2 U670 ( .A1(n775), .A2(G902), .ZN(n565) );
  XNOR2_X1 U671 ( .A(KEYINPUT74), .B(G469), .ZN(n564) );
  XNOR2_X2 U672 ( .A(n565), .B(n564), .ZN(n635) );
  NAND2_X1 U673 ( .A1(n566), .A2(G210), .ZN(n567) );
  XNOR2_X1 U674 ( .A(n568), .B(n567), .ZN(n571) );
  XNOR2_X1 U675 ( .A(n569), .B(G137), .ZN(n570) );
  XNOR2_X1 U676 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U677 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U678 ( .A(n575), .B(n574), .ZN(n756) );
  INV_X1 U679 ( .A(G472), .ZN(n754) );
  XNOR2_X1 U680 ( .A(n799), .B(KEYINPUT6), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n576), .A2(G221), .ZN(n581) );
  XNOR2_X1 U682 ( .A(G119), .B(G128), .ZN(n578) );
  XNOR2_X1 U683 ( .A(n581), .B(n580), .ZN(n585) );
  INV_X1 U684 ( .A(n582), .ZN(n583) );
  XNOR2_X1 U685 ( .A(n584), .B(n583), .ZN(n684) );
  INV_X1 U686 ( .A(G217), .ZN(n739) );
  XNOR2_X1 U687 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n587) );
  XNOR2_X1 U688 ( .A(n587), .B(KEYINPUT81), .ZN(n589) );
  XNOR2_X1 U689 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n588) );
  XNOR2_X1 U690 ( .A(n589), .B(n588), .ZN(n590) );
  AND2_X1 U691 ( .A1(n634), .A2(n599), .ZN(n592) );
  NAND2_X1 U692 ( .A1(n368), .A2(n592), .ZN(n712) );
  XNOR2_X1 U693 ( .A(n712), .B(G101), .ZN(G3) );
  NAND2_X1 U694 ( .A1(n593), .A2(n599), .ZN(n594) );
  OR2_X1 U695 ( .A1(n595), .A2(n594), .ZN(n598) );
  XNOR2_X1 U696 ( .A(KEYINPUT84), .B(KEYINPUT32), .ZN(n596) );
  XNOR2_X1 U697 ( .A(n596), .B(KEYINPUT66), .ZN(n597) );
  XNOR2_X1 U698 ( .A(n598), .B(n597), .ZN(n697) );
  XNOR2_X1 U699 ( .A(n697), .B(G119), .ZN(G21) );
  INV_X1 U700 ( .A(n599), .ZN(n699) );
  INV_X1 U701 ( .A(n647), .ZN(n600) );
  NAND2_X1 U702 ( .A1(n600), .A2(n646), .ZN(n602) );
  INV_X1 U703 ( .A(KEYINPUT101), .ZN(n601) );
  XNOR2_X1 U704 ( .A(n602), .B(n601), .ZN(n834) );
  INV_X1 U705 ( .A(n796), .ZN(n633) );
  NOR2_X1 U706 ( .A1(G900), .A2(n603), .ZN(n604) );
  AND2_X1 U707 ( .A1(n604), .A2(n822), .ZN(n606) );
  INV_X1 U708 ( .A(KEYINPUT106), .ZN(n605) );
  XNOR2_X1 U709 ( .A(n606), .B(n605), .ZN(n610) );
  INV_X1 U710 ( .A(n607), .ZN(n608) );
  NAND2_X1 U711 ( .A1(n822), .A2(n608), .ZN(n609) );
  NAND2_X1 U712 ( .A1(n610), .A2(n609), .ZN(n636) );
  AND2_X1 U713 ( .A1(n633), .A2(n636), .ZN(n611) );
  NOR2_X1 U714 ( .A1(n834), .A2(n623), .ZN(n612) );
  AND2_X1 U715 ( .A1(n699), .A2(n612), .ZN(n674) );
  INV_X1 U716 ( .A(n674), .ZN(n614) );
  OR2_X1 U717 ( .A1(n382), .A2(n640), .ZN(n613) );
  OR2_X1 U718 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U719 ( .A(n615), .B(KEYINPUT43), .ZN(n619) );
  XNOR2_X1 U720 ( .A(n616), .B(n617), .ZN(n649) );
  INV_X1 U721 ( .A(n649), .ZN(n618) );
  NAND2_X1 U722 ( .A1(n619), .A2(n618), .ZN(n680) );
  XNOR2_X1 U723 ( .A(n680), .B(G140), .ZN(G42) );
  XNOR2_X1 U724 ( .A(n649), .B(KEYINPUT38), .ZN(n807) );
  INV_X1 U725 ( .A(KEYINPUT111), .ZN(n620) );
  XNOR2_X1 U726 ( .A(n621), .B(n620), .ZN(n812) );
  OR2_X1 U727 ( .A1(n812), .A2(n811), .ZN(n622) );
  INV_X1 U728 ( .A(n635), .ZN(n624) );
  INV_X1 U729 ( .A(KEYINPUT110), .ZN(n625) );
  NAND2_X1 U730 ( .A1(n805), .A2(n628), .ZN(n627) );
  XNOR2_X1 U731 ( .A(n627), .B(KEYINPUT42), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(G137), .ZN(G39) );
  NOR2_X1 U733 ( .A1(n668), .A2(n834), .ZN(n629) );
  XOR2_X1 U734 ( .A(G146), .B(n629), .Z(G48) );
  XOR2_X1 U735 ( .A(G128), .B(KEYINPUT29), .Z(n632) );
  INV_X1 U736 ( .A(n646), .ZN(n630) );
  NAND2_X1 U737 ( .A1(n630), .A2(n647), .ZN(n837) );
  NOR2_X1 U738 ( .A1(n668), .A2(n837), .ZN(n631) );
  XOR2_X1 U739 ( .A(n632), .B(n631), .Z(G30) );
  NAND2_X1 U740 ( .A1(n635), .A2(n654), .ZN(n707) );
  XNOR2_X1 U741 ( .A(n707), .B(KEYINPUT107), .ZN(n637) );
  NAND2_X1 U742 ( .A1(n637), .A2(n636), .ZN(n639) );
  OR2_X1 U743 ( .A1(n695), .A2(n640), .ZN(n642) );
  XNOR2_X1 U744 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n641) );
  XNOR2_X1 U745 ( .A(n642), .B(n641), .ZN(n643) );
  INV_X1 U746 ( .A(n643), .ZN(n644) );
  OR2_X1 U747 ( .A1(n647), .A2(n646), .ZN(n648) );
  INV_X1 U748 ( .A(n648), .ZN(n705) );
  AND2_X1 U749 ( .A1(n705), .A2(n649), .ZN(n650) );
  XNOR2_X1 U750 ( .A(n653), .B(KEYINPUT39), .ZN(n659) );
  XNOR2_X1 U751 ( .A(n837), .B(KEYINPUT102), .ZN(n663) );
  OR2_X1 U752 ( .A1(n659), .A2(n663), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n681), .B(G134), .ZN(G36) );
  BUF_X1 U754 ( .A(n655), .Z(n709) );
  INV_X1 U755 ( .A(n709), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n710), .A2(n837), .ZN(n657) );
  XOR2_X1 U757 ( .A(G116), .B(n657), .Z(G18) );
  NOR2_X1 U758 ( .A1(n710), .A2(n834), .ZN(n658) );
  XOR2_X1 U759 ( .A(G113), .B(n658), .Z(G15) );
  NAND2_X1 U760 ( .A1(n730), .A2(n660), .ZN(n662) );
  INV_X1 U761 ( .A(KEYINPUT85), .ZN(n669) );
  NAND2_X1 U762 ( .A1(n668), .A2(n669), .ZN(n665) );
  AND2_X1 U763 ( .A1(n663), .A2(n834), .ZN(n813) );
  INV_X1 U764 ( .A(KEYINPUT47), .ZN(n666) );
  NOR2_X1 U765 ( .A1(n813), .A2(n666), .ZN(n664) );
  NAND2_X1 U766 ( .A1(n669), .A2(n666), .ZN(n667) );
  INV_X1 U767 ( .A(n668), .ZN(n672) );
  OR2_X1 U768 ( .A1(n813), .A2(KEYINPUT47), .ZN(n670) );
  NAND2_X1 U769 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U770 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U771 ( .A(n675), .B(KEYINPUT36), .ZN(n677) );
  INV_X1 U772 ( .A(n382), .ZN(n793) );
  OR2_X1 U773 ( .A1(n677), .A2(n793), .ZN(n843) );
  INV_X1 U774 ( .A(KEYINPUT48), .ZN(n679) );
  AND2_X1 U775 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U776 ( .A(n683), .B(n684), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n736), .B(n686), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n685), .A2(n532), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n686), .B(G227), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n687), .A2(G900), .ZN(n688) );
  NAND2_X1 U781 ( .A1(n688), .A2(G953), .ZN(n689) );
  XNOR2_X1 U782 ( .A(n689), .B(KEYINPUT126), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(G72) );
  NAND2_X1 U784 ( .A1(n693), .A2(G953), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n692), .A2(n694), .ZN(n729) );
  INV_X1 U786 ( .A(n717), .ZN(n706) );
  XNOR2_X1 U787 ( .A(n698), .B(KEYINPUT105), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U789 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n701) );
  INV_X1 U790 ( .A(KEYINPUT34), .ZN(n704) );
  NOR2_X1 U791 ( .A1(n707), .A2(n799), .ZN(n708) );
  NAND2_X1 U792 ( .A1(n709), .A2(n708), .ZN(n838) );
  INV_X1 U793 ( .A(n813), .ZN(n711) );
  INV_X1 U794 ( .A(KEYINPUT44), .ZN(n714) );
  NAND2_X1 U795 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U796 ( .A(n716), .B(KEYINPUT69), .ZN(n719) );
  INV_X1 U797 ( .A(n717), .ZN(n718) );
  NAND2_X1 U798 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U800 ( .A1(n735), .A2(n532), .ZN(n727) );
  XOR2_X1 U801 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n724) );
  NAND2_X1 U802 ( .A1(G224), .A2(G953), .ZN(n723) );
  XNOR2_X1 U803 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U804 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U805 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U806 ( .A(n729), .B(n728), .Z(G69) );
  XNOR2_X1 U807 ( .A(G131), .B(KEYINPUT127), .ZN(n731) );
  XOR2_X1 U808 ( .A(n731), .B(n730), .Z(G33) );
  INV_X1 U809 ( .A(KEYINPUT124), .ZN(n744) );
  NOR2_X1 U810 ( .A1(n732), .A2(KEYINPUT2), .ZN(n734) );
  INV_X1 U811 ( .A(KEYINPUT2), .ZN(n781) );
  NAND2_X1 U812 ( .A1(n733), .A2(n781), .ZN(n789) );
  NAND2_X1 U813 ( .A1(n737), .A2(KEYINPUT87), .ZN(n738) );
  NOR2_X1 U814 ( .A1(n774), .A2(n739), .ZN(n741) );
  XNOR2_X1 U815 ( .A(n741), .B(n740), .ZN(n743) );
  INV_X1 U816 ( .A(G952), .ZN(n742) );
  INV_X1 U817 ( .A(G210), .ZN(n745) );
  XNOR2_X1 U818 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n746) );
  XOR2_X1 U819 ( .A(n746), .B(KEYINPUT55), .Z(n747) );
  NAND2_X1 U820 ( .A1(n749), .A2(n770), .ZN(n752) );
  XOR2_X1 U821 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n750) );
  XNOR2_X1 U822 ( .A(n750), .B(KEYINPUT88), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n752), .B(n751), .ZN(G51) );
  XOR2_X1 U824 ( .A(G122), .B(n753), .Z(G24) );
  NOR2_X1 U825 ( .A1(n774), .A2(n754), .ZN(n758) );
  XNOR2_X1 U826 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U828 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U829 ( .A1(n759), .A2(n770), .ZN(n760) );
  XNOR2_X1 U830 ( .A(n760), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U831 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U832 ( .A(n764), .B(n763), .ZN(n765) );
  INV_X1 U833 ( .A(n770), .ZN(n779) );
  NOR2_X1 U834 ( .A1(n765), .A2(n779), .ZN(G63) );
  NOR2_X1 U835 ( .A1(n774), .A2(n766), .ZN(n769) );
  XNOR2_X1 U836 ( .A(n769), .B(n768), .ZN(n771) );
  NAND2_X1 U837 ( .A1(n771), .A2(n770), .ZN(n773) );
  XOR2_X1 U838 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n772) );
  XNOR2_X1 U839 ( .A(n773), .B(n772), .ZN(G60) );
  XNOR2_X1 U840 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n776) );
  XNOR2_X1 U841 ( .A(n776), .B(KEYINPUT58), .ZN(n777) );
  XNOR2_X1 U842 ( .A(n775), .B(n777), .ZN(n778) );
  NAND2_X1 U843 ( .A1(n781), .A2(KEYINPUT86), .ZN(n782) );
  NAND2_X1 U844 ( .A1(n780), .A2(n782), .ZN(n786) );
  AND2_X1 U845 ( .A1(n783), .A2(KEYINPUT86), .ZN(n784) );
  NAND2_X1 U846 ( .A1(n735), .A2(n784), .ZN(n785) );
  NAND2_X1 U847 ( .A1(n786), .A2(n785), .ZN(n791) );
  INV_X1 U848 ( .A(KEYINPUT86), .ZN(n787) );
  NAND2_X1 U849 ( .A1(n787), .A2(KEYINPUT2), .ZN(n788) );
  AND2_X1 U850 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U851 ( .A1(n791), .A2(n790), .ZN(n831) );
  NAND2_X1 U852 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U853 ( .A(n794), .B(KEYINPUT116), .ZN(n795) );
  XNOR2_X1 U854 ( .A(KEYINPUT50), .B(n795), .ZN(n801) );
  XNOR2_X1 U855 ( .A(n797), .B(KEYINPUT49), .ZN(n798) );
  NOR2_X1 U856 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U857 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U858 ( .A(KEYINPUT117), .B(n802), .Z(n803) );
  XNOR2_X1 U859 ( .A(n804), .B(KEYINPUT51), .ZN(n806) );
  INV_X1 U860 ( .A(n805), .ZN(n826) );
  NOR2_X1 U861 ( .A1(n806), .A2(n826), .ZN(n819) );
  NOR2_X1 U862 ( .A1(n351), .A2(n808), .ZN(n809) );
  XNOR2_X1 U863 ( .A(n809), .B(KEYINPUT118), .ZN(n810) );
  NOR2_X1 U864 ( .A1(n811), .A2(n810), .ZN(n815) );
  NOR2_X1 U865 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U866 ( .A1(n815), .A2(n814), .ZN(n817) );
  NOR2_X1 U867 ( .A1(n817), .A2(n381), .ZN(n818) );
  NOR2_X1 U868 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U869 ( .A(n820), .B(KEYINPUT52), .ZN(n821) );
  XNOR2_X1 U870 ( .A(n821), .B(KEYINPUT119), .ZN(n824) );
  AND2_X1 U871 ( .A1(n822), .A2(G952), .ZN(n823) );
  NAND2_X1 U872 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U873 ( .A1(n825), .A2(n532), .ZN(n829) );
  NOR2_X1 U874 ( .A1(n381), .A2(n826), .ZN(n827) );
  XNOR2_X1 U875 ( .A(n827), .B(KEYINPUT120), .ZN(n828) );
  NOR2_X1 U876 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U877 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U878 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n832) );
  XNOR2_X1 U879 ( .A(n833), .B(n832), .ZN(G75) );
  XOR2_X1 U880 ( .A(G104), .B(KEYINPUT113), .Z(n836) );
  OR2_X1 U881 ( .A1(n838), .A2(n834), .ZN(n835) );
  XNOR2_X1 U882 ( .A(n836), .B(n835), .ZN(G6) );
  XNOR2_X1 U883 ( .A(G107), .B(KEYINPUT27), .ZN(n842) );
  XOR2_X1 U884 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n840) );
  OR2_X1 U885 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U886 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U887 ( .A(n842), .B(n841), .ZN(G9) );
  XOR2_X1 U888 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n845) );
  XOR2_X1 U889 ( .A(G125), .B(n843), .Z(n844) );
  XNOR2_X1 U890 ( .A(n845), .B(n844), .ZN(G27) );
endmodule

