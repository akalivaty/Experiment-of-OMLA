

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742;

  NAND2_X1 U379 ( .A1(n570), .A2(n590), .ZN(n656) );
  NOR2_X1 U380 ( .A1(n547), .A2(n546), .ZN(n634) );
  NOR2_X1 U381 ( .A1(n656), .A2(n655), .ZN(n596) );
  XNOR2_X2 U382 ( .A(n527), .B(n433), .ZN(n655) );
  XNOR2_X2 U383 ( .A(G119), .B(KEYINPUT71), .ZN(n468) );
  NAND2_X1 U384 ( .A1(n741), .A2(n739), .ZN(n431) );
  XNOR2_X2 U385 ( .A(n572), .B(KEYINPUT22), .ZN(n583) );
  NOR2_X2 U386 ( .A1(G902), .A2(n695), .ZN(n520) );
  INV_X8 U387 ( .A(G953), .ZN(n728) );
  NOR2_X1 U388 ( .A1(n737), .A2(n626), .ZN(n429) );
  XNOR2_X1 U389 ( .A(n432), .B(n366), .ZN(n741) );
  XNOR2_X1 U390 ( .A(n445), .B(G478), .ZN(n546) );
  XNOR2_X1 U391 ( .A(n726), .B(n476), .ZN(n516) );
  XNOR2_X1 U392 ( .A(n434), .B(n710), .ZN(n515) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n479) );
  XNOR2_X1 U394 ( .A(n399), .B(n398), .ZN(n478) );
  XNOR2_X1 U395 ( .A(n468), .B(n400), .ZN(n399) );
  XNOR2_X1 U396 ( .A(G137), .B(G140), .ZN(n512) );
  XNOR2_X1 U397 ( .A(n518), .B(G469), .ZN(n519) );
  NOR2_X1 U398 ( .A1(n617), .A2(G902), .ZN(n485) );
  XNOR2_X1 U399 ( .A(n723), .B(n454), .ZN(n455) );
  XOR2_X1 U400 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n460) );
  XNOR2_X1 U401 ( .A(n410), .B(G101), .ZN(n477) );
  INV_X1 U402 ( .A(KEYINPUT67), .ZN(n410) );
  XNOR2_X1 U403 ( .A(n467), .B(G113), .ZN(n398) );
  XNOR2_X1 U404 ( .A(n476), .B(G125), .ZN(n463) );
  NAND2_X1 U405 ( .A1(n387), .A2(n386), .ZN(n388) );
  INV_X1 U406 ( .A(n639), .ZN(n389) );
  XNOR2_X1 U407 ( .A(n378), .B(n516), .ZN(n617) );
  XNOR2_X1 U408 ( .A(n484), .B(n420), .ZN(n378) );
  INV_X1 U409 ( .A(n477), .ZN(n420) );
  XNOR2_X1 U410 ( .A(n483), .B(n375), .ZN(n484) );
  XNOR2_X1 U411 ( .A(n463), .B(n401), .ZN(n723) );
  XNOR2_X1 U412 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n401) );
  XNOR2_X1 U413 ( .A(G119), .B(KEYINPUT24), .ZN(n491) );
  XOR2_X1 U414 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n441) );
  XNOR2_X1 U415 ( .A(n514), .B(n515), .ZN(n517) );
  XNOR2_X1 U416 ( .A(n724), .B(n513), .ZN(n514) );
  AND2_X1 U417 ( .A1(G227), .A2(n728), .ZN(n513) );
  XNOR2_X1 U418 ( .A(n374), .B(n470), .ZN(n693) );
  XNOR2_X1 U419 ( .A(n417), .B(n377), .ZN(n470) );
  XNOR2_X1 U420 ( .A(n709), .B(n515), .ZN(n374) );
  XNOR2_X1 U421 ( .A(n380), .B(n463), .ZN(n417) );
  NOR2_X1 U422 ( .A1(n671), .A2(n674), .ZN(n473) );
  AND2_X1 U423 ( .A1(n574), .A2(n533), .ZN(n534) );
  AND2_X1 U424 ( .A1(n650), .A2(n598), .ZN(n379) );
  INV_X1 U425 ( .A(KEYINPUT1), .ZN(n433) );
  NOR2_X1 U426 ( .A1(n421), .A2(n526), .ZN(n428) );
  XNOR2_X1 U427 ( .A(n505), .B(n504), .ZN(n652) );
  XNOR2_X1 U428 ( .A(n503), .B(n502), .ZN(n504) );
  INV_X1 U429 ( .A(KEYINPUT25), .ZN(n502) );
  NAND2_X1 U430 ( .A1(n700), .A2(G472), .ZN(n385) );
  XNOR2_X1 U431 ( .A(n416), .B(n367), .ZN(n415) );
  NAND2_X1 U432 ( .A1(n700), .A2(G475), .ZN(n416) );
  XNOR2_X1 U433 ( .A(G143), .B(G128), .ZN(n461) );
  XNOR2_X1 U434 ( .A(G113), .B(G131), .ZN(n452) );
  XOR2_X1 U435 ( .A(G104), .B(G143), .Z(n453) );
  XNOR2_X1 U436 ( .A(G122), .B(G140), .ZN(n448) );
  XNOR2_X1 U437 ( .A(n482), .B(n376), .ZN(n375) );
  INV_X1 U438 ( .A(KEYINPUT5), .ZN(n376) );
  XOR2_X1 U439 ( .A(G137), .B(KEYINPUT99), .Z(n481) );
  XNOR2_X1 U440 ( .A(n475), .B(n474), .ZN(n726) );
  XOR2_X1 U441 ( .A(G131), .B(KEYINPUT4), .Z(n474) );
  XNOR2_X1 U442 ( .A(n461), .B(G134), .ZN(n475) );
  XNOR2_X1 U443 ( .A(n461), .B(n418), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n462), .B(KEYINPUT4), .ZN(n418) );
  INV_X1 U445 ( .A(KEYINPUT77), .ZN(n462) );
  XNOR2_X1 U446 ( .A(n477), .B(KEYINPUT72), .ZN(n434) );
  XNOR2_X1 U447 ( .A(n464), .B(n465), .ZN(n377) );
  XNOR2_X1 U448 ( .A(KEYINPUT92), .B(KEYINPUT76), .ZN(n459) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n488) );
  XNOR2_X1 U450 ( .A(n597), .B(n419), .ZN(n574) );
  INV_X1 U451 ( .A(KEYINPUT6), .ZN(n419) );
  XNOR2_X1 U452 ( .A(n478), .B(n469), .ZN(n709) );
  XNOR2_X1 U453 ( .A(n466), .B(G107), .ZN(n710) );
  XNOR2_X1 U454 ( .A(G104), .B(G110), .ZN(n466) );
  XNOR2_X1 U455 ( .A(G116), .B(G107), .ZN(n436) );
  NAND2_X1 U456 ( .A1(n393), .A2(n392), .ZN(n613) );
  NAND2_X1 U457 ( .A1(n396), .A2(n394), .ZN(n393) );
  NAND2_X1 U458 ( .A1(n388), .A2(n364), .ZN(n392) );
  NAND2_X1 U459 ( .A1(n391), .A2(n390), .ZN(n612) );
  XNOR2_X1 U460 ( .A(n531), .B(n530), .ZN(n607) );
  INV_X1 U461 ( .A(KEYINPUT39), .ZN(n530) );
  NOR2_X1 U462 ( .A1(n541), .A2(n529), .ZN(n531) );
  NAND2_X1 U463 ( .A1(n424), .A2(n422), .ZN(n593) );
  AND2_X1 U464 ( .A1(n426), .A2(n423), .ZN(n422) );
  XNOR2_X1 U465 ( .A(n457), .B(n458), .ZN(n547) );
  XNOR2_X1 U466 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U467 ( .A(n524), .B(n523), .ZN(n739) );
  XNOR2_X1 U468 ( .A(n522), .B(KEYINPUT108), .ZN(n523) );
  XNOR2_X1 U469 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U470 ( .A(n582), .B(n581), .ZN(n737) );
  XNOR2_X1 U471 ( .A(n580), .B(KEYINPUT85), .ZN(n581) );
  INV_X1 U472 ( .A(KEYINPUT35), .ZN(n580) );
  AND2_X1 U473 ( .A1(n584), .A2(n362), .ZN(n626) );
  NAND2_X1 U474 ( .A1(n384), .A2(n414), .ZN(n383) );
  XNOR2_X1 U475 ( .A(n385), .B(n618), .ZN(n384) );
  NAND2_X1 U476 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U477 ( .A(KEYINPUT118), .ZN(n406) );
  INV_X1 U478 ( .A(KEYINPUT56), .ZN(n402) );
  AND2_X1 U479 ( .A1(n381), .A2(n552), .ZN(n357) );
  AND2_X1 U480 ( .A1(n411), .A2(n639), .ZN(n358) );
  AND2_X1 U481 ( .A1(G210), .A2(n472), .ZN(n359) );
  AND2_X1 U482 ( .A1(n638), .A2(n630), .ZN(n360) );
  AND2_X1 U483 ( .A1(n547), .A2(n546), .ZN(n361) );
  AND2_X1 U484 ( .A1(n658), .A2(n652), .ZN(n362) );
  OR2_X1 U485 ( .A1(n389), .A2(n555), .ZN(n363) );
  INV_X1 U486 ( .A(G146), .ZN(n476) );
  AND2_X1 U487 ( .A1(n358), .A2(n555), .ZN(n364) );
  INV_X1 U488 ( .A(n411), .ZN(n641) );
  XOR2_X1 U489 ( .A(G472), .B(KEYINPUT74), .Z(n365) );
  XOR2_X1 U490 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n366) );
  XOR2_X1 U491 ( .A(n698), .B(n697), .Z(n367) );
  XOR2_X1 U492 ( .A(n695), .B(n694), .Z(n368) );
  XOR2_X1 U493 ( .A(n693), .B(n435), .Z(n369) );
  XNOR2_X1 U494 ( .A(KEYINPUT46), .B(KEYINPUT86), .ZN(n370) );
  XOR2_X1 U495 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n371) );
  NOR2_X1 U496 ( .A1(G952), .A2(n728), .ZN(n708) );
  INV_X1 U497 ( .A(n708), .ZN(n414) );
  XOR2_X1 U498 ( .A(KEYINPUT63), .B(KEYINPUT109), .Z(n372) );
  XOR2_X1 U499 ( .A(n699), .B(KEYINPUT60), .Z(n373) );
  XNOR2_X1 U500 ( .A(n413), .B(n373), .ZN(G60) );
  NAND2_X1 U501 ( .A1(n587), .A2(n573), .ZN(n430) );
  NAND2_X1 U502 ( .A1(n593), .A2(n428), .ZN(n541) );
  XNOR2_X1 U503 ( .A(n379), .B(KEYINPUT34), .ZN(n579) );
  NAND2_X1 U504 ( .A1(n738), .A2(n429), .ZN(n586) );
  XNOR2_X2 U505 ( .A(n430), .B(KEYINPUT32), .ZN(n738) );
  INV_X1 U506 ( .A(n412), .ZN(n535) );
  NAND2_X1 U507 ( .A1(n412), .A2(n668), .ZN(n544) );
  XNOR2_X2 U508 ( .A(n471), .B(n359), .ZN(n412) );
  XNOR2_X1 U509 ( .A(n382), .B(KEYINPUT75), .ZN(n381) );
  AND2_X1 U510 ( .A1(n549), .A2(n631), .ZN(n382) );
  XNOR2_X1 U511 ( .A(n383), .B(n372), .ZN(G57) );
  NOR2_X1 U512 ( .A1(n634), .A2(n361), .ZN(n548) );
  NOR2_X1 U513 ( .A1(n554), .A2(n363), .ZN(n394) );
  INV_X1 U514 ( .A(n554), .ZN(n386) );
  INV_X1 U515 ( .A(n553), .ZN(n387) );
  AND2_X1 U516 ( .A1(n388), .A2(n555), .ZN(n395) );
  NOR2_X1 U517 ( .A1(n554), .A2(n555), .ZN(n397) );
  NAND2_X1 U518 ( .A1(n395), .A2(n411), .ZN(n390) );
  NAND2_X1 U519 ( .A1(n396), .A2(n397), .ZN(n391) );
  NOR2_X1 U520 ( .A1(n553), .A2(n641), .ZN(n396) );
  XNOR2_X2 U521 ( .A(G116), .B(KEYINPUT91), .ZN(n400) );
  XNOR2_X1 U522 ( .A(n403), .B(n402), .ZN(G51) );
  NAND2_X1 U523 ( .A1(n404), .A2(n414), .ZN(n403) );
  XNOR2_X1 U524 ( .A(n405), .B(n369), .ZN(n404) );
  NAND2_X1 U525 ( .A1(n700), .A2(G210), .ZN(n405) );
  XNOR2_X1 U526 ( .A(n407), .B(n406), .ZN(G54) );
  NAND2_X1 U527 ( .A1(n408), .A2(n414), .ZN(n407) );
  XNOR2_X1 U528 ( .A(n409), .B(n368), .ZN(n408) );
  NAND2_X1 U529 ( .A1(n700), .A2(G469), .ZN(n409) );
  XNOR2_X1 U530 ( .A(n535), .B(KEYINPUT38), .ZN(n669) );
  NAND2_X1 U531 ( .A1(n542), .A2(n412), .ZN(n630) );
  OR2_X1 U532 ( .A1(n559), .A2(n412), .ZN(n411) );
  INV_X1 U533 ( .A(n597), .ZN(n658) );
  XNOR2_X1 U534 ( .A(n525), .B(KEYINPUT30), .ZN(n421) );
  NAND2_X1 U535 ( .A1(n656), .A2(n427), .ZN(n423) );
  NAND2_X1 U536 ( .A1(n425), .A2(n527), .ZN(n424) );
  NOR2_X1 U537 ( .A1(n656), .A2(n427), .ZN(n425) );
  NAND2_X1 U538 ( .A1(n528), .A2(n427), .ZN(n426) );
  INV_X1 U539 ( .A(KEYINPUT98), .ZN(n427) );
  NOR2_X2 U540 ( .A1(n583), .A2(n574), .ZN(n587) );
  XNOR2_X2 U541 ( .A(n431), .B(n370), .ZN(n554) );
  NAND2_X1 U542 ( .A1(n607), .A2(n361), .ZN(n432) );
  XNOR2_X2 U543 ( .A(n520), .B(n519), .ZN(n527) );
  XNOR2_X1 U544 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n435) );
  INV_X1 U545 ( .A(KEYINPUT48), .ZN(n555) );
  AND2_X1 U546 ( .A1(n532), .A2(n361), .ZN(n533) );
  XNOR2_X1 U547 ( .A(KEYINPUT16), .B(G122), .ZN(n469) );
  XNOR2_X1 U548 ( .A(n723), .B(n495), .ZN(n498) );
  XNOR2_X1 U549 ( .A(KEYINPUT36), .B(KEYINPUT88), .ZN(n536) );
  XOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .Z(n611) );
  XNOR2_X1 U551 ( .A(n436), .B(KEYINPUT7), .ZN(n437) );
  XOR2_X1 U552 ( .A(n437), .B(KEYINPUT9), .Z(n439) );
  XNOR2_X1 U553 ( .A(n475), .B(G122), .ZN(n438) );
  XNOR2_X1 U554 ( .A(n439), .B(n438), .ZN(n444) );
  NAND2_X1 U555 ( .A1(G234), .A2(n728), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U557 ( .A(KEYINPUT81), .B(n442), .Z(n496) );
  NAND2_X1 U558 ( .A1(G217), .A2(n496), .ZN(n443) );
  XOR2_X1 U559 ( .A(n444), .B(n443), .Z(n702) );
  NOR2_X1 U560 ( .A1(G902), .A2(n702), .ZN(n445) );
  INV_X1 U561 ( .A(n546), .ZN(n539) );
  XNOR2_X1 U562 ( .A(KEYINPUT13), .B(G475), .ZN(n458) );
  XOR2_X1 U563 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n447) );
  NAND2_X1 U564 ( .A1(G214), .A2(n479), .ZN(n446) );
  XNOR2_X1 U565 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U566 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n449) );
  XNOR2_X1 U567 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U568 ( .A(n451), .B(n450), .Z(n456) );
  XNOR2_X1 U569 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U570 ( .A(n456), .B(n455), .ZN(n696) );
  NOR2_X1 U571 ( .A1(G902), .A2(n696), .ZN(n457) );
  OR2_X1 U572 ( .A1(n539), .A2(n547), .ZN(n671) );
  XNOR2_X1 U573 ( .A(n460), .B(n459), .ZN(n464) );
  NAND2_X1 U574 ( .A1(G224), .A2(n728), .ZN(n465) );
  INV_X1 U575 ( .A(KEYINPUT3), .ZN(n467) );
  INV_X1 U576 ( .A(n611), .ZN(n499) );
  NAND2_X1 U577 ( .A1(n693), .A2(n499), .ZN(n471) );
  OR2_X1 U578 ( .A1(G237), .A2(G902), .ZN(n472) );
  NAND2_X1 U579 ( .A1(G214), .A2(n472), .ZN(n668) );
  NAND2_X1 U580 ( .A1(n669), .A2(n668), .ZN(n674) );
  XNOR2_X1 U581 ( .A(n473), .B(KEYINPUT41), .ZN(n667) );
  INV_X1 U582 ( .A(n478), .ZN(n483) );
  NAND2_X1 U583 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U584 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X2 U585 ( .A(n485), .B(n365), .ZN(n597) );
  NOR2_X1 U586 ( .A1(G900), .A2(n728), .ZN(n486) );
  NAND2_X1 U587 ( .A1(n486), .A2(G902), .ZN(n487) );
  NAND2_X1 U588 ( .A1(G952), .A2(n728), .ZN(n561) );
  NAND2_X1 U589 ( .A1(n487), .A2(n561), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n488), .B(KEYINPUT14), .ZN(n563) );
  NAND2_X1 U591 ( .A1(n489), .A2(n563), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G128), .B(G110), .ZN(n490) );
  XNOR2_X1 U593 ( .A(n490), .B(n512), .ZN(n494) );
  XOR2_X1 U594 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n492) );
  XNOR2_X1 U595 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U596 ( .A1(n496), .A2(G221), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n498), .B(n497), .ZN(n704) );
  NOR2_X1 U598 ( .A1(G902), .A2(n704), .ZN(n505) );
  NAND2_X1 U599 ( .A1(n499), .A2(G234), .ZN(n501) );
  XNOR2_X1 U600 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n500) );
  XNOR2_X1 U601 ( .A(n501), .B(n500), .ZN(n506) );
  NAND2_X1 U602 ( .A1(G217), .A2(n506), .ZN(n503) );
  NAND2_X1 U603 ( .A1(n506), .A2(G221), .ZN(n507) );
  XNOR2_X1 U604 ( .A(n507), .B(KEYINPUT21), .ZN(n508) );
  XNOR2_X1 U605 ( .A(KEYINPUT97), .B(n508), .ZN(n570) );
  NAND2_X1 U606 ( .A1(n652), .A2(n570), .ZN(n509) );
  NOR2_X1 U607 ( .A1(n526), .A2(n509), .ZN(n532) );
  AND2_X1 U608 ( .A1(n597), .A2(n532), .ZN(n511) );
  XNOR2_X1 U609 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n510) );
  XNOR2_X1 U610 ( .A(n511), .B(n510), .ZN(n521) );
  XNOR2_X1 U611 ( .A(KEYINPUT94), .B(n512), .ZN(n724) );
  XNOR2_X1 U612 ( .A(n517), .B(n516), .ZN(n695) );
  INV_X1 U613 ( .A(KEYINPUT70), .ZN(n518) );
  NAND2_X1 U614 ( .A1(n521), .A2(n527), .ZN(n545) );
  NOR2_X1 U615 ( .A1(n667), .A2(n545), .ZN(n524) );
  INV_X1 U616 ( .A(KEYINPUT42), .ZN(n522) );
  NAND2_X1 U617 ( .A1(n597), .A2(n668), .ZN(n525) );
  INV_X1 U618 ( .A(n652), .ZN(n590) );
  INV_X1 U619 ( .A(n527), .ZN(n528) );
  INV_X1 U620 ( .A(n669), .ZN(n529) );
  NAND2_X1 U621 ( .A1(n534), .A2(n668), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n556), .A2(n535), .ZN(n537) );
  INV_X1 U623 ( .A(n655), .ZN(n589) );
  NAND2_X1 U624 ( .A1(n538), .A2(n589), .ZN(n638) );
  NAND2_X1 U625 ( .A1(n547), .A2(n539), .ZN(n540) );
  XNOR2_X1 U626 ( .A(n540), .B(KEYINPUT104), .ZN(n577) );
  NOR2_X1 U627 ( .A1(n577), .A2(n541), .ZN(n542) );
  INV_X1 U628 ( .A(KEYINPUT19), .ZN(n543) );
  XNOR2_X1 U629 ( .A(n544), .B(n543), .ZN(n566) );
  NOR2_X1 U630 ( .A1(n545), .A2(n566), .ZN(n631) );
  XNOR2_X1 U631 ( .A(n548), .B(KEYINPUT102), .ZN(n673) );
  XNOR2_X1 U632 ( .A(KEYINPUT80), .B(n673), .ZN(n601) );
  NOR2_X1 U633 ( .A1(KEYINPUT47), .A2(n601), .ZN(n549) );
  INV_X1 U634 ( .A(n673), .ZN(n550) );
  NAND2_X1 U635 ( .A1(n550), .A2(n631), .ZN(n551) );
  NAND2_X1 U636 ( .A1(n551), .A2(KEYINPUT47), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n360), .A2(n357), .ZN(n553) );
  XOR2_X1 U638 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n558) );
  NOR2_X1 U639 ( .A1(n556), .A2(n589), .ZN(n557) );
  XNOR2_X1 U640 ( .A(n558), .B(n557), .ZN(n559) );
  NOR2_X1 U641 ( .A1(G898), .A2(n728), .ZN(n560) );
  XOR2_X1 U642 ( .A(KEYINPUT93), .B(n560), .Z(n713) );
  NAND2_X1 U643 ( .A1(n713), .A2(G902), .ZN(n562) );
  AND2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n564) );
  INV_X1 U645 ( .A(n563), .ZN(n684) );
  OR2_X1 U646 ( .A1(n564), .A2(n684), .ZN(n565) );
  NOR2_X2 U647 ( .A1(n566), .A2(n565), .ZN(n569) );
  XOR2_X1 U648 ( .A(KEYINPUT0), .B(KEYINPUT66), .Z(n567) );
  XNOR2_X1 U649 ( .A(KEYINPUT89), .B(n567), .ZN(n568) );
  XNOR2_X2 U650 ( .A(n569), .B(n568), .ZN(n598) );
  INV_X1 U651 ( .A(n570), .ZN(n651) );
  NOR2_X1 U652 ( .A1(n671), .A2(n651), .ZN(n571) );
  NAND2_X1 U653 ( .A1(n598), .A2(n571), .ZN(n572) );
  NOR2_X1 U654 ( .A1(n590), .A2(n655), .ZN(n573) );
  NAND2_X1 U655 ( .A1(n596), .A2(n574), .ZN(n576) );
  XOR2_X1 U656 ( .A(KEYINPUT103), .B(KEYINPUT33), .Z(n575) );
  XNOR2_X1 U657 ( .A(n576), .B(n575), .ZN(n650) );
  XOR2_X1 U658 ( .A(n577), .B(KEYINPUT78), .Z(n578) );
  NAND2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n582) );
  NOR2_X1 U660 ( .A1(n589), .A2(n583), .ZN(n584) );
  NOR2_X2 U661 ( .A1(n586), .A2(KEYINPUT73), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT44), .ZN(n605) );
  NAND2_X1 U663 ( .A1(n586), .A2(KEYINPUT73), .ZN(n592) );
  XNOR2_X1 U664 ( .A(KEYINPUT87), .B(n587), .ZN(n588) );
  NOR2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n619) );
  NAND2_X1 U667 ( .A1(n592), .A2(n619), .ZN(n603) );
  INV_X1 U668 ( .A(n593), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n658), .A2(n598), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n622) );
  AND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n664) );
  NAND2_X1 U672 ( .A1(n598), .A2(n664), .ZN(n599) );
  XNOR2_X1 U673 ( .A(KEYINPUT31), .B(n599), .ZN(n635) );
  NOR2_X1 U674 ( .A1(n622), .A2(n635), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X2 U678 ( .A(n606), .B(n371), .ZN(n646) );
  NAND2_X1 U679 ( .A1(n607), .A2(n634), .ZN(n639) );
  NAND2_X1 U680 ( .A1(KEYINPUT2), .A2(n639), .ZN(n608) );
  XOR2_X1 U681 ( .A(KEYINPUT79), .B(n608), .Z(n609) );
  NOR2_X1 U682 ( .A1(n646), .A2(n609), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n612), .A2(n610), .ZN(n645) );
  NAND2_X1 U684 ( .A1(n611), .A2(n645), .ZN(n616) );
  XNOR2_X2 U685 ( .A(n613), .B(KEYINPUT83), .ZN(n642) );
  NOR2_X1 U686 ( .A1(n642), .A2(n646), .ZN(n614) );
  NOR2_X1 U687 ( .A1(KEYINPUT2), .A2(n614), .ZN(n615) );
  NOR2_X4 U688 ( .A1(n616), .A2(n615), .ZN(n700) );
  XOR2_X1 U689 ( .A(KEYINPUT62), .B(n617), .Z(n618) );
  XNOR2_X1 U690 ( .A(G101), .B(n619), .ZN(G3) );
  NAND2_X1 U691 ( .A1(n622), .A2(n361), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n620), .B(KEYINPUT110), .ZN(n621) );
  XNOR2_X1 U693 ( .A(G104), .B(n621), .ZN(G6) );
  XOR2_X1 U694 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n624) );
  NAND2_X1 U695 ( .A1(n622), .A2(n634), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U697 ( .A(G107), .B(n625), .ZN(G9) );
  XOR2_X1 U698 ( .A(G110), .B(n626), .Z(G12) );
  XOR2_X1 U699 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n628) );
  NAND2_X1 U700 ( .A1(n631), .A2(n634), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XOR2_X1 U702 ( .A(G128), .B(n629), .Z(G30) );
  XNOR2_X1 U703 ( .A(G143), .B(n630), .ZN(G45) );
  NAND2_X1 U704 ( .A1(n631), .A2(n361), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(G146), .ZN(G48) );
  NAND2_X1 U706 ( .A1(n635), .A2(n361), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(G113), .ZN(G15) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(G116), .ZN(G18) );
  XOR2_X1 U710 ( .A(G125), .B(KEYINPUT37), .Z(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G27) );
  XNOR2_X1 U712 ( .A(G134), .B(KEYINPUT112), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(G36) );
  XOR2_X1 U714 ( .A(G140), .B(n641), .Z(G42) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n649) );
  INV_X1 U718 ( .A(n646), .ZN(n718) );
  NOR2_X1 U719 ( .A1(KEYINPUT2), .A2(n718), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n647), .B(KEYINPUT82), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n690) );
  INV_X1 U722 ( .A(n650), .ZN(n678) );
  OR2_X1 U723 ( .A1(n678), .A2(n667), .ZN(n687) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n654) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(n661) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT50), .B(n657), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT114), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(KEYINPUT51), .B(n665), .Z(n666) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n680) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT115), .B(n672), .Z(n676) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U742 ( .A(KEYINPUT52), .B(n681), .Z(n682) );
  XOR2_X1 U743 ( .A(KEYINPUT116), .B(n682), .Z(n683) );
  NOR2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n685), .A2(G952), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U747 ( .A(KEYINPUT117), .B(n688), .Z(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U749 ( .A1(n728), .A2(n691), .ZN(n692) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(n692), .Z(G75) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XOR2_X1 U752 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n698) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT90), .ZN(n697) );
  XNOR2_X1 U754 ( .A(KEYINPUT65), .B(KEYINPUT119), .ZN(n699) );
  NAND2_X1 U755 ( .A1(G478), .A2(n700), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U757 ( .A1(n708), .A2(n703), .ZN(G63) );
  XNOR2_X1 U758 ( .A(n704), .B(KEYINPUT120), .ZN(n706) );
  NAND2_X1 U759 ( .A1(G217), .A2(n700), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n708), .A2(n707), .ZN(G66) );
  XOR2_X1 U762 ( .A(KEYINPUT122), .B(n709), .Z(n712) );
  XNOR2_X1 U763 ( .A(G101), .B(n710), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n714) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n722) );
  XOR2_X1 U766 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n716) );
  NAND2_X1 U767 ( .A1(G224), .A2(G953), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(G898), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n718), .A2(n728), .ZN(n719) );
  NAND2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(G69) );
  XOR2_X1 U773 ( .A(n724), .B(n723), .Z(n725) );
  XOR2_X1 U774 ( .A(n726), .B(n725), .Z(n730) );
  XOR2_X1 U775 ( .A(n730), .B(KEYINPUT123), .Z(n727) );
  XNOR2_X1 U776 ( .A(n727), .B(n642), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n736) );
  XNOR2_X1 U778 ( .A(n730), .B(G227), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n731), .B(KEYINPUT124), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G900), .ZN(n733) );
  XOR2_X1 U781 ( .A(KEYINPUT125), .B(n733), .Z(n734) );
  NAND2_X1 U782 ( .A1(G953), .A2(n734), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U784 ( .A(n737), .B(G122), .Z(G24) );
  XNOR2_X1 U785 ( .A(n738), .B(G119), .ZN(G21) );
  XNOR2_X1 U786 ( .A(G137), .B(KEYINPUT126), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n740), .B(n739), .ZN(G39) );
  XOR2_X1 U788 ( .A(n741), .B(G131), .Z(n742) );
  XNOR2_X1 U789 ( .A(KEYINPUT127), .B(n742), .ZN(G33) );
endmodule

