//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(KEYINPUT68), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(KEYINPUT68), .B2(new_n457), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n461), .B2(new_n462), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n460), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n471), .A2(new_n479), .ZN(G160));
  AOI21_X1  g055(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT71), .Z(new_n483));
  AOI21_X1  g058(.A(new_n460), .B1(new_n472), .B2(new_n474), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT72), .Z(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n475), .A2(new_n476), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(new_n508), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n503), .A2(new_n510), .B1(new_n511), .B2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  INV_X1    g091(.A(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT74), .B1(new_n512), .B2(new_n513), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n524), .A2(new_n525), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n529), .B1(new_n509), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n520), .A2(new_n527), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n503), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n524), .A2(new_n525), .A3(G543), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n518), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n535), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n519), .A2(G81), .B1(new_n526), .B2(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n503), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND4_X1  g126(.A1(new_n524), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n526), .A2(new_n555), .A3(G53), .A4(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT77), .B1(new_n552), .B2(new_n556), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n552), .A2(new_n560), .A3(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n554), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n563), .A2(new_n503), .B1(new_n564), .B2(new_n518), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  OAI21_X1  g142(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n509), .A2(G87), .A3(new_n517), .ZN(new_n569));
  INV_X1    g144(.A(G49), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n537), .ZN(G288));
  NAND2_X1  g146(.A1(new_n509), .A2(G61), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n509), .A2(new_n574), .A3(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n503), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n509), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G48), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n514), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n519), .A2(G85), .B1(new_n526), .B2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n503), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n509), .A2(G66), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n592), .A2(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G286), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(G299), .B(KEYINPUT80), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G280));
  XNOR2_X1  g180(.A(KEYINPUT81), .B(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(G860), .B2(new_n606), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g185(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  NAND3_X1  g187(.A1(new_n475), .A2(new_n476), .A3(new_n465), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n481), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n460), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n484), .B(KEYINPUT72), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n619), .B1(new_n620), .B2(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n617), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n625), .A3(new_n626), .ZN(G156));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(G401));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT84), .Z(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n646), .B2(KEYINPUT85), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(KEYINPUT85), .B2(new_n646), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2084), .B(G2090), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n646), .B(KEYINPUT17), .Z(new_n650));
  INV_X1    g225(.A(new_n644), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n644), .A2(new_n649), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n666), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n670), .C1(new_n663), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(G171), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G5), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G1961), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT97), .Z(new_n684));
  NOR2_X1   g259(.A1(G29), .A2(G33), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT25), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n475), .A2(new_n476), .A3(G127), .ZN(new_n688));
  NAND2_X1  g263(.A1(G115), .A2(G2104), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n460), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g265(.A(new_n687), .B(new_n690), .C1(G139), .C2(new_n481), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n685), .B1(new_n691), .B2(G29), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(G2072), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT90), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n679), .A2(G4), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n598), .B2(new_n679), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1348), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(G2072), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  NOR4_X1   g274(.A1(new_n684), .A2(new_n694), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G2084), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(KEYINPUT24), .B2(G34), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(KEYINPUT24), .B2(G34), .ZN(new_n704));
  INV_X1    g279(.A(G160), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(G29), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n681), .A2(new_n682), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G21), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G168), .B2(G16), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G1966), .ZN(new_n710));
  NAND2_X1  g285(.A1(G162), .A2(G29), .ZN(new_n711));
  OR2_X1    g286(.A1(G29), .A2(G35), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT29), .B(G2090), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n702), .A2(G32), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n485), .A2(G129), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT92), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT94), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT26), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n717), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n707), .B(new_n716), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n715), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n713), .A2(new_n730), .B1(G1966), .B2(new_n709), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n702), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n485), .A2(G128), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(G116), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n481), .B2(G140), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2067), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n731), .B(new_n741), .C1(new_n701), .C2(new_n706), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n546), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT89), .B(G1341), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n702), .B1(new_n748), .B2(G28), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(KEYINPUT96), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(G28), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n749), .B2(KEYINPUT96), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n747), .B1(new_n750), .B2(new_n752), .C1(new_n624), .C2(new_n702), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  NAND2_X1  g329(.A1(G164), .A2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G27), .B2(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n746), .B(new_n757), .C1(new_n754), .C2(new_n756), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n729), .A2(new_n742), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n679), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n727), .A2(new_n728), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT95), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n700), .A2(new_n759), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G6), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n580), .B2(G16), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n679), .A2(G22), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G166), .B2(new_n679), .ZN(new_n775));
  INV_X1    g350(.A(G1971), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n679), .A2(G23), .ZN(new_n778));
  INV_X1    g353(.A(G288), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n679), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AND4_X1   g357(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT34), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n481), .A2(G131), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n460), .A2(G107), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n789));
  INV_X1    g364(.A(G119), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n787), .B1(new_n788), .B2(new_n789), .C1(new_n622), .C2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G25), .B(new_n791), .S(G29), .Z(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT35), .B(G1991), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT87), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n792), .B(new_n794), .Z(new_n795));
  INV_X1    g370(.A(G1986), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n679), .A2(G24), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G290), .B2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n796), .B2(new_n798), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n785), .A2(new_n786), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n785), .A2(new_n803), .A3(new_n786), .A4(new_n800), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n766), .B1(new_n802), .B2(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  NAND2_X1  g381(.A1(new_n598), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT38), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n503), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n518), .A2(new_n811), .B1(new_n537), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n546), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n814), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n545), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n808), .B(new_n818), .Z(new_n819));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n820));
  AOI21_X1  g395(.A(G860), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n691), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n726), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n721), .B(new_n725), .C1(new_n826), .C2(new_n691), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n739), .B(G164), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(G118), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(G2105), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n481), .B2(G142), .ZN(new_n839));
  INV_X1    g414(.A(G130), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n622), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n791), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n614), .B(KEYINPUT99), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n845), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n835), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n832), .A2(new_n848), .A3(new_n847), .A4(new_n834), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n489), .B(new_n705), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n624), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g437(.A(G288), .B(KEYINPUT103), .ZN(new_n863));
  XNOR2_X1  g438(.A(G305), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G290), .B(G303), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n867));
  XOR2_X1   g442(.A(new_n866), .B(new_n867), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n608), .B(new_n818), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n598), .B1(KEYINPUT102), .B2(G299), .ZN(new_n871));
  AND2_X1   g446(.A1(G299), .A2(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n871), .A2(new_n872), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(KEYINPUT41), .A3(new_n873), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n869), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n868), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n868), .B1(new_n882), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g459(.A(G868), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(G868), .B2(new_n814), .ZN(G295));
  OAI21_X1  g461(.A(new_n885), .B1(G868), .B2(new_n814), .ZN(G331));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n818), .A2(G301), .ZN(new_n889));
  OAI21_X1  g464(.A(G171), .B1(new_n815), .B2(new_n817), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n889), .A2(G168), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G168), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n878), .A3(new_n880), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n873), .B(new_n879), .C1(new_n891), .C2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n896), .B2(new_n866), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n898));
  INV_X1    g473(.A(new_n866), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n899), .A3(new_n895), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n898), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n888), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT44), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(G397));
  NAND2_X1  g483(.A1(new_n499), .A2(new_n501), .ZN(new_n909));
  INV_X1    g484(.A(new_n496), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT106), .B(G1384), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT107), .B1(G164), .B2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n477), .A2(new_n478), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G2105), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n463), .A2(new_n469), .A3(new_n466), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n469), .B1(new_n463), .B2(new_n466), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n923), .A3(G40), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT109), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(G1996), .A3(new_n726), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT110), .Z(new_n928));
  AND2_X1   g503(.A1(new_n791), .A2(new_n794), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n791), .A2(new_n794), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n739), .A2(G2067), .ZN(new_n933));
  INV_X1    g508(.A(G2067), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n734), .A2(new_n934), .A3(new_n738), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n926), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n925), .A2(G1996), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n721), .A3(new_n725), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n932), .B1(new_n926), .B2(new_n936), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n925), .ZN(new_n943));
  NOR2_X1   g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT48), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n928), .A2(new_n931), .A3(new_n942), .A4(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n938), .B(KEYINPUT46), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n926), .B1(new_n726), .B2(new_n936), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n947), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n926), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n928), .A2(new_n930), .A3(new_n942), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(new_n935), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT62), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n911), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT112), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n920), .A2(new_n923), .A3(G40), .A4(new_n701), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1966), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n471), .A2(new_n479), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n909), .B2(new_n910), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n917), .B1(G164), .B2(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n971), .A2(new_n973), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n963), .B1(new_n981), .B2(G168), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n911), .B2(new_n965), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n924), .ZN(new_n984));
  AOI21_X1  g559(.A(G1966), .B1(new_n984), .B2(new_n978), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n972), .B1(new_n969), .B2(new_n970), .ZN(new_n986));
  OAI21_X1  g561(.A(G286), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n962), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT51), .B(new_n963), .C1(new_n981), .C2(G168), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n988), .A2(KEYINPUT121), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT121), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n971), .A2(new_n973), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n980), .A2(new_n974), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(G168), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n987), .A3(G8), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT51), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n982), .A2(new_n962), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n961), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT121), .B1(new_n988), .B2(new_n989), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n991), .A3(new_n997), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n911), .A2(KEYINPUT45), .A3(new_n914), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n984), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n776), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n971), .A2(new_n976), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(G2090), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n509), .A2(G62), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G75), .A2(G543), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n503), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n1011));
  INV_X1    g586(.A(new_n508), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT73), .B1(new_n507), .B2(G543), .ZN(new_n1013));
  OAI211_X1 g588(.A(G88), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G50), .A2(G543), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n514), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT55), .B(G8), .C1(new_n1010), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(G303), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1020), .A3(KEYINPUT114), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1007), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n977), .A2(G40), .A3(new_n920), .A4(new_n923), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G288), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1032), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT115), .B(G1976), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n1029), .A3(new_n1036), .A4(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n576), .B2(new_n579), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n572), .A2(KEYINPUT78), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G73), .A2(G543), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n575), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G651), .ZN(new_n1043));
  INV_X1    g618(.A(new_n579), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1046), .A3(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT49), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1030), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1038), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n984), .B2(new_n1003), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n976), .A2(new_n967), .A3(new_n966), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2090), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1025), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1024), .A3(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1028), .A2(new_n1051), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1006), .A2(new_n682), .ZN(new_n1059));
  INV_X1    g634(.A(new_n980), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2078), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n976), .A2(new_n1003), .A3(new_n754), .A4(new_n979), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1060), .A2(new_n1062), .B1(new_n1063), .B2(new_n1061), .ZN(new_n1064));
  AOI21_X1  g639(.A(G301), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n999), .A2(new_n1002), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n558), .A2(new_n559), .ZN(new_n1069));
  INV_X1    g644(.A(new_n561), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n560), .B1(new_n552), .B2(KEYINPUT9), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n565), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1068), .B1(new_n1073), .B2(KEYINPUT116), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NAND3_X1  g650(.A1(G299), .A2(new_n1075), .A3(KEYINPUT57), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1053), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n976), .A2(new_n1003), .A3(new_n979), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n1029), .B2(G2067), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n976), .A2(new_n1084), .A3(new_n934), .A4(new_n977), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n924), .B1(new_n969), .B2(new_n970), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(G1348), .B2(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1088), .A2(KEYINPUT118), .A3(new_n598), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT118), .B1(new_n1088), .B2(new_n598), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(G299), .B2(new_n1075), .ZN(new_n1092));
  AOI211_X1 g667(.A(KEYINPUT116), .B(new_n1068), .C1(new_n562), .C2(new_n566), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1089), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1081), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1081), .B2(new_n1094), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1006), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n598), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1103), .A4(new_n1086), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n542), .B(new_n544), .C1(KEYINPUT119), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1996), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n976), .A2(new_n1003), .A3(new_n1107), .A4(new_n979), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1029), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT120), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1111), .B(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n598), .B1(new_n1088), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1086), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1104), .B(new_n1115), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1082), .A2(new_n1096), .B1(new_n1100), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n990), .A2(new_n998), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1059), .A2(G301), .A3(new_n1064), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n479), .A2(new_n975), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT123), .B1(new_n921), .B2(new_n922), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n468), .A2(new_n1128), .A3(new_n470), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT124), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1126), .A2(new_n1132), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1062), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G164), .A2(new_n913), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(KEYINPUT45), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1131), .A2(new_n918), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1063), .A2(new_n1061), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1137), .B(new_n1138), .C1(G1961), .C2(new_n1087), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1125), .B1(new_n1139), .B2(G171), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1059), .A2(new_n1064), .A3(KEYINPUT125), .A4(G301), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1124), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1143));
  NOR2_X1   g718(.A1(new_n1139), .A2(G171), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1065), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1058), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1120), .A2(new_n1121), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1050), .A2(new_n1047), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G288), .A2(G1976), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(new_n1045), .B2(new_n580), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1051), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1150), .A2(new_n1030), .B1(new_n1151), .B2(new_n1028), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n981), .A2(new_n963), .A3(G286), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT63), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1027), .B1(new_n1007), .B2(G8), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n1028), .A3(new_n1051), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1028), .A2(new_n1051), .A3(new_n1057), .A4(new_n1153), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1067), .A2(new_n1147), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n796), .B1(new_n582), .B2(new_n584), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n943), .B1(new_n1163), .B2(new_n944), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT108), .Z(new_n1165));
  AND4_X1   g740(.A1(new_n931), .A2(new_n928), .A3(new_n942), .A4(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1162), .A2(KEYINPUT126), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT126), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n960), .B1(new_n1167), .B2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g744(.A(G319), .B1(new_n641), .B2(new_n642), .ZN(new_n1171));
  NOR3_X1   g745(.A1(G229), .A2(G227), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n861), .B(new_n1172), .C1(new_n901), .C2(new_n902), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


