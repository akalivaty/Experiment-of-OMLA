

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XOR2_X1 U325 ( .A(G211GAT), .B(KEYINPUT88), .Z(n293) );
  XOR2_X1 U326 ( .A(KEYINPUT10), .B(G99GAT), .Z(n294) );
  XNOR2_X1 U327 ( .A(n523), .B(n522), .ZN(n553) );
  XNOR2_X1 U328 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n505) );
  XNOR2_X1 U329 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U330 ( .A(n449), .B(n318), .ZN(n319) );
  XNOR2_X1 U331 ( .A(n381), .B(G50GAT), .ZN(n382) );
  AND2_X1 U332 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U333 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U334 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U335 ( .A(n441), .B(KEYINPUT73), .ZN(n443) );
  NOR2_X1 U336 ( .A1(n414), .A2(n579), .ZN(n557) );
  XNOR2_X1 U337 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n522) );
  XNOR2_X1 U338 ( .A(n442), .B(n395), .ZN(n396) );
  XNOR2_X1 U339 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U340 ( .A(KEYINPUT26), .B(n415), .Z(n578) );
  XNOR2_X1 U341 ( .A(n397), .B(n396), .ZN(n414) );
  XNOR2_X1 U342 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U343 ( .A1(n559), .A2(n558), .ZN(n566) );
  XNOR2_X1 U344 ( .A(n454), .B(n453), .ZN(n584) );
  XOR2_X1 U345 ( .A(n338), .B(n337), .Z(n573) );
  INV_X1 U346 ( .A(G29GAT), .ZN(n457) );
  XNOR2_X1 U347 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U348 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  XOR2_X1 U349 ( .A(G57GAT), .B(G120GAT), .Z(n296) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(G1GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U352 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n298) );
  XNOR2_X1 U353 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U355 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U356 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n302) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT5), .B(n303), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U361 ( .A(G85GAT), .B(G162GAT), .Z(n307) );
  XNOR2_X1 U362 ( .A(G29GAT), .B(G148GAT), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U364 ( .A(n309), .B(n308), .Z(n316) );
  XOR2_X1 U365 ( .A(G127GAT), .B(KEYINPUT81), .Z(n311) );
  XNOR2_X1 U366 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n407) );
  XOR2_X1 U368 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n313) );
  XNOR2_X1 U369 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U371 ( .A(G141GAT), .B(n314), .Z(n378) );
  XNOR2_X1 U372 ( .A(n407), .B(n378), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n555) );
  XNOR2_X1 U374 ( .A(G190GAT), .B(G134GAT), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n294), .B(n317), .ZN(n320) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G92GAT), .Z(n449) );
  AND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XOR2_X1 U378 ( .A(KEYINPUT11), .B(n321), .Z(n324) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(G162GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n322), .B(KEYINPUT74), .ZN(n394) );
  XNOR2_X1 U381 ( .A(n394), .B(KEYINPUT66), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U383 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n326) );
  XNOR2_X1 U384 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  NAND2_X1 U386 ( .A1(n328), .A2(n327), .ZN(n332) );
  INV_X1 U387 ( .A(n327), .ZN(n330) );
  INV_X1 U388 ( .A(n328), .ZN(n329) );
  NAND2_X1 U389 ( .A1(n330), .A2(n329), .ZN(n331) );
  NAND2_X1 U390 ( .A1(n332), .A2(n331), .ZN(n338) );
  XNOR2_X1 U391 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n333), .B(G29GAT), .ZN(n334) );
  XOR2_X1 U393 ( .A(n334), .B(KEYINPUT7), .Z(n336) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G50GAT), .ZN(n335) );
  XOR2_X1 U395 ( .A(n336), .B(n335), .Z(n439) );
  INV_X1 U396 ( .A(n439), .ZN(n337) );
  INV_X1 U397 ( .A(n573), .ZN(n548) );
  XOR2_X1 U398 ( .A(KEYINPUT36), .B(n548), .Z(n591) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G211GAT), .Z(n340) );
  XNOR2_X1 U400 ( .A(G127GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT13), .Z(n444) );
  XOR2_X1 U403 ( .A(n341), .B(n444), .Z(n343) );
  XNOR2_X1 U404 ( .A(G183GAT), .B(G78GAT), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n349) );
  XOR2_X1 U406 ( .A(G1GAT), .B(G8GAT), .Z(n345) );
  XNOR2_X1 U407 ( .A(G22GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n435) );
  XOR2_X1 U409 ( .A(n435), .B(KEYINPUT77), .Z(n347) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n349), .B(n348), .Z(n357) );
  XOR2_X1 U413 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n351) );
  XNOR2_X1 U414 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U416 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n353) );
  XNOR2_X1 U417 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U420 ( .A(n357), .B(n356), .Z(n587) );
  INV_X1 U421 ( .A(n587), .ZN(n512) );
  XNOR2_X1 U422 ( .A(KEYINPUT17), .B(KEYINPUT83), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n358), .B(KEYINPUT18), .ZN(n359) );
  XOR2_X1 U424 ( .A(n359), .B(KEYINPUT19), .Z(n361) );
  XNOR2_X1 U425 ( .A(G183GAT), .B(G190GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n402) );
  XOR2_X1 U427 ( .A(G176GAT), .B(G64GAT), .Z(n440) );
  XNOR2_X1 U428 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n293), .B(n362), .ZN(n380) );
  XOR2_X1 U430 ( .A(n440), .B(n380), .Z(n364) );
  XNOR2_X1 U431 ( .A(G36GAT), .B(G218GAT), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U433 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n366) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U436 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U437 ( .A(KEYINPUT76), .B(G92GAT), .Z(n370) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U439 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(n371), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n402), .B(n374), .ZN(n552) );
  XOR2_X1 U443 ( .A(KEYINPUT27), .B(n552), .Z(n416) );
  INV_X1 U444 ( .A(n416), .ZN(n375) );
  NOR2_X1 U445 ( .A1(n555), .A2(n375), .ZN(n538) );
  INV_X1 U446 ( .A(KEYINPUT28), .ZN(n398) );
  XOR2_X1 U447 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n377) );
  XNOR2_X1 U448 ( .A(G22GAT), .B(KEYINPUT90), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n377), .B(n376), .ZN(n379) );
  XOR2_X1 U450 ( .A(n379), .B(n378), .Z(n385) );
  XOR2_X1 U451 ( .A(n380), .B(KEYINPUT87), .Z(n383) );
  NAND2_X1 U452 ( .A1(G228GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U454 ( .A(n386), .B(KEYINPUT24), .Z(n397) );
  INV_X1 U455 ( .A(G106GAT), .ZN(n387) );
  NAND2_X1 U456 ( .A1(n387), .A2(G148GAT), .ZN(n390) );
  INV_X1 U457 ( .A(G148GAT), .ZN(n388) );
  NAND2_X1 U458 ( .A1(n388), .A2(G106GAT), .ZN(n389) );
  NAND2_X1 U459 ( .A1(n390), .A2(n389), .ZN(n392) );
  XNOR2_X1 U460 ( .A(G204GAT), .B(G78GAT), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U462 ( .A(KEYINPUT71), .B(n393), .Z(n442) );
  XNOR2_X1 U463 ( .A(n394), .B(KEYINPUT86), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n398), .B(n414), .ZN(n501) );
  NAND2_X1 U465 ( .A1(n538), .A2(n501), .ZN(n525) );
  XOR2_X1 U466 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n400) );
  XNOR2_X1 U467 ( .A(G43GAT), .B(KEYINPUT84), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n411) );
  XOR2_X1 U470 ( .A(G169GAT), .B(G113GAT), .Z(n431) );
  XNOR2_X1 U471 ( .A(G99GAT), .B(G71GAT), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n403), .B(G120GAT), .ZN(n450) );
  XOR2_X1 U473 ( .A(n431), .B(n450), .Z(n405) );
  NAND2_X1 U474 ( .A1(G227GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U475 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U476 ( .A(n406), .B(G176GAT), .Z(n409) );
  XNOR2_X1 U477 ( .A(G15GAT), .B(n407), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n558) );
  XNOR2_X1 U480 ( .A(KEYINPUT85), .B(n558), .ZN(n412) );
  NOR2_X1 U481 ( .A1(n525), .A2(n412), .ZN(n413) );
  XOR2_X1 U482 ( .A(KEYINPUT96), .B(n413), .Z(n424) );
  NAND2_X1 U483 ( .A1(n414), .A2(n558), .ZN(n415) );
  NAND2_X1 U484 ( .A1(n416), .A2(n578), .ZN(n420) );
  NOR2_X1 U485 ( .A1(n558), .A2(n552), .ZN(n417) );
  NOR2_X1 U486 ( .A1(n414), .A2(n417), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n418), .B(KEYINPUT25), .ZN(n419) );
  NAND2_X1 U488 ( .A1(n420), .A2(n419), .ZN(n421) );
  NAND2_X1 U489 ( .A1(n421), .A2(n555), .ZN(n422) );
  XOR2_X1 U490 ( .A(KEYINPUT97), .B(n422), .Z(n423) );
  NAND2_X1 U491 ( .A1(n424), .A2(n423), .ZN(n465) );
  NAND2_X1 U492 ( .A1(n512), .A2(n465), .ZN(n425) );
  XOR2_X1 U493 ( .A(KEYINPUT101), .B(n425), .Z(n426) );
  NOR2_X1 U494 ( .A1(n591), .A2(n426), .ZN(n427) );
  XNOR2_X1 U495 ( .A(KEYINPUT37), .B(n427), .ZN(n494) );
  XOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n429) );
  XNOR2_X1 U497 ( .A(G197GAT), .B(G141GAT), .ZN(n428) );
  XNOR2_X1 U498 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U499 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U500 ( .A1(G229GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U501 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U502 ( .A(n434), .B(KEYINPUT29), .Z(n437) );
  XNOR2_X1 U503 ( .A(n435), .B(KEYINPUT30), .ZN(n436) );
  XNOR2_X1 U504 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U505 ( .A(n439), .B(n438), .Z(n581) );
  INV_X1 U506 ( .A(n581), .ZN(n481) );
  XOR2_X1 U507 ( .A(KEYINPUT70), .B(n481), .Z(n560) );
  XOR2_X1 U508 ( .A(n440), .B(KEYINPUT32), .Z(n441) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n454) );
  XOR2_X1 U510 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n447) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U512 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U513 ( .A(KEYINPUT31), .B(n448), .Z(n452) );
  XOR2_X1 U514 ( .A(n450), .B(n449), .Z(n451) );
  NAND2_X1 U515 ( .A1(n560), .A2(n584), .ZN(n467) );
  NOR2_X1 U516 ( .A1(n494), .A2(n467), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n455) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n479) );
  NOR2_X1 U519 ( .A1(n555), .A2(n479), .ZN(n460) );
  XNOR2_X1 U520 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n458) );
  INV_X1 U521 ( .A(G43GAT), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n558), .A2(n479), .ZN(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT40), .B(n461), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  NAND2_X1 U525 ( .A1(n573), .A2(n587), .ZN(n464) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n464), .Z(n466) );
  NAND2_X1 U527 ( .A1(n466), .A2(n465), .ZN(n482) );
  OR2_X1 U528 ( .A1(n467), .A2(n482), .ZN(n476) );
  NOR2_X1 U529 ( .A1(n555), .A2(n476), .ZN(n468) );
  XOR2_X1 U530 ( .A(n468), .B(KEYINPUT34), .Z(n469) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n469), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n552), .A2(n476), .ZN(n470) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(n470), .Z(n471) );
  XNOR2_X1 U534 ( .A(G8GAT), .B(n471), .ZN(G1325GAT) );
  NOR2_X1 U535 ( .A1(n476), .A2(n558), .ZN(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n473) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT100), .ZN(n472) );
  XNOR2_X1 U538 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U539 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n501), .A2(n476), .ZN(n477) );
  XOR2_X1 U541 ( .A(G22GAT), .B(n477), .Z(G1327GAT) );
  NOR2_X1 U542 ( .A1(n552), .A2(n479), .ZN(n478) );
  XOR2_X1 U543 ( .A(G36GAT), .B(n478), .Z(G1329GAT) );
  NOR2_X1 U544 ( .A1(n501), .A2(n479), .ZN(n480) );
  XOR2_X1 U545 ( .A(G50GAT), .B(n480), .Z(G1331GAT) );
  XNOR2_X1 U546 ( .A(KEYINPUT41), .B(n584), .ZN(n504) );
  NAND2_X1 U547 ( .A1(n481), .A2(n504), .ZN(n493) );
  NOR2_X1 U548 ( .A1(n482), .A2(n493), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n483), .B(KEYINPUT105), .ZN(n490) );
  NOR2_X1 U550 ( .A1(n555), .A2(n490), .ZN(n485) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n484) );
  XNOR2_X1 U552 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U553 ( .A(G57GAT), .B(n486), .Z(G1332GAT) );
  NOR2_X1 U554 ( .A1(n552), .A2(n490), .ZN(n487) );
  XOR2_X1 U555 ( .A(G64GAT), .B(n487), .Z(G1333GAT) );
  NOR2_X1 U556 ( .A1(n558), .A2(n490), .ZN(n488) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(n488), .Z(n489) );
  XNOR2_X1 U558 ( .A(G71GAT), .B(n489), .ZN(G1334GAT) );
  NOR2_X1 U559 ( .A1(n501), .A2(n490), .ZN(n492) );
  XNOR2_X1 U560 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n492), .B(n491), .ZN(G1335GAT) );
  OR2_X1 U562 ( .A1(n494), .A2(n493), .ZN(n500) );
  NOR2_X1 U563 ( .A1(n555), .A2(n500), .ZN(n496) );
  XNOR2_X1 U564 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n496), .B(n495), .ZN(G1336GAT) );
  NOR2_X1 U566 ( .A1(n552), .A2(n500), .ZN(n497) );
  XOR2_X1 U567 ( .A(G92GAT), .B(n497), .Z(G1337GAT) );
  NOR2_X1 U568 ( .A1(n558), .A2(n500), .ZN(n498) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(n498), .Z(n499) );
  XNOR2_X1 U570 ( .A(G99GAT), .B(n499), .ZN(G1338GAT) );
  NOR2_X1 U571 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U572 ( .A(KEYINPUT44), .B(n502), .Z(n503) );
  XNOR2_X1 U573 ( .A(G106GAT), .B(n503), .ZN(G1339GAT) );
  NAND2_X1 U574 ( .A1(n504), .A2(n581), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n587), .B(KEYINPUT109), .ZN(n567) );
  NAND2_X1 U576 ( .A1(n507), .A2(n567), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(KEYINPUT111), .ZN(n509) );
  NAND2_X1 U578 ( .A1(n509), .A2(n573), .ZN(n511) );
  XNOR2_X1 U579 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n510) );
  XNOR2_X1 U580 ( .A(n511), .B(n510), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n591), .A2(n512), .ZN(n515) );
  XNOR2_X1 U582 ( .A(KEYINPUT113), .B(KEYINPUT45), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n513), .B(KEYINPUT65), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n518) );
  INV_X1 U585 ( .A(n560), .ZN(n516) );
  AND2_X1 U586 ( .A1(n584), .A2(n516), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n519), .B(KEYINPUT114), .ZN(n520) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n523) );
  OR2_X1 U589 ( .A1(n558), .A2(n553), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n560), .A2(n531), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U594 ( .A1(n531), .A2(n504), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n530) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT115), .Z(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  INV_X1 U598 ( .A(n531), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n567), .A2(n535), .ZN(n533) );
  XNOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U603 ( .A1(n573), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n538), .A2(n578), .ZN(n539) );
  NOR2_X1 U607 ( .A1(n553), .A2(n539), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n581), .A2(n549), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n540), .B(KEYINPUT118), .ZN(n541) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n543) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(n544), .Z(n546) );
  NAND2_X1 U615 ( .A1(n549), .A2(n504), .ZN(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n587), .A2(n549), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT121), .Z(n551) );
  NAND2_X1 U620 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U621 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n554), .B(KEYINPUT54), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n579) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT55), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n566), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT122), .B(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  NAND2_X1 U630 ( .A1(n566), .A2(n504), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  INV_X1 U633 ( .A(n566), .ZN(n572) );
  NOR2_X1 U634 ( .A1(n567), .A2(n572), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n571) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(G1351GAT) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(KEYINPUT126), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(n577), .Z(n583) );
  INV_X1 U645 ( .A(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U650 ( .A(n588), .ZN(n590) );
  OR2_X1 U651 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

