

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n734) );
  NOR2_X1 U561 ( .A1(G651), .A2(n618), .ZN(n641) );
  XNOR2_X1 U562 ( .A(n761), .B(KEYINPUT30), .ZN(n762) );
  INV_X1 U563 ( .A(KEYINPUT101), .ZN(n763) );
  NAND2_X1 U564 ( .A1(n724), .A2(n723), .ZN(n777) );
  NAND2_X1 U565 ( .A1(n777), .A2(G8), .ZN(n799) );
  XNOR2_X1 U566 ( .A(n690), .B(n689), .ZN(n723) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n649) );
  AND2_X1 U568 ( .A1(n885), .A2(G137), .ZN(n530) );
  AND2_X1 U569 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U570 ( .A(G2104), .ZN(n526) );
  NOR2_X1 U571 ( .A1(n526), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U572 ( .A(n523), .B(KEYINPUT64), .ZN(n886) );
  NAND2_X1 U573 ( .A1(n886), .A2(G101), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n524), .Z(n532) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n525), .Z(n885) );
  AND2_X1 U577 ( .A1(n526), .A2(G2105), .ZN(n881) );
  NAND2_X1 U578 ( .A1(G125), .A2(n881), .ZN(n528) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U580 ( .A1(G113), .A2(n882), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n531) );
  INV_X1 U583 ( .A(G651), .ZN(n536) );
  NOR2_X1 U584 ( .A1(G543), .A2(n536), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n533), .Z(n639) );
  NAND2_X1 U586 ( .A1(G64), .A2(n639), .ZN(n535) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n618) );
  NAND2_X1 U588 ( .A1(G52), .A2(n641), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X1 U590 ( .A1(n618), .A2(n536), .ZN(n645) );
  NAND2_X1 U591 ( .A1(G77), .A2(n645), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G90), .A2(n649), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(G171) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G69), .ZN(G235) );
  INV_X1 U598 ( .A(G132), .ZN(G219) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  NAND2_X1 U600 ( .A1(G7), .A2(G661), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n542), .B(KEYINPUT10), .ZN(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT70), .B(n543), .ZN(G223) );
  INV_X1 U603 ( .A(G223), .ZN(n830) );
  NAND2_X1 U604 ( .A1(n830), .A2(G567), .ZN(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT71), .ZN(n545) );
  XNOR2_X1 U606 ( .A(KEYINPUT11), .B(n545), .ZN(G234) );
  NAND2_X1 U607 ( .A1(G56), .A2(n639), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT14), .B(n546), .Z(n552) );
  NAND2_X1 U609 ( .A1(n649), .A2(G81), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT12), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G68), .A2(n645), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT13), .B(n550), .Z(n551) );
  NOR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n641), .A2(G43), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n972) );
  INV_X1 U617 ( .A(n972), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n555), .A2(G860), .ZN(G153) );
  XOR2_X1 U619 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U620 ( .A1(G92), .A2(n649), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G66), .A2(n639), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G54), .A2(n641), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G79), .A2(n645), .ZN(n558) );
  XNOR2_X1 U625 ( .A(KEYINPUT73), .B(n558), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT15), .ZN(n900) );
  INV_X1 U629 ( .A(n900), .ZN(n975) );
  INV_X1 U630 ( .A(G868), .ZN(n665) );
  NAND2_X1 U631 ( .A1(n975), .A2(n665), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT74), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G301), .A2(G868), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT75), .B(n567), .Z(G284) );
  NAND2_X1 U636 ( .A1(G63), .A2(n639), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G51), .A2(n641), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U639 ( .A(KEYINPUT6), .B(n570), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G89), .A2(n649), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT4), .ZN(n572) );
  XNOR2_X1 U642 ( .A(n572), .B(KEYINPUT76), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G76), .A2(n645), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U645 ( .A(n575), .B(KEYINPUT5), .Z(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U647 ( .A(KEYINPUT7), .B(n578), .Z(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT77), .B(n579), .Z(G168) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(n639), .A2(G65), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G78), .A2(n645), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G91), .A2(n649), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n641), .A2(G53), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n582), .Z(n583) );
  NOR2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT69), .B(n587), .Z(G299) );
  NAND2_X1 U659 ( .A1(G286), .A2(G868), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G299), .A2(n665), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(G297) );
  INV_X1 U662 ( .A(G559), .ZN(n590) );
  NOR2_X1 U663 ( .A1(G860), .A2(n590), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT78), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n975), .A2(n592), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT79), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U668 ( .A1(G868), .A2(n972), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n900), .A2(G868), .ZN(n595) );
  NOR2_X1 U670 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G123), .A2(n881), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT18), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT80), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G111), .A2(n882), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G135), .A2(n885), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G99), .A2(n886), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n931) );
  XNOR2_X1 U681 ( .A(n931), .B(G2096), .ZN(n607) );
  INV_X1 U682 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G67), .A2(n639), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G55), .A2(n641), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U687 ( .A(KEYINPUT82), .B(n610), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G80), .A2(n645), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G93), .A2(n649), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  OR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n664) );
  NAND2_X1 U692 ( .A1(n900), .A2(G559), .ZN(n661) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(n972), .Z(n615) );
  XNOR2_X1 U694 ( .A(n661), .B(n615), .ZN(n616) );
  NOR2_X1 U695 ( .A1(G860), .A2(n616), .ZN(n617) );
  XOR2_X1 U696 ( .A(n664), .B(n617), .Z(G145) );
  NAND2_X1 U697 ( .A1(G49), .A2(n641), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G87), .A2(n618), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n639), .A2(n621), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G74), .A2(G651), .ZN(n622) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(n622), .Z(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U704 ( .A1(G61), .A2(n639), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G86), .A2(n649), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT84), .B(n627), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n645), .A2(G73), .ZN(n628) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n628), .Z(n629) );
  NOR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n641), .A2(G48), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G75), .A2(n645), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G88), .A2(n649), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G62), .A2(n639), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G50), .A2(n641), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(G166) );
  NAND2_X1 U720 ( .A1(G60), .A2(n639), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n640), .B(KEYINPUT66), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G47), .A2(n641), .ZN(n642) );
  XOR2_X1 U723 ( .A(KEYINPUT67), .B(n642), .Z(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G72), .A2(n645), .ZN(n646) );
  XNOR2_X1 U726 ( .A(KEYINPUT65), .B(n646), .ZN(n647) );
  NOR2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n649), .A2(G85), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(G290) );
  XOR2_X1 U730 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n652) );
  XNOR2_X1 U731 ( .A(G305), .B(n652), .ZN(n653) );
  XOR2_X1 U732 ( .A(n653), .B(KEYINPUT85), .Z(n655) );
  XNOR2_X1 U733 ( .A(G166), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U735 ( .A(n664), .B(n656), .Z(n658) );
  INV_X1 U736 ( .A(G299), .ZN(n737) );
  XNOR2_X1 U737 ( .A(n972), .B(n737), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U739 ( .A(n659), .B(G290), .Z(n660) );
  XNOR2_X1 U740 ( .A(G288), .B(n660), .ZN(n902) );
  XOR2_X1 U741 ( .A(n902), .B(n661), .Z(n662) );
  XNOR2_X1 U742 ( .A(KEYINPUT88), .B(n662), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U745 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n672) );
  XNOR2_X1 U753 ( .A(KEYINPUT22), .B(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n673), .A2(G96), .ZN(n674) );
  NOR2_X1 U755 ( .A1(n674), .A2(G218), .ZN(n675) );
  XNOR2_X1 U756 ( .A(n675), .B(KEYINPUT89), .ZN(n837) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n837), .ZN(n679) );
  NAND2_X1 U758 ( .A1(G120), .A2(G108), .ZN(n676) );
  NOR2_X1 U759 ( .A1(G235), .A2(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G57), .A2(n677), .ZN(n836) );
  NAND2_X1 U761 ( .A1(G567), .A2(n836), .ZN(n678) );
  NAND2_X1 U762 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U763 ( .A(KEYINPUT90), .B(n680), .Z(G319) );
  INV_X1 U764 ( .A(G319), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n834) );
  NAND2_X1 U767 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U768 ( .A1(G138), .A2(n885), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G102), .A2(n886), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G126), .A2(n881), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G114), .A2(n882), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U774 ( .A1(n688), .A2(n687), .ZN(G164) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n724) );
  INV_X1 U777 ( .A(KEYINPUT91), .ZN(n690) );
  AND2_X1 U778 ( .A1(G40), .A2(G160), .ZN(n689) );
  INV_X1 U779 ( .A(n723), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n724), .A2(n691), .ZN(n825) );
  XNOR2_X1 U781 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n702) );
  NAND2_X1 U782 ( .A1(G128), .A2(n881), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G116), .A2(n882), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U785 ( .A(KEYINPUT35), .B(n694), .ZN(n700) );
  NAND2_X1 U786 ( .A1(G140), .A2(n885), .ZN(n696) );
  NAND2_X1 U787 ( .A1(G104), .A2(n886), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n698) );
  XOR2_X1 U789 ( .A(KEYINPUT34), .B(KEYINPUT92), .Z(n697) );
  XNOR2_X1 U790 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n702), .B(n701), .ZN(n864) );
  XNOR2_X1 U793 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NOR2_X1 U794 ( .A1(n864), .A2(n822), .ZN(n927) );
  NAND2_X1 U795 ( .A1(n825), .A2(n927), .ZN(n820) );
  NAND2_X1 U796 ( .A1(G119), .A2(n881), .ZN(n704) );
  NAND2_X1 U797 ( .A1(G107), .A2(n882), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n886), .A2(G95), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n705), .B(KEYINPUT94), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n885), .A2(G131), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n868) );
  INV_X1 U804 ( .A(G1991), .ZN(n814) );
  NOR2_X1 U805 ( .A1(n868), .A2(n814), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n886), .A2(G105), .ZN(n710) );
  XNOR2_X1 U807 ( .A(n710), .B(KEYINPUT38), .ZN(n717) );
  NAND2_X1 U808 ( .A1(G141), .A2(n885), .ZN(n712) );
  NAND2_X1 U809 ( .A1(G117), .A2(n882), .ZN(n711) );
  NAND2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G129), .A2(n881), .ZN(n713) );
  XNOR2_X1 U812 ( .A(KEYINPUT95), .B(n713), .ZN(n714) );
  NOR2_X1 U813 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n865) );
  AND2_X1 U815 ( .A1(n865), .A2(G1996), .ZN(n718) );
  NOR2_X1 U816 ( .A1(n719), .A2(n718), .ZN(n933) );
  INV_X1 U817 ( .A(n825), .ZN(n720) );
  NOR2_X1 U818 ( .A1(n933), .A2(n720), .ZN(n817) );
  INV_X1 U819 ( .A(n817), .ZN(n721) );
  NAND2_X1 U820 ( .A1(n820), .A2(n721), .ZN(n722) );
  XNOR2_X1 U821 ( .A(KEYINPUT96), .B(n722), .ZN(n811) );
  OR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n793) );
  XNOR2_X1 U823 ( .A(n793), .B(KEYINPUT24), .ZN(n725) );
  NOR2_X1 U824 ( .A1(n799), .A2(n725), .ZN(n726) );
  XNOR2_X1 U825 ( .A(n726), .B(KEYINPUT97), .ZN(n791) );
  NOR2_X1 U826 ( .A1(G1966), .A2(n799), .ZN(n771) );
  XOR2_X1 U827 ( .A(G2078), .B(KEYINPUT25), .Z(n959) );
  XOR2_X1 U828 ( .A(KEYINPUT98), .B(n777), .Z(n745) );
  INV_X1 U829 ( .A(n745), .ZN(n731) );
  NOR2_X1 U830 ( .A1(n959), .A2(n731), .ZN(n728) );
  INV_X1 U831 ( .A(n777), .ZN(n738) );
  NOR2_X1 U832 ( .A1(n738), .A2(G1961), .ZN(n727) );
  NOR2_X1 U833 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U834 ( .A(KEYINPUT99), .B(n729), .ZN(n759) );
  NAND2_X1 U835 ( .A1(n759), .A2(G171), .ZN(n758) );
  NAND2_X1 U836 ( .A1(G2072), .A2(n745), .ZN(n730) );
  XNOR2_X1 U837 ( .A(n730), .B(KEYINPUT27), .ZN(n733) );
  AND2_X1 U838 ( .A1(n731), .A2(G1956), .ZN(n732) );
  NOR2_X1 U839 ( .A1(n733), .A2(n732), .ZN(n736) );
  NOR2_X1 U840 ( .A1(n737), .A2(n736), .ZN(n735) );
  XNOR2_X1 U841 ( .A(n735), .B(n734), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n737), .A2(n736), .ZN(n753) );
  AND2_X1 U843 ( .A1(n738), .A2(G1996), .ZN(n740) );
  XOR2_X1 U844 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n739) );
  XNOR2_X1 U845 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U846 ( .A1(n777), .A2(G1341), .ZN(n741) );
  NAND2_X1 U847 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U848 ( .A1(n972), .A2(n743), .ZN(n744) );
  OR2_X1 U849 ( .A1(n900), .A2(n744), .ZN(n751) );
  NAND2_X1 U850 ( .A1(n900), .A2(n744), .ZN(n749) );
  NAND2_X1 U851 ( .A1(G2067), .A2(n745), .ZN(n747) );
  NAND2_X1 U852 ( .A1(G1348), .A2(n777), .ZN(n746) );
  NAND2_X1 U853 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U854 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U855 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U856 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U857 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U858 ( .A(KEYINPUT29), .B(n756), .Z(n757) );
  NAND2_X1 U859 ( .A1(n758), .A2(n757), .ZN(n769) );
  NOR2_X1 U860 ( .A1(G171), .A2(n759), .ZN(n766) );
  NOR2_X1 U861 ( .A1(G2084), .A2(n777), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n771), .A2(n773), .ZN(n760) );
  NAND2_X1 U863 ( .A1(G8), .A2(n760), .ZN(n761) );
  NOR2_X1 U864 ( .A1(G168), .A2(n762), .ZN(n764) );
  XNOR2_X1 U865 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U866 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U867 ( .A(KEYINPUT31), .B(n767), .Z(n768) );
  NAND2_X1 U868 ( .A1(n769), .A2(n768), .ZN(n776) );
  INV_X1 U869 ( .A(n776), .ZN(n770) );
  NOR2_X1 U870 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U871 ( .A(n772), .B(KEYINPUT102), .ZN(n775) );
  NAND2_X1 U872 ( .A1(n773), .A2(G8), .ZN(n774) );
  NAND2_X1 U873 ( .A1(n775), .A2(n774), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n776), .A2(G286), .ZN(n782) );
  NOR2_X1 U875 ( .A1(G1971), .A2(n799), .ZN(n779) );
  NOR2_X1 U876 ( .A1(G2090), .A2(n777), .ZN(n778) );
  NOR2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U878 ( .A1(n780), .A2(G303), .ZN(n781) );
  NAND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U880 ( .A1(G8), .A2(n783), .ZN(n784) );
  XNOR2_X1 U881 ( .A(n784), .B(KEYINPUT32), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n795) );
  NOR2_X1 U883 ( .A1(G2090), .A2(G303), .ZN(n787) );
  NAND2_X1 U884 ( .A1(G8), .A2(n787), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n795), .A2(n788), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n789), .A2(n799), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n809) );
  NAND2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n988) );
  NOR2_X1 U890 ( .A1(G1976), .A2(G288), .ZN(n801) );
  NOR2_X1 U891 ( .A1(G1971), .A2(G303), .ZN(n794) );
  NOR2_X1 U892 ( .A1(n801), .A2(n794), .ZN(n982) );
  NAND2_X1 U893 ( .A1(n795), .A2(n982), .ZN(n797) );
  AND2_X1 U894 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NOR2_X1 U895 ( .A1(n984), .A2(n799), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  INV_X1 U897 ( .A(KEYINPUT33), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n798), .A2(n803), .ZN(n806) );
  INV_X1 U899 ( .A(n799), .ZN(n800) );
  NAND2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U902 ( .A(n804), .B(KEYINPUT103), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n988), .A2(n807), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n813) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U908 ( .A1(n980), .A2(n825), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n828) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n865), .ZN(n944) );
  AND2_X1 U911 ( .A1(n814), .A2(n868), .ZN(n935) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n935), .A2(n815), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U915 ( .A1(n944), .A2(n818), .ZN(n819) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n864), .A2(n822), .ZN(n926) );
  NAND2_X1 U919 ( .A1(n823), .A2(n926), .ZN(n824) );
  XNOR2_X1 U920 ( .A(KEYINPUT104), .B(n824), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n829), .ZN(G329) );
  NAND2_X1 U924 ( .A1(n830), .A2(G2106), .ZN(n831) );
  XOR2_X1 U925 ( .A(KEYINPUT111), .B(n831), .Z(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U927 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n833) );
  XNOR2_X1 U929 ( .A(KEYINPUT112), .B(n833), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G188) );
  XNOR2_X1 U931 ( .A(G120), .B(KEYINPUT113), .ZN(G236) );
  XOR2_X1 U932 ( .A(G108), .B(KEYINPUT120), .Z(G238) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U937 ( .A(G1961), .B(KEYINPUT114), .ZN(n847) );
  XOR2_X1 U938 ( .A(G1956), .B(G1971), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1976), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U941 ( .A(G1981), .B(G1966), .Z(n841) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U944 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2474), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U948 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2084), .B(G2078), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U957 ( .A1(n882), .A2(G112), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G100), .A2(n886), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n881), .A2(G124), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G136), .A2(n885), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(n861), .Z(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U966 ( .A(G160), .B(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n867), .B(n931), .Z(n870) );
  XNOR2_X1 U969 ( .A(n868), .B(G162), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n898) );
  NAND2_X1 U971 ( .A1(G139), .A2(n885), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G103), .A2(n886), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U974 ( .A1(n882), .A2(G115), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT116), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G127), .A2(n881), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(KEYINPUT117), .B(n876), .ZN(n877) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n877), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT118), .B(n880), .Z(n938) );
  NAND2_X1 U982 ( .A1(G130), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G118), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G142), .A2(n885), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G106), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(n889), .B(KEYINPUT45), .Z(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(KEYINPUT48), .B(n892), .Z(n893) );
  XOR2_X1 U991 ( .A(n893), .B(KEYINPUT46), .Z(n895) );
  XNOR2_X1 U992 ( .A(G164), .B(KEYINPUT119), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n938), .B(n896), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G171), .B(n900), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(G286), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U1001 ( .A(G2430), .B(G2454), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n918) );
  XOR2_X1 U1004 ( .A(G2446), .B(KEYINPUT105), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G2435), .B(G2451), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n916) );
  XOR2_X1 U1007 ( .A(KEYINPUT106), .B(G2443), .Z(n910) );
  XNOR2_X1 U1008 ( .A(G2438), .B(KEYINPUT109), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1010 ( .A(KEYINPUT108), .B(G2427), .Z(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT107), .B(KEYINPUT110), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1013 ( .A(n914), .B(n913), .Z(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n919), .A2(G14), .ZN(n925) );
  NAND2_X1 U1017 ( .A1(n925), .A2(G319), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G57), .ZN(G237) );
  INV_X1 U1025 ( .A(n925), .ZN(G401) );
  INV_X1 U1026 ( .A(n926), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n937) );
  XNOR2_X1 U1028 ( .A(G2084), .B(G160), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT121), .B(n929), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n949) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n940) );
  XNOR2_X1 U1035 ( .A(G2072), .B(n938), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(KEYINPUT122), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n942), .B(KEYINPUT50), .ZN(n947) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n945), .Z(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n950), .ZN(n951) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n1023), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n952), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1048 ( .A(G2084), .B(G34), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(KEYINPUT54), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n969) );
  XOR2_X1 U1052 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n967) );
  XOR2_X1 U1053 ( .A(G2067), .B(G26), .Z(n956) );
  NAND2_X1 U1054 ( .A1(n956), .A2(G28), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(G1996), .B(G32), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G1991), .B(G25), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(G27), .B(n959), .ZN(n960) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1063 ( .A(n967), .B(n966), .Z(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n1024) );
  NOR2_X1 U1065 ( .A1(G29), .A2(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n1024), .A2(n970), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(G11), .A2(n971), .ZN(n1028) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XOR2_X1 U1069 ( .A(G171), .B(G1961), .Z(n974) );
  XNOR2_X1 U1070 ( .A(n972), .B(G1341), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n993) );
  XNOR2_X1 U1072 ( .A(G1348), .B(KEYINPUT124), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(n976), .B(n975), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(G1956), .B(G299), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n986) );
  AND2_X1 U1076 ( .A1(G303), .A2(G1971), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n991) );
  XOR2_X1 U1081 ( .A(G1966), .B(G168), .Z(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n989), .B(KEYINPUT57), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1021) );
  INV_X1 U1087 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(G4), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT125), .B(G1341), .Z(n1001) );
  XNOR2_X1 U1095 ( .A(G19), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(n1005), .B(KEYINPUT60), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G21), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1006) );
  NOR2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G1976), .B(G23), .ZN(n1011) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1010) );
  NOR2_X1 U1105 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1012) );
  NAND2_X1 U1107 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1109 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT127), .ZN(n1026) );
  OR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

