//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n202), .A2(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(G8gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n202), .A2(G1gat), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(new_n205), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT83), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n211), .A3(KEYINPUT83), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G64gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G57gat), .ZN(new_n218));
  INV_X1    g017(.A(G57gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G64gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT9), .ZN(new_n222));
  NAND2_X1  g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  OR2_X1    g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT85), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT85), .B1(new_n218), .B2(new_n220), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT86), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT86), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n226), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT21), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(G183gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n239), .A2(G231gat), .A3(G233gat), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G231gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n240), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n238), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G155gat), .ZN(new_n245));
  INV_X1    g044(.A(G211gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n241), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n241), .B2(new_n244), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT21), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OR3_X1    g053(.A1(new_n249), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n249), .B2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(KEYINPUT87), .A2(G85gat), .A3(G92gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G99gat), .A2(G106gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT8), .ZN(new_n263));
  INV_X1    g062(.A(G85gat), .ZN(new_n264));
  INV_X1    g063(.A(G92gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(KEYINPUT87), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n261), .A2(new_n263), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G99gat), .B(G106gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n272));
  AOI22_X1  g071(.A1(KEYINPUT8), .A2(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(new_n269), .A3(new_n261), .A4(new_n267), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(new_n272), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(G29gat), .A2(G36gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT14), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G29gat), .A2(G36gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G43gat), .B(G50gat), .Z(new_n287));
  INV_X1    g086(.A(KEYINPUT15), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n281), .B(KEYINPUT82), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n289), .A2(new_n280), .A3(new_n284), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT17), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(new_n286), .B2(new_n291), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n277), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G190gat), .B(G218gat), .Z(new_n297));
  AND3_X1   g096(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n275), .A2(new_n276), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n292), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n296), .B2(new_n300), .ZN(new_n302));
  XNOR2_X1  g101(.A(G134gat), .B(G162gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n297), .B(new_n305), .C1(new_n296), .C2(new_n300), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n301), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n296), .A2(new_n297), .A3(new_n300), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n258), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT11), .B(G169gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(G197gat), .ZN(new_n315));
  XOR2_X1   g114(.A(G113gat), .B(G141gat), .Z(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(KEYINPUT12), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n212), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n293), .B2(new_n295), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n214), .A2(new_n215), .A3(new_n292), .ZN(new_n322));
  NAND2_X1  g121(.A1(G229gat), .A2(G233gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT18), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT18), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n321), .A2(new_n326), .A3(new_n322), .A4(new_n323), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n329));
  INV_X1    g128(.A(new_n292), .ZN(new_n330));
  INV_X1    g129(.A(new_n215), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT83), .B1(new_n208), .B2(new_n211), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n322), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n323), .B(KEYINPUT13), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n329), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI211_X1 g136(.A(KEYINPUT84), .B(new_n335), .C1(new_n333), .C2(new_n322), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n319), .B1(new_n328), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n327), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(new_n318), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT85), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n221), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G57gat), .B(G64gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT86), .B1(new_n349), .B2(new_n228), .ZN(new_n350));
  INV_X1    g149(.A(new_n234), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n225), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n277), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT90), .B1(new_n235), .B2(new_n299), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n235), .A2(new_n274), .A3(new_n271), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n235), .A2(KEYINPUT10), .A3(new_n299), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G230gat), .A2(G233gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n363));
  INV_X1    g162(.A(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G120gat), .B(G148gat), .ZN(new_n367));
  INV_X1    g166(.A(G176gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G204gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n362), .A2(new_n365), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n344), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT71), .B(G71gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G15gat), .B(G43gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT33), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G169gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n368), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(KEYINPUT65), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT23), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G183gat), .ZN(new_n391));
  INV_X1    g190(.A(G190gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT24), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n394), .A2(KEYINPUT24), .ZN(new_n396));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT64), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n399), .A2(new_n400), .B1(new_n386), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n390), .A2(new_n395), .A3(new_n396), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT23), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n395), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n403), .A2(KEYINPUT25), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n399), .A2(new_n400), .B1(new_n386), .B2(KEYINPUT26), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n387), .A2(new_n389), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(KEYINPUT26), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT27), .B(G183gat), .Z(new_n415));
  INV_X1    g214(.A(KEYINPUT66), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n391), .A2(KEYINPUT27), .ZN(new_n418));
  AOI21_X1  g217(.A(G190gat), .B1(new_n418), .B2(KEYINPUT66), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT28), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n415), .A2(new_n421), .A3(G190gat), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n394), .B(new_n413), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n410), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(G113gat), .A2(G120gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT1), .ZN(new_n426));
  NAND2_X1  g225(.A1(G113gat), .A2(G120gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT68), .ZN(new_n429));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT70), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n424), .A2(KEYINPUT70), .A3(new_n431), .ZN(new_n435));
  INV_X1    g234(.A(new_n430), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n429), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n410), .A2(new_n423), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT69), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n410), .A2(new_n423), .A3(new_n440), .A4(new_n437), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n434), .A2(new_n435), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT32), .B(new_n384), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(new_n435), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT70), .B1(new_n424), .B2(new_n431), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n443), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT32), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(KEYINPUT33), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n444), .B1(new_n451), .B2(new_n380), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT34), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT34), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n442), .A2(new_n454), .A3(new_n443), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  OAI22_X1  g257(.A1(new_n442), .A2(new_n443), .B1(KEYINPUT32), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n381), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n460), .A2(new_n444), .A3(new_n453), .A4(new_n455), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(G22gat), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G155gat), .B(G162gat), .Z(new_n465));
  XOR2_X1   g264(.A(KEYINPUT76), .B(KEYINPUT2), .Z(new_n466));
  XNOR2_X1  g265(.A(G141gat), .B(G148gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G141gat), .B(G148gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G155gat), .B(G162gat), .ZN(new_n470));
  INV_X1    g269(.A(G162gat), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT2), .B1(new_n471), .B2(KEYINPUT77), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(KEYINPUT73), .A2(G218gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(KEYINPUT73), .A2(G218gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(G211gat), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT22), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G197gat), .B(G204gat), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G211gat), .B(G218gat), .Z(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n478), .B2(new_n477), .ZN(new_n485));
  INV_X1    g284(.A(new_n483), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT74), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n483), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n474), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n490), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(G228gat), .B(G233gat), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G50gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G228gat), .A2(G233gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n497), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT80), .B1(new_n482), .B2(new_n483), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT29), .B1(new_n504), .B2(new_n487), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n486), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT3), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n502), .B(new_n503), .C1(new_n507), .C2(new_n474), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n499), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n501), .B1(new_n499), .B2(new_n508), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n464), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n499), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n500), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n499), .A2(new_n501), .A3(new_n508), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n463), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n457), .A2(new_n461), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n495), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT29), .B1(new_n410), .B2(new_n423), .ZN(new_n519));
  AND2_X1   g318(.A1(G226gat), .A2(G233gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n424), .A2(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n424), .A2(new_n520), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n524), .B(new_n495), .C1(new_n520), .C2(new_n519), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT75), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G8gat), .B(G36gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(new_n217), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n265), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n530), .ZN(new_n533));
  INV_X1    g332(.A(new_n523), .ZN(new_n534));
  INV_X1    g333(.A(new_n525), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n537), .B(new_n530), .C1(new_n523), .C2(new_n525), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n437), .A2(new_n474), .ZN(new_n544));
  AND2_X1   g343(.A1(G225gat), .A2(G233gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n468), .A2(new_n473), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT3), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n496), .A2(new_n431), .A3(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n437), .B2(new_n474), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n546), .B(new_n549), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT5), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n431), .A2(new_n547), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n544), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n556), .B2(new_n545), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT0), .B(G57gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G85gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(G1gat), .B(G29gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  NOR2_X1   g361(.A1(new_n545), .A2(KEYINPUT5), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n549), .B(new_n563), .C1(new_n550), .C2(new_n552), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n558), .A2(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n558), .A2(KEYINPUT78), .A3(new_n562), .A4(new_n564), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n567), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n517), .A2(new_n542), .A3(new_n543), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n580), .A2(new_n563), .B1(new_n553), .B2(new_n557), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n578), .B1(new_n581), .B2(new_n562), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n568), .A2(KEYINPUT79), .A3(new_n569), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n574), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n538), .A3(new_n532), .A4(new_n540), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n457), .A2(new_n461), .A3(new_n516), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT35), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n577), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT75), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT37), .B1(new_n591), .B2(new_n526), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n523), .A2(new_n525), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n592), .B(KEYINPUT38), .C1(KEYINPUT37), .C2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n523), .A2(new_n525), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n533), .B1(KEYINPUT37), .B2(new_n595), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(new_n575), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n579), .A2(new_n545), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n569), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n545), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n603), .B(KEYINPUT39), .C1(new_n545), .C2(new_n556), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(KEYINPUT40), .A3(new_n604), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n541), .A2(new_n609), .A3(new_n570), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n599), .A2(new_n610), .A3(new_n516), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n452), .A2(new_n456), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n460), .A2(new_n444), .B1(new_n453), .B2(new_n455), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n457), .A2(new_n461), .A3(KEYINPUT36), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n516), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n611), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT81), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n590), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n590), .B2(new_n620), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n313), .B(new_n376), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT91), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n590), .A2(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT81), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n590), .A2(new_n620), .A3(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT91), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n629), .A2(new_n630), .A3(new_n313), .A4(new_n376), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n586), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(G8gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT92), .B1(new_n632), .B2(new_n541), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n639));
  AOI211_X1 g438(.A(new_n639), .B(new_n542), .C1(new_n625), .C2(new_n631), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT16), .B(G8gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(KEYINPUT42), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n637), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n632), .ZN(new_n647));
  NOR4_X1   g446(.A1(new_n647), .A2(new_n636), .A3(new_n542), .A4(new_n642), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT93), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT93), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n638), .A2(new_n640), .A3(new_n644), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n637), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(G1325gat));
  NOR2_X1   g453(.A1(new_n613), .A2(new_n614), .ZN(new_n655));
  AOI21_X1  g454(.A(G15gat), .B1(new_n632), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n632), .A2(G15gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n617), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(G1326gat));
  NAND2_X1  g458(.A1(new_n632), .A2(new_n618), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT43), .B(G22gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n312), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n627), .B2(new_n628), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n258), .A2(new_n376), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n667), .A2(G29gat), .A3(new_n586), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(KEYINPUT94), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(KEYINPUT94), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n663), .B1(new_n590), .B2(new_n620), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n664), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n622), .A2(new_n623), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n673), .B(KEYINPUT44), .C1(new_n678), .C2(new_n663), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n679), .A3(new_n666), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n586), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n672), .A2(new_n681), .A3(new_n682), .ZN(G1328gat));
  OR3_X1    g482(.A1(new_n667), .A2(G36gat), .A3(new_n542), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT96), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n680), .A2(new_n542), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G36gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n689), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT96), .B1(new_n691), .B2(new_n685), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1329gat));
  NAND2_X1  g492(.A1(new_n658), .A2(G43gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n655), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n667), .A2(new_n695), .ZN(new_n696));
  OAI22_X1  g495(.A1(new_n680), .A2(new_n694), .B1(new_n696), .B2(G43gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g497(.A(G50gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n516), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n677), .A2(new_n679), .A3(new_n666), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT97), .B(KEYINPUT48), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n667), .B2(new_n516), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT98), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n701), .A2(new_n703), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT99), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT48), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n708), .B2(KEYINPUT48), .ZN(new_n711));
  OAI22_X1  g510(.A1(new_n706), .A2(new_n707), .B1(new_n710), .B2(new_n711), .ZN(G1331gat));
  AND4_X1   g511(.A1(new_n313), .A2(new_n626), .A3(new_n375), .A4(new_n344), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n633), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n541), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT100), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  AOI21_X1  g519(.A(G71gat), .B1(new_n713), .B2(new_n655), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n713), .A2(G71gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n658), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g523(.A1(new_n713), .A2(new_n618), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT101), .B(G78gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT102), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n725), .B(new_n727), .ZN(G1335gat));
  NAND2_X1  g527(.A1(new_n258), .A2(new_n344), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n677), .A2(new_n679), .A3(new_n375), .A4(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n731), .A2(new_n264), .A3(new_n586), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n674), .A2(new_n730), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT51), .ZN(new_n734));
  INV_X1    g533(.A(new_n375), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736), .B2(new_n633), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT103), .ZN(G1336gat));
  OAI21_X1  g538(.A(G92gat), .B1(new_n731), .B2(new_n542), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT104), .B(G92gat), .C1(new_n731), .C2(new_n542), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT51), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n542), .A2(G92gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n375), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n736), .A2(new_n746), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT106), .B(KEYINPUT52), .Z(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n731), .B2(new_n617), .ZN(new_n754));
  INV_X1    g553(.A(G99gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n755), .A3(new_n655), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1338gat));
  OAI21_X1  g556(.A(G106gat), .B1(new_n731), .B2(new_n516), .ZN(new_n758));
  INV_X1    g557(.A(new_n734), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n735), .A2(new_n516), .A3(G106gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n760), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(G1339gat));
  NAND3_X1  g566(.A1(new_n358), .A2(new_n364), .A3(new_n359), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n362), .A2(KEYINPUT54), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n364), .B1(new_n358), .B2(new_n359), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n373), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(KEYINPUT55), .A3(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n773), .A2(new_n312), .A3(new_n374), .ZN(new_n774));
  INV_X1    g573(.A(new_n317), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n334), .A2(new_n336), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n342), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n360), .A2(new_n771), .A3(new_n361), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n768), .A2(KEYINPUT54), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n371), .B(new_n780), .C1(new_n781), .C2(new_n770), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT55), .B1(new_n769), .B2(new_n772), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT108), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n774), .A2(new_n779), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n785), .B(KEYINPUT55), .C1(new_n769), .C2(new_n772), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT108), .B1(new_n782), .B2(new_n783), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n794), .A2(KEYINPUT109), .A3(new_n779), .A4(new_n774), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n343), .A2(new_n374), .A3(new_n773), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n797), .A2(new_n793), .A3(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n375), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n663), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n257), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n258), .A2(new_n312), .A3(new_n375), .A4(new_n343), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n588), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n542), .A2(new_n633), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n343), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(G113gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(G113gat), .ZN(new_n813));
  MUX2_X1   g612(.A(new_n810), .B(new_n812), .S(new_n813), .Z(G1340gat));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n375), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g615(.A1(new_n809), .A2(new_n257), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g617(.A1(new_n541), .A2(new_n663), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT111), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(G134gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n633), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT112), .Z(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n808), .B2(new_n663), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n633), .B1(new_n802), .B2(new_n803), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n516), .B1(new_n830), .B2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(G141gat), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n658), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n542), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n835), .B2(new_n344), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n807), .A2(new_n617), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT113), .Z(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n343), .B(new_n374), .C1(new_n784), .C2(KEYINPUT114), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n787), .B1(new_n841), .B2(new_n773), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n799), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n663), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n796), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n258), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n791), .A2(new_n795), .B1(new_n843), .B2(new_n663), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT115), .B1(new_n848), .B2(new_n257), .ZN(new_n849));
  INV_X1    g648(.A(new_n803), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n516), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n618), .B1(new_n802), .B2(new_n803), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n852), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n839), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT117), .B1(new_n857), .B2(new_n343), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n851), .A2(new_n853), .B1(new_n855), .B2(new_n852), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NOR4_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n344), .A4(new_n839), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n836), .B1(new_n862), .B2(G141gat), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n831), .A2(new_n834), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n832), .A3(new_n343), .A4(new_n542), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n832), .B1(new_n857), .B2(new_n343), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n828), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT118), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n835), .A2(new_n344), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT58), .B1(new_n870), .B2(new_n866), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n858), .A2(new_n861), .A3(new_n832), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n836), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n874), .ZN(G1344gat));
  NAND3_X1  g674(.A1(new_n773), .A2(new_n312), .A3(new_n374), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n792), .A3(new_n793), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n779), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n257), .B1(new_n880), .B2(new_n844), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n852), .B(new_n618), .C1(new_n881), .C2(new_n803), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n855), .A2(KEYINPUT57), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n375), .A3(new_n838), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT121), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n887), .A3(new_n375), .A4(new_n838), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(G148gat), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT59), .B1(new_n857), .B2(new_n375), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n889), .A2(new_n890), .B1(G148gat), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n831), .A2(new_n834), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n893), .A2(G148gat), .A3(new_n735), .A4(new_n541), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n892), .A2(new_n894), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n864), .A2(new_n257), .A3(new_n542), .ZN(new_n896));
  INV_X1    g695(.A(G155gat), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n258), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(new_n857), .B2(new_n898), .ZN(G1346gat));
  XNOR2_X1  g698(.A(KEYINPUT77), .B(G162gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n893), .B2(new_n820), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n857), .A2(new_n312), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n542), .A2(new_n633), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n805), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT123), .Z(new_n907));
  OAI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n344), .ZN(new_n908));
  INV_X1    g707(.A(new_n906), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n385), .A3(new_n343), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n909), .B2(new_n375), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n907), .A2(new_n735), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n907), .B2(new_n258), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n906), .A2(new_n258), .A3(new_n415), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT60), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n909), .A2(new_n392), .A3(new_n312), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n906), .B(KEYINPUT123), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n312), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(G190gat), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT61), .B(new_n392), .C1(new_n926), .C2(new_n312), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  AND2_X1   g729(.A1(new_n617), .A2(new_n905), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n884), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n343), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G197gat), .ZN(new_n934));
  INV_X1    g733(.A(new_n855), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n931), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(G197gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n344), .B2(new_n937), .ZN(G1352gat));
  NOR3_X1   g737(.A1(new_n936), .A2(G204gat), .A3(new_n735), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT62), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n884), .A2(new_n375), .A3(new_n931), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n370), .B2(new_n941), .ZN(G1353gat));
  INV_X1    g741(.A(new_n936), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n246), .A3(new_n257), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n932), .A2(new_n257), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  NAND3_X1  g747(.A1(new_n312), .A2(new_n475), .A3(new_n476), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT126), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n943), .A2(new_n312), .ZN(new_n953));
  INV_X1    g752(.A(G218gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT125), .B(G218gat), .C1(new_n943), .C2(new_n312), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1355gat));
endmodule


