//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT74), .A4(G104), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n191), .A2(KEYINPUT74), .A3(G104), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT4), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G101), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT75), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n190), .B1(new_n191), .B2(G104), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(KEYINPUT74), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n203), .B2(new_n192), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n197), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n199), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(KEYINPUT0), .B2(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n211), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n220), .A2(new_n211), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n208), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n211), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n214), .A2(new_n212), .B1(new_n217), .B2(new_n219), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n224), .B(KEYINPUT67), .C1(new_n225), .C2(new_n211), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n196), .A2(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n203), .A2(new_n200), .A3(new_n192), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n207), .A2(new_n223), .A3(new_n226), .A4(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G131), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n232));
  INV_X1    g046(.A(G134), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G137), .ZN(new_n234));
  INV_X1    g048(.A(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT11), .A3(G134), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT66), .A4(new_n237), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n231), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT65), .A2(G131), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT65), .A2(G131), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(new_n236), .A3(new_n237), .A4(new_n234), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n194), .A2(G107), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n191), .A2(G104), .ZN(new_n250));
  OAI21_X1  g064(.A(G101), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n220), .A2(new_n210), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n216), .A2(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n217), .A3(new_n219), .A4(KEYINPUT76), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT76), .B1(new_n258), .B2(new_n255), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n228), .B(new_n251), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT10), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n228), .A2(new_n251), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n220), .A2(new_n210), .B1(KEYINPUT1), .B2(new_n253), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n255), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n230), .A2(new_n248), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G140), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(G227), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n268), .B(new_n270), .Z(new_n271));
  AND2_X1   g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n248), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n199), .A2(new_n206), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n229), .A2(new_n223), .A3(new_n226), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n261), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n262), .A2(new_n265), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n273), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n264), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n254), .B1(new_n258), .B2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n228), .A2(new_n251), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n260), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n242), .B2(new_n247), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT12), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n260), .A2(new_n285), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT12), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n273), .A2(new_n290), .A3(new_n287), .A4(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n267), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n271), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n272), .A2(new_n280), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n189), .B1(new_n295), .B2(G469), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT72), .B(G902), .Z(new_n297));
  NAND4_X1  g111(.A1(new_n267), .A2(new_n289), .A3(new_n271), .A4(new_n292), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n271), .B1(new_n280), .B2(new_n267), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n187), .B(new_n297), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n297), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n230), .A2(new_n248), .A3(new_n266), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n248), .B1(new_n230), .B2(new_n266), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n294), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n304), .B1(new_n307), .B2(new_n298), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT78), .B1(new_n308), .B2(new_n187), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n296), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G210), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G116), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT2), .B(G113), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G113), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n326));
  INV_X1    g140(.A(new_n319), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G116), .B(G119), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n324), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n262), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n329), .B(new_n323), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n229), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n333), .B(new_n334), .C1(new_n274), .C2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n229), .A2(new_n336), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n339), .A2(new_n207), .B1(new_n262), .B2(new_n332), .ZN(new_n340));
  INV_X1    g154(.A(new_n334), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT80), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n338), .B(KEYINPUT6), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G125), .B1(new_n221), .B2(new_n222), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n281), .B2(new_n282), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n344), .B2(new_n346), .ZN(new_n349));
  INV_X1    g163(.A(G224), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G953), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n344), .A2(new_n346), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT81), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n333), .B1(new_n274), .B2(new_n337), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(KEYINPUT80), .A3(new_n360), .A4(new_n341), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n343), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n363));
  NOR2_X1   g177(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n353), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n344), .A2(new_n346), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT7), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n351), .A2(KEYINPUT85), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n351), .A2(KEYINPUT85), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n354), .A2(KEYINPUT86), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT86), .B1(new_n354), .B2(new_n370), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n338), .B(new_n366), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n374));
  OAI21_X1  g188(.A(G113), .B1(new_n330), .B2(new_n319), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT82), .B(G113), .C1(new_n330), .C2(new_n319), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n324), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n284), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n334), .B(KEYINPUT8), .ZN(new_n383));
  INV_X1    g197(.A(new_n331), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n381), .B1(new_n384), .B2(new_n375), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(new_n262), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n374), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n383), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n332), .B2(new_n284), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n375), .A2(new_n376), .B1(KEYINPUT5), .B2(new_n329), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n324), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n389), .B(KEYINPUT83), .C1(new_n284), .C2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n188), .B1(new_n373), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n317), .B1(new_n362), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n343), .A2(new_n358), .A3(new_n361), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n371), .A2(new_n372), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n392), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n338), .A4(new_n366), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n399), .A3(new_n188), .A4(new_n316), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n315), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n194), .ZN(new_n403));
  XNOR2_X1  g217(.A(G125), .B(G140), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n216), .ZN(new_n405));
  NOR2_X1   g219(.A1(G237), .A2(G953), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G214), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n218), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(G143), .A3(G214), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT18), .A2(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n406), .A2(G143), .A3(G214), .ZN(new_n412));
  AOI21_X1  g226(.A(G143), .B1(new_n406), .B2(G214), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT18), .B(G131), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT65), .B(G131), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n412), .B2(new_n413), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n245), .A3(new_n409), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G125), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n345), .A2(G140), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT16), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n345), .A2(KEYINPUT16), .A3(G140), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n216), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT17), .B(new_n416), .C1(new_n412), .C2(new_n413), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n425), .A3(G146), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n403), .B(new_n415), .C1(new_n420), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT87), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(new_n427), .A3(new_n429), .A4(new_n428), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n403), .A4(new_n415), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n403), .B1(new_n434), .B2(new_n415), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n188), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G475), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n432), .A2(new_n436), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n417), .A2(new_n418), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n404), .A2(KEYINPUT19), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n404), .A2(KEYINPUT19), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n443), .B(new_n429), .C1(new_n446), .C2(G146), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n415), .ZN(new_n448));
  INV_X1    g262(.A(new_n403), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT88), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT89), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n432), .A2(new_n436), .B1(new_n449), .B2(new_n448), .ZN(new_n458));
  INV_X1    g272(.A(new_n453), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n457), .B(KEYINPUT20), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n461), .A3(new_n453), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n441), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n218), .A2(G128), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n210), .A2(G143), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT91), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n466), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n233), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n320), .A2(G122), .ZN(new_n472));
  INV_X1    g286(.A(G122), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G116), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n474), .A3(new_n191), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n191), .B1(new_n472), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(new_n466), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n218), .A2(G128), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n466), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n233), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n469), .A2(new_n470), .A3(new_n233), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n210), .A2(G143), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT91), .B1(new_n486), .B2(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n488));
  AOI21_X1  g302(.A(G134), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(KEYINPUT14), .C1(new_n473), .C2(G116), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT14), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n320), .A3(G122), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n474), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n472), .B2(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g310(.A(G107), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n475), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT93), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n473), .B2(G116), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT92), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(new_n492), .A3(new_n474), .A4(new_n494), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n476), .B1(new_n502), .B2(G107), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n487), .A2(G134), .A3(new_n488), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n471), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n484), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G217), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n311), .A2(new_n509), .A3(G953), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT94), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n465), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n506), .B1(new_n503), .B2(new_n505), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n514), .A2(new_n515), .B1(new_n483), .B2(new_n478), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT95), .A3(new_n511), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n512), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n297), .ZN(new_n520));
  INV_X1    g334(.A(G478), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT15), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n519), .B(new_n297), .C1(KEYINPUT15), .C2(new_n521), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n269), .A2(G952), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(G234), .B2(G237), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n269), .B(new_n297), .C1(G234), .C2(G237), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n401), .A2(new_n464), .A3(new_n525), .A4(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT96), .B1(new_n313), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n312), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n301), .A2(new_n302), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n308), .A2(KEYINPUT78), .A3(new_n187), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n537), .B2(new_n296), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n523), .A2(new_n524), .A3(new_n531), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n457), .B1(new_n454), .B2(KEYINPUT20), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n460), .A2(new_n462), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n440), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n538), .A2(new_n539), .A3(new_n544), .A4(new_n401), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n533), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n221), .A2(new_n222), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT11), .B1(new_n235), .B2(G134), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n235), .A2(G134), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT66), .B1(new_n551), .B2(new_n236), .ZN(new_n552));
  INV_X1    g366(.A(new_n241), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n548), .B1(new_n554), .B2(new_n246), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n233), .A2(G137), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n556), .B2(new_n550), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n246), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n283), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n547), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n223), .B(new_n226), .C1(new_n242), .C2(new_n247), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n557), .B(new_n562), .C1(new_n238), .C2(new_n416), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n246), .B2(new_n557), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n564), .A2(new_n565), .B1(new_n281), .B2(new_n282), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n566), .A3(KEYINPUT30), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(new_n336), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n406), .A2(G210), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT27), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT26), .B(G101), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n561), .A2(new_n566), .A3(new_n335), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n568), .A2(KEYINPUT31), .A3(new_n572), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT28), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n248), .A2(new_n548), .B1(new_n283), .B2(new_n558), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n573), .A2(new_n579), .B1(new_n580), .B2(new_n336), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n561), .A2(new_n566), .A3(KEYINPUT28), .A4(new_n335), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(G472), .A2(G902), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(KEYINPUT69), .Z(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n587), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n561), .A2(new_n566), .A3(new_n335), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n335), .B1(new_n561), .B2(new_n566), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n594), .B(KEYINPUT28), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n561), .A2(new_n566), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n336), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n579), .B1(new_n599), .B2(new_n573), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT71), .B1(new_n573), .B2(new_n579), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n572), .A2(KEYINPUT29), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n297), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n573), .A2(new_n579), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n580), .A2(new_n336), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n572), .A3(new_n606), .A4(new_n582), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT29), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n572), .B1(new_n568), .B2(new_n573), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n589), .A2(new_n593), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT22), .B(G137), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT23), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n318), .B2(G128), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n618), .B(new_n619), .C1(G119), .C2(new_n210), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT73), .B(G110), .Z(new_n621));
  XNOR2_X1  g435(.A(G119), .B(G128), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT24), .B(G110), .Z(new_n623));
  OAI22_X1  g437(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n422), .A2(new_n423), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n624), .B(new_n429), .C1(G146), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n427), .A2(new_n429), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n620), .A2(G110), .B1(new_n622), .B2(new_n623), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n616), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n629), .A3(new_n616), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT25), .B1(new_n633), .B2(new_n304), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n509), .B1(new_n297), .B2(G234), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n304), .B1(new_n631), .B2(new_n632), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT25), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n635), .A2(G902), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n613), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n546), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G101), .ZN(G3));
  NOR2_X1   g461(.A1(new_n592), .A2(new_n587), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n585), .A2(new_n297), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(G472), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n538), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n516), .B2(new_n511), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n519), .A2(new_n652), .B1(new_n518), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n521), .B1(new_n654), .B2(new_n297), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n519), .A2(new_n521), .A3(new_n297), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT97), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n530), .B(new_n315), .C1(new_n395), .C2(new_n400), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  AOI221_X4 g474(.A(new_n304), .B1(new_n518), .B2(new_n653), .C1(new_n519), .C2(new_n652), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n660), .B(new_n656), .C1(new_n661), .C2(new_n521), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n658), .A2(new_n659), .A3(new_n543), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT34), .B(G104), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  AOI21_X1  g480(.A(new_n441), .B1(new_n523), .B2(new_n524), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n456), .A2(new_n463), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT98), .B1(new_n541), .B2(new_n542), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n659), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n651), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT35), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G107), .ZN(G9));
  NAND2_X1  g491(.A1(new_n626), .A2(new_n629), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n616), .A2(KEYINPUT36), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n634), .A2(new_n639), .B1(new_n641), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n650), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n546), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n527), .B1(new_n528), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n671), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n315), .B(new_n681), .C1(new_n395), .C2(new_n400), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n613), .A3(new_n538), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XOR2_X1   g506(.A(new_n688), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n538), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT40), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n395), .A2(new_n400), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  INV_X1    g511(.A(new_n574), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n572), .B1(new_n599), .B2(new_n573), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n188), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G472), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n589), .A2(new_n593), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n315), .B1(new_n523), .B2(new_n524), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n703), .A2(new_n543), .A3(new_n681), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n697), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n695), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT101), .B(G143), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G45));
  AND3_X1   g524(.A1(new_n538), .A2(new_n613), .A3(new_n690), .ZN(new_n711));
  INV_X1    g525(.A(new_n688), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n543), .A2(new_n658), .A3(new_n662), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  AND4_X1   g529(.A1(new_n543), .A2(new_n658), .A3(new_n659), .A4(new_n662), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n307), .A2(new_n298), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n187), .B1(new_n717), .B2(new_n297), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n534), .B(new_n718), .C1(new_n535), .C2(new_n536), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n716), .A2(new_n645), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT102), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n613), .A3(new_n644), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n673), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n320), .ZN(G18));
  NOR3_X1   g540(.A1(new_n540), .A2(new_n543), .A3(new_n681), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n719), .A3(new_n613), .A4(new_n401), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  INV_X1    g543(.A(new_n572), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n602), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n578), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n588), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT103), .B(G472), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n592), .B2(new_n304), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n733), .A2(new_n736), .A3(new_n644), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n703), .A2(new_n543), .A3(new_n696), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n719), .A4(new_n531), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  INV_X1    g554(.A(new_n718), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n401), .A2(new_n537), .A3(new_n312), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n733), .A2(new_n736), .A3(new_n682), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n713), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NAND2_X1  g560(.A1(new_n272), .A2(new_n280), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n293), .A2(new_n294), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n295), .A2(KEYINPUT104), .A3(G469), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n189), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n537), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n395), .A2(new_n314), .A3(new_n400), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n534), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT42), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT32), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n592), .B2(new_n587), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n589), .A2(new_n612), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n644), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT105), .B1(new_n760), .B2(new_n644), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n713), .B(new_n757), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n613), .A2(new_n754), .A3(new_n756), .A4(new_n644), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n658), .A2(new_n543), .A3(new_n662), .A4(new_n712), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n763), .A2(KEYINPUT106), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT106), .B1(new_n763), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  AND2_X1   g585(.A1(new_n754), .A2(new_n756), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n645), .A2(new_n772), .A3(new_n689), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(new_n755), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n295), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(G469), .ZN(new_n778));
  INV_X1    g592(.A(new_n189), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(G469), .C1(new_n777), .C2(G902), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n537), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n312), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n693), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n658), .A2(new_n464), .A3(new_n662), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT107), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(new_n650), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n682), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n775), .B(new_n785), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n235), .ZN(G39));
  NAND2_X1  g609(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n783), .A2(new_n312), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n766), .A2(new_n644), .A3(new_n613), .A4(new_n755), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT108), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND2_X1  g618(.A1(new_n537), .A2(new_n741), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n534), .A3(new_n755), .ZN(new_n806));
  INV_X1    g620(.A(new_n702), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n644), .A3(new_n527), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n658), .A2(new_n543), .A3(new_n662), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n788), .A2(new_n527), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n737), .ZN(new_n812));
  INV_X1    g626(.A(new_n742), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n526), .B(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n788), .A2(new_n527), .A3(new_n806), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT48), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n761), .A2(new_n762), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n816), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n719), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n697), .A3(new_n314), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n812), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n811), .A2(new_n737), .ZN(new_n827));
  INV_X1    g641(.A(new_n824), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n743), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n816), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n543), .B(new_n808), .C1(new_n658), .C2(new_n662), .ZN(new_n833));
  INV_X1    g647(.A(new_n800), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n537), .A2(new_n534), .A3(new_n741), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n755), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n833), .B1(new_n836), .B2(new_n812), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n830), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n812), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(KEYINPUT115), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(KEYINPUT51), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT51), .B1(new_n839), .B2(KEYINPUT115), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n832), .A3(new_n830), .A4(new_n837), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n822), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT111), .B1(new_n525), .B2(new_n543), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n809), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n658), .A2(KEYINPUT111), .A3(new_n662), .A4(new_n543), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n644), .A2(new_n538), .A3(new_n650), .A4(new_n659), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n533), .B(new_n545), .C1(new_n645), .C2(new_n683), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT110), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n739), .B(new_n728), .C1(new_n663), .C2(new_n724), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n725), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n727), .A2(new_n613), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n537), .A2(new_n312), .A3(new_n531), .A4(new_n741), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n703), .A2(new_n696), .A3(new_n543), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n856), .A2(new_n813), .B1(new_n859), .B2(new_n737), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n645), .A2(new_n672), .A3(new_n659), .A4(new_n719), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n720), .A3(new_n861), .A4(KEYINPUT110), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n852), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n681), .A2(KEYINPUT112), .A3(new_n712), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT112), .B1(new_n681), .B2(new_n712), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n534), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n738), .A3(new_n702), .A4(new_n754), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n714), .A2(new_n745), .A3(new_n691), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n711), .B1(new_n713), .B2(new_n689), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .A3(new_n745), .A4(new_n867), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n525), .A2(new_n440), .A3(new_n682), .A4(new_n712), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n755), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n669), .A2(new_n670), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n613), .A3(new_n538), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n773), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n713), .A2(new_n831), .A3(new_n772), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n770), .A2(new_n863), .A3(new_n873), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n852), .A2(new_n882), .A3(new_n878), .A4(new_n879), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n854), .A2(new_n725), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n763), .A2(new_n767), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n886), .A2(KEYINPUT113), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT113), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n885), .B(new_n873), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n883), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n881), .B(new_n882), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(KEYINPUT54), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n844), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT116), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n844), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  OR2_X1    g711(.A1(G952), .A2(G953), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n786), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n644), .A3(new_n312), .A4(new_n314), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT109), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n805), .B(KEYINPUT49), .Z(new_n905));
  NOR2_X1   g719(.A1(new_n697), .A2(new_n702), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n899), .A2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n269), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n297), .B1(new_n883), .B2(new_n890), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n911), .B2(new_n317), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n343), .A2(new_n361), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n358), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n910), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n912), .B2(new_n915), .ZN(G51));
  XNOR2_X1  g731(.A(new_n189), .B(KEYINPUT57), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n884), .B1(new_n883), .B2(new_n890), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n891), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n921), .A3(new_n717), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n911), .A2(G469), .A3(new_n777), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n920), .B2(new_n717), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n910), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(KEYINPUT118), .B(new_n910), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G54));
  AND3_X1   g744(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n910), .B1(new_n931), .B2(new_n451), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n451), .B2(new_n931), .ZN(G60));
  NOR2_X1   g747(.A1(new_n891), .A2(new_n919), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n654), .B(KEYINPUT119), .Z(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n910), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT120), .ZN(new_n940));
  INV_X1    g754(.A(new_n893), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(new_n883), .A2(new_n890), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT60), .B1(new_n509), .B2(new_n188), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n509), .A2(new_n188), .A3(KEYINPUT60), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n909), .B1(new_n947), .B2(new_n633), .ZN(new_n948));
  INV_X1    g762(.A(new_n680), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n947), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT61), .ZN(G66));
  OR3_X1    g766(.A1(new_n863), .A2(KEYINPUT122), .A3(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT122), .B1(new_n863), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n529), .B2(new_n350), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n913), .B1(G898), .B2(new_n269), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n560), .A2(new_n567), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n446), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT123), .Z(new_n961));
  NOR2_X1   g775(.A1(new_n694), .A2(new_n755), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n848), .A2(new_n645), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n803), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n794), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n871), .A2(new_n745), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n708), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  AND3_X1   g783(.A1(new_n964), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n961), .B1(new_n970), .B2(G953), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n785), .A2(new_n738), .A3(new_n819), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n972), .A2(new_n773), .A3(new_n967), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n803), .A2(new_n770), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n269), .B1(new_n974), .B2(new_n794), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n687), .A2(G953), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n960), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT124), .B1(new_n975), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n961), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n980), .B(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(new_n568), .A2(new_n573), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n572), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n964), .A2(new_n969), .A3(new_n965), .A4(new_n863), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  AOI21_X1  g804(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT126), .Z(new_n992));
  OR2_X1    g806(.A1(new_n974), .A2(new_n794), .ZN(new_n993));
  INV_X1    g807(.A(new_n863), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(new_n730), .A3(new_n573), .A4(new_n568), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n990), .B1(new_n698), .B2(new_n610), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n892), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n910), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n992), .A2(new_n1000), .ZN(G57));
endmodule


