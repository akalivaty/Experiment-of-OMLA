//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n207), .A2(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G97), .A2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n218), .B(new_n223), .C1(G58), .C2(G232), .ZN(new_n224));
  INV_X1    g0024(.A(new_n210), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  AOI211_X1 g0027(.A(new_n214), .B(new_n227), .C1(new_n213), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G226), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n217), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  INV_X1    g0039(.A(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n216), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT69), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n250));
  OAI21_X1  g0050(.A(G58), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT8), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n248), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT69), .B1(new_n255), .B2(G58), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n247), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n203), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n210), .B2(new_n246), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT71), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(new_n266), .A3(G13), .A4(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n267), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT70), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n261), .A2(new_n276), .A3(new_n263), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(new_n271), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n202), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n265), .A2(new_n275), .A3(new_n277), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n266), .A2(KEYINPUT67), .A3(G274), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n292), .B1(new_n240), .B2(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n262), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n289), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G226), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT67), .B1(new_n296), .B2(new_n262), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n208), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(G1), .B1(new_n283), .B2(new_n288), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n298), .B1(new_n299), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT72), .B1(new_n281), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n308), .A2(G179), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n290), .A2(G232), .A3(new_n291), .ZN(new_n315));
  INV_X1    g0115(.A(G107), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n315), .B1(new_n316), .B2(new_n290), .C1(new_n293), .C2(new_n222), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n297), .ZN(new_n318));
  INV_X1    g0118(.A(new_n289), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n305), .B1(new_n300), .B2(new_n303), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G244), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n318), .A2(G190), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n323), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n289), .B1(new_n317), .B2(new_n297), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n321), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n274), .A2(G77), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n279), .A2(new_n240), .ZN(new_n331));
  INV_X1    g0131(.A(new_n247), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  INV_X1    g0134(.A(new_n258), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n332), .A2(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G20), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n240), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n263), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n326), .A2(new_n329), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n308), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G190), .B2(new_n308), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT74), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n281), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n264), .A2(KEYINPUT70), .B1(new_n202), .B2(new_n279), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n349), .A2(KEYINPUT74), .A3(new_n275), .A4(new_n277), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n348), .A2(KEYINPUT9), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT9), .B1(new_n348), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT10), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n346), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  AOI211_X1 g0156(.A(new_n314), .B(new_n343), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT16), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT78), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT78), .A3(G33), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(G20), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n290), .B2(G20), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n221), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n252), .A2(new_n221), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n370), .B2(new_n201), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n335), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n358), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n375));
  INV_X1    g0175(.A(new_n263), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n362), .A2(G33), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n361), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n366), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n368), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n373), .B1(new_n380), .B2(G68), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n376), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT79), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n358), .C1(new_n369), .C2(new_n373), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n375), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n254), .A2(new_n256), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n273), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n279), .B2(new_n386), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT80), .ZN(new_n389));
  INV_X1    g0189(.A(G232), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n307), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n320), .A2(KEYINPUT80), .A3(G232), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n289), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n290), .A2(G226), .A3(G1698), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n290), .A2(G223), .A3(new_n291), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n297), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(G190), .A3(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n320), .A2(KEYINPUT80), .A3(G232), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT80), .B1(new_n320), .B2(G232), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n319), .B(new_n398), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G200), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n385), .A2(new_n388), .A3(new_n399), .A4(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n385), .A2(new_n388), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(G169), .ZN(new_n408));
  INV_X1    g0208(.A(G179), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n402), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT18), .B1(new_n407), .B2(new_n410), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n405), .A2(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n377), .A2(new_n361), .A3(G226), .A4(new_n291), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n377), .A2(new_n361), .A3(G232), .A4(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT75), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT75), .A4(new_n418), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n297), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n289), .B1(new_n320), .B2(G238), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n415), .B1(new_n428), .B2(G179), .ZN(new_n429));
  OAI21_X1  g0229(.A(G169), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n423), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n431), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(G169), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n429), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n272), .A2(G68), .A3(new_n267), .ZN(new_n440));
  XOR2_X1   g0240(.A(new_n440), .B(KEYINPUT76), .Z(new_n441));
  AOI22_X1  g0241(.A1(new_n247), .A2(G77), .B1(new_n258), .B2(G50), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n337), .B2(G68), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n263), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT11), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n279), .A2(new_n221), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT12), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n439), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n428), .A2(G190), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n436), .A2(G200), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n451), .A2(new_n452), .A3(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n328), .A2(new_n309), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n327), .A2(new_n409), .A3(new_n321), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n340), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n413), .A2(new_n450), .A3(new_n453), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n357), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n316), .A2(G20), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT23), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n377), .A2(new_n361), .A3(new_n337), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n290), .A2(new_n465), .A3(new_n337), .A4(G87), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n247), .A2(G116), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n263), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT81), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n246), .B2(G1), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n266), .A2(KEYINPUT81), .A3(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n278), .A2(new_n376), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n272), .A2(KEYINPUT82), .A3(new_n474), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n278), .A2(G107), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n482), .B(KEYINPUT25), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n377), .A2(new_n361), .A3(G250), .A4(new_n291), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT86), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT86), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n290), .A2(new_n487), .A3(G250), .A4(new_n291), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G294), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n297), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n266), .A2(G45), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n496), .C1(new_n287), .C2(KEYINPUT5), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G264), .A3(new_n304), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT66), .B(G41), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT5), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(new_n304), .A3(G274), .A4(new_n494), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G169), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT87), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n493), .A2(G179), .A3(new_n498), .A4(new_n502), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n484), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT88), .B(new_n484), .C1(new_n507), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n472), .A2(new_n481), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n486), .A2(new_n488), .A3(new_n491), .A4(new_n490), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n501), .A2(new_n494), .B1(new_n300), .B2(new_n303), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n297), .A2(new_n515), .B1(new_n516), .B2(G264), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G190), .A3(new_n502), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n503), .A2(G200), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n514), .A2(new_n483), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n497), .A2(G257), .A3(new_n304), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n521), .A2(new_n502), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n377), .A2(new_n361), .A3(G244), .A4(new_n291), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n291), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n297), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n409), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n480), .A2(G97), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n279), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT6), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n316), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n316), .A2(KEYINPUT6), .A3(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n258), .A2(G77), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n378), .A2(new_n337), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n542), .B(new_n543), .C1(new_n545), .C2(new_n316), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n263), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n533), .A2(new_n535), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n522), .A2(new_n530), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n309), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n532), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n344), .B1(new_n522), .B2(new_n530), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n480), .A2(G97), .B1(new_n546), .B2(new_n263), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n522), .A2(G190), .A3(new_n530), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n535), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n377), .A2(new_n361), .A3(G238), .A4(new_n291), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n377), .A2(new_n361), .A3(G244), .A4(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n297), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n282), .A2(new_n288), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n296), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n301), .B1(new_n208), .B2(new_n302), .ZN(new_n565));
  OAI211_X1 g0365(.A(G250), .B(new_n495), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G190), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n344), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n480), .A2(G87), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n337), .ZN(new_n573));
  INV_X1    g0373(.A(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n538), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n290), .A2(new_n337), .A3(G68), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n332), .B2(new_n534), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT83), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n578), .A2(new_n579), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n263), .B1(new_n279), .B2(new_n333), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n571), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n333), .B1(new_n478), .B2(new_n479), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n263), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n279), .A2(new_n333), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n586), .A2(new_n589), .B1(G179), .B2(new_n567), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n568), .A2(G169), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n570), .A2(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n269), .A2(new_n216), .A3(new_n271), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT85), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n269), .A2(KEYINPUT85), .A3(new_n216), .A4(new_n271), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n272), .A2(G116), .A3(new_n474), .A4(new_n475), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n528), .B(new_n337), .C1(G33), .C2(new_n534), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n216), .A2(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n263), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n599), .A2(new_n263), .A3(KEYINPUT20), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n377), .A2(new_n361), .A3(G264), .A4(G1698), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n377), .A2(new_n361), .A3(G257), .A4(new_n291), .ZN(new_n609));
  XOR2_X1   g0409(.A(KEYINPUT84), .B(G303), .Z(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n290), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n297), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n497), .A2(G270), .A3(new_n304), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n502), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  INV_X1    g0415(.A(G190), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n607), .B(new_n615), .C1(new_n616), .C2(new_n614), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n606), .A2(G169), .A3(new_n614), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n614), .A2(new_n409), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n606), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n606), .A2(new_n614), .A3(KEYINPUT21), .A4(G169), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n617), .A2(new_n620), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n557), .A2(new_n592), .A3(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n460), .A2(new_n513), .A3(new_n520), .A4(new_n625), .ZN(G372));
  NAND3_X1  g0426(.A1(new_n571), .A2(KEYINPUT90), .A3(new_n584), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT90), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n574), .B1(new_n478), .B2(new_n479), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n589), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT89), .B1(new_n566), .B2(new_n563), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n566), .A2(KEYINPUT89), .A3(new_n563), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n562), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n627), .A2(new_n630), .A3(new_n635), .A4(new_n569), .ZN(new_n636));
  INV_X1    g0436(.A(new_n333), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n480), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n584), .B1(new_n409), .B2(new_n568), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n309), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n504), .A2(new_n506), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n484), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n554), .A2(new_n535), .B1(new_n309), .B2(new_n549), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n552), .B1(G190), .B2(new_n531), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n533), .A2(new_n535), .A3(new_n547), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n647), .A2(new_n532), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n642), .A2(new_n646), .A3(new_n650), .A4(new_n520), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT26), .B1(new_n592), .B2(new_n551), .ZN(new_n652));
  INV_X1    g0452(.A(new_n551), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n641), .A4(new_n636), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n651), .A2(new_n652), .A3(new_n641), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n460), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n453), .A2(new_n456), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n450), .A2(new_n659), .B1(new_n405), .B2(new_n406), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n411), .A2(new_n412), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n354), .A2(new_n356), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n658), .B1(new_n662), .B2(new_n314), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n354), .A2(new_n356), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n314), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(KEYINPUT91), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(G369));
  INV_X1    g0470(.A(new_n643), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n268), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n266), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n607), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n671), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n624), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT92), .Z(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n484), .A2(new_n678), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n513), .A2(new_n520), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n509), .A2(new_n679), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT93), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT93), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n686), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n645), .A2(new_n678), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n643), .A2(new_n678), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n211), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n499), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n575), .A2(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n206), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT95), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n642), .A2(new_n653), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n711), .A2(KEYINPUT26), .B1(new_n639), .B2(new_n640), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n592), .A2(new_n551), .A3(KEYINPUT26), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n642), .A2(new_n520), .A3(new_n650), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n671), .B1(new_n511), .B2(new_n512), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n712), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n710), .B1(new_n716), .B2(new_n679), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n656), .A2(new_n679), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n513), .A2(new_n520), .A3(new_n625), .A4(new_n679), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT94), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n566), .A2(KEYINPUT89), .A3(new_n563), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n631), .ZN(new_n725));
  AOI21_X1  g0525(.A(G179), .B1(new_n725), .B2(new_n562), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n503), .A3(new_n549), .A4(new_n614), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n517), .A2(new_n568), .A3(new_n530), .A4(new_n522), .ZN(new_n729));
  INV_X1    g0529(.A(new_n621), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n517), .A2(new_n568), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT30), .A3(new_n531), .A4(new_n621), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT31), .B1(new_n734), .B2(new_n678), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n723), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n678), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(KEYINPUT94), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n722), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n709), .B1(new_n721), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n720), .A2(KEYINPUT95), .A3(new_n744), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n708), .B1(new_n748), .B2(G1), .ZN(G364));
  NAND3_X1  g0549(.A1(G20), .A2(G190), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n409), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G326), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n337), .A2(G190), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G179), .A3(G200), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT33), .B(G317), .Z(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n337), .A2(new_n409), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(new_n344), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n756), .B1(new_n763), .B2(G322), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n616), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n337), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n753), .A2(new_n409), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n753), .A2(new_n409), .A3(new_n344), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n290), .B(new_n770), .C1(G329), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n757), .A2(new_n616), .A3(new_n344), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G311), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n750), .A2(G179), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G303), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n764), .A2(new_n773), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n763), .A2(G58), .B1(G77), .B2(new_n775), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT98), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n771), .A2(new_n372), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  INV_X1    g0584(.A(new_n751), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n290), .B1(new_n754), .B2(new_n221), .C1(new_n202), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n768), .A2(new_n316), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n766), .A2(new_n534), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n781), .A2(new_n782), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n777), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n574), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n779), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n262), .B1(G20), .B2(new_n309), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n702), .A2(new_n290), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n207), .A2(G45), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n241), .C2(new_n288), .ZN(new_n801));
  INV_X1    g0601(.A(G355), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n290), .A2(new_n211), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(G116), .B2(new_n211), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n793), .A2(new_n794), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n266), .B1(new_n672), .B2(G45), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n703), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n797), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n805), .B(new_n808), .C1(new_n682), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n683), .A2(new_n684), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n810), .B1(new_n813), .B2(new_n808), .ZN(G396));
  INV_X1    g0614(.A(new_n754), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G150), .B1(G137), .B2(new_n751), .ZN(new_n816));
  INV_X1    g0616(.A(G143), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n372), .B2(new_n774), .C1(new_n762), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n768), .A2(new_n221), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n766), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n822), .A2(G58), .B1(new_n772), .B2(G132), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n378), .B1(new_n777), .B2(G50), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n819), .A2(new_n821), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n777), .A2(G107), .B1(new_n751), .B2(G303), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n216), .B2(new_n774), .C1(new_n769), .C2(new_n754), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n763), .B2(G294), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n574), .A2(new_n768), .B1(new_n771), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT99), .Z(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n378), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n825), .B1(new_n788), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n794), .A2(new_n795), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n833), .A2(new_n794), .B1(new_n240), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n456), .A2(new_n678), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n340), .A2(new_n678), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n342), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n838), .B2(new_n456), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n835), .B(new_n808), .C1(new_n839), .C2(new_n796), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n718), .B(new_n839), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n745), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(KEYINPUT100), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(KEYINPUT100), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n841), .A2(new_n745), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n840), .B1(new_n846), .B2(new_n808), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n735), .A2(new_n736), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n722), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n460), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT40), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n382), .B1(KEYINPUT16), .B2(new_n381), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n388), .ZN(new_n853));
  INV_X1    g0653(.A(new_n676), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n410), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n404), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n407), .A2(new_n410), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n407), .B2(new_n854), .ZN(new_n860));
  AOI211_X1 g0660(.A(KEYINPUT101), .B(new_n676), .C1(new_n385), .C2(new_n388), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n404), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n676), .B1(new_n852), .B2(new_n388), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n413), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n439), .A2(new_n449), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n451), .A2(new_n452), .A3(new_n448), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n449), .A2(new_n678), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n449), .B(new_n678), .C1(new_n453), .C2(new_n439), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n849), .A2(new_n839), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n851), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n862), .A2(new_n863), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n858), .A2(new_n404), .ZN(new_n880));
  INV_X1    g0680(.A(new_n863), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n880), .B(new_n881), .C1(new_n861), .C2(new_n860), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n860), .A2(new_n861), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n879), .A2(new_n882), .B1(new_n413), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n885));
  OAI21_X1  g0685(.A(new_n878), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n875), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n838), .A2(new_n456), .ZN(new_n888));
  INV_X1    g0688(.A(new_n836), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n886), .A2(new_n891), .A3(KEYINPUT40), .A4(new_n849), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n877), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n850), .B(new_n893), .Z(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(G330), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n656), .A2(new_n679), .A3(new_n839), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n889), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n875), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n898), .A2(new_n869), .B1(new_n661), .B2(new_n854), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT39), .B1(new_n867), .B2(new_n868), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT103), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n878), .B(new_n902), .C1(new_n884), .C2(new_n885), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(KEYINPUT39), .C1(new_n867), .C2(new_n868), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n870), .A2(new_n678), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n357), .B(new_n458), .C1(new_n717), .C2(new_n719), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n669), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n895), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n266), .B2(new_n672), .ZN(new_n913));
  OAI211_X1 g0713(.A(G20), .B(new_n208), .C1(new_n541), .C2(KEYINPUT35), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n216), .B(new_n914), .C1(KEYINPUT35), .C2(new_n541), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OAI21_X1  g0716(.A(G77), .B1(new_n252), .B2(new_n221), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n917), .A2(new_n206), .B1(G50), .B2(new_n221), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G1), .A3(new_n268), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n916), .A3(new_n919), .ZN(G367));
  INV_X1    g0720(.A(new_n808), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n378), .B1(new_n774), .B2(new_n769), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(G311), .B2(new_n751), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT46), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n777), .A2(G116), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n923), .B1(new_n924), .B2(new_n925), .C1(new_n926), .C2(new_n771), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n924), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n928), .B1(new_n534), .B2(new_n768), .C1(new_n316), .C2(new_n766), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n754), .A2(new_n767), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n762), .A2(new_n610), .ZN(new_n931));
  NOR4_X1   g0731(.A1(new_n927), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n290), .B1(new_n791), .B2(new_n252), .ZN(new_n933));
  INV_X1    g0733(.A(G137), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n240), .A2(new_n768), .B1(new_n771), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G50), .C2(new_n775), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n766), .A2(new_n221), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(G150), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n938), .B1(new_n817), .B2(new_n785), .C1(new_n762), .C2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n815), .A2(G159), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n932), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT47), .Z(new_n946));
  AOI21_X1  g0746(.A(new_n921), .B1(new_n946), .B2(new_n794), .ZN(new_n947));
  INV_X1    g0747(.A(new_n799), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n798), .B1(new_n211), .B2(new_n333), .C1(new_n236), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n627), .A2(new_n630), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n678), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n642), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n641), .B2(new_n951), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n947), .B(new_n949), .C1(new_n809), .C2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n806), .B(KEYINPUT108), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n650), .B1(new_n649), .B2(new_n679), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n653), .A2(new_n678), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n699), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n691), .B2(new_n693), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n959), .B1(new_n961), .B2(new_n698), .ZN(new_n962));
  AND2_X1   g0762(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n959), .B(new_n966), .C1(new_n961), .C2(new_n698), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT45), .B1(new_n700), .B2(new_n958), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n688), .A2(new_n692), .A3(new_n689), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n692), .B1(new_n688), .B2(new_n689), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n699), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n698), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n958), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n964), .B(new_n967), .C1(new_n968), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n696), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n973), .A2(new_n974), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n978), .A2(new_n979), .B1(new_n963), .B2(new_n962), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n697), .A3(new_n967), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n691), .A2(new_n693), .A3(new_n960), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n971), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n686), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n685), .A2(new_n971), .A3(new_n982), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n746), .B2(new_n747), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n977), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n748), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n703), .B(KEYINPUT41), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n955), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT106), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n699), .B(new_n958), .C1(new_n969), .C2(new_n970), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(KEYINPUT42), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT42), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n961), .A2(KEYINPUT106), .A3(new_n995), .A4(new_n958), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n513), .A2(new_n956), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n678), .B1(new_n999), .B2(new_n551), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT105), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT105), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n997), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n696), .A2(new_n958), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n953), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT43), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1006), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1004), .B1(new_n998), .B2(new_n1001), .ZN(new_n1013));
  AOI211_X1 g0813(.A(KEYINPUT105), .B(new_n1000), .C1(new_n993), .C2(KEYINPUT42), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n994), .B(new_n996), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1011), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1012), .A2(new_n1017), .B1(KEYINPUT43), .B2(new_n953), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1008), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1015), .A2(new_n1007), .A3(new_n1016), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1019), .A2(new_n1010), .A3(new_n1009), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n954), .B1(new_n991), .B2(new_n1022), .ZN(G387));
  NAND3_X1  g0823(.A1(new_n748), .A2(new_n985), .A3(new_n984), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n746), .A2(new_n986), .A3(new_n747), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n703), .A3(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n815), .A2(G311), .B1(G322), .B2(new_n751), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n610), .B2(new_n774), .C1(new_n762), .C2(new_n926), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n769), .B2(new_n766), .C1(new_n767), .C2(new_n791), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT49), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n290), .B1(new_n772), .B2(G326), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n216), .C2(new_n768), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n768), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(G97), .B1(new_n772), .B2(G150), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n333), .B2(new_n766), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n762), .A2(new_n202), .B1(new_n372), .B2(new_n785), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT110), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n386), .A2(new_n754), .B1(new_n221), .B2(new_n774), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1036), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n1038), .B2(new_n1039), .C1(new_n240), .C2(new_n791), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1033), .B1(new_n378), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n799), .B1(new_n233), .B2(new_n288), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n705), .B2(new_n803), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G116), .B(new_n575), .C1(G68), .C2(G77), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n334), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT50), .B1(new_n334), .B2(G50), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1045), .A2(new_n288), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(G107), .B2(new_n211), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1042), .A2(new_n794), .B1(new_n798), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n808), .C1(new_n694), .C2(new_n809), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n955), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1026), .B(new_n1052), .C1(new_n986), .C2(new_n1053), .ZN(G393));
  NOR2_X1   g0854(.A1(new_n976), .A2(new_n696), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n697), .B1(new_n980), .B2(new_n967), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1024), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n703), .A3(new_n988), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n977), .A2(new_n981), .A3(new_n955), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n762), .A2(new_n829), .B1(new_n926), .B2(new_n785), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n290), .B1(new_n777), .B2(G283), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n767), .B2(new_n774), .C1(new_n610), .C2(new_n754), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n787), .B(new_n1063), .C1(G322), .C2(new_n772), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(new_n216), .C2(new_n766), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT113), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n762), .A2(new_n372), .B1(new_n939), .B2(new_n785), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n378), .B1(new_n777), .B2(G68), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n574), .B2(new_n768), .C1(new_n817), .C2(new_n771), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(KEYINPUT112), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n766), .A2(new_n240), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n754), .A2(new_n202), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n1070), .C2(KEYINPUT112), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1068), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n334), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n775), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n794), .B1(new_n1066), .B2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n798), .B1(new_n534), .B2(new_n211), .C1(new_n244), .C2(new_n948), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n808), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT111), .Z(new_n1081));
  OAI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(new_n809), .C2(new_n958), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1058), .A2(new_n1059), .A3(new_n1082), .ZN(G390));
  INV_X1    g0883(.A(new_n907), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n898), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1085), .A2(new_n903), .A3(new_n901), .A4(new_n905), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n716), .A2(new_n679), .A3(new_n888), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n889), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n875), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n886), .A2(new_n1084), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n340), .B1(new_n324), .B2(new_n325), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1093), .A2(new_n329), .B1(new_n340), .B2(new_n678), .ZN(new_n1094));
  OAI211_X1 g0894(.A(G330), .B(new_n889), .C1(new_n1094), .C2(new_n457), .ZN(new_n1095));
  AOI221_X4 g0895(.A(new_n1095), .B1(new_n873), .B2(new_n874), .C1(new_n722), .C2(new_n848), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1095), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n743), .A2(new_n875), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1086), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n357), .A2(G330), .A3(new_n458), .A4(new_n849), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n669), .A2(new_n909), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n875), .B1(new_n849), .B2(new_n1099), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1088), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n875), .B1(new_n743), .B2(new_n1099), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n897), .B1(new_n1106), .B2(new_n1096), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT114), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT114), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n897), .C1(new_n1106), .C2(new_n1096), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1105), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1098), .B(new_n1101), .C1(new_n1103), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1105), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1103), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1086), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1096), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n703), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n955), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n774), .A2(new_n534), .B1(new_n754), .B2(new_n316), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n763), .B2(G116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n751), .A2(G283), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n820), .B(new_n1072), .C1(G294), .C2(new_n772), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n792), .A2(new_n290), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n791), .A2(new_n939), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT53), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n290), .B1(new_n754), .B2(new_n934), .C1(new_n1130), .C2(new_n785), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G125), .C2(new_n772), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n766), .A2(new_n372), .B1(new_n768), .B2(new_n202), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n763), .A2(G132), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n774), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1126), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n794), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n921), .B1(new_n386), .B2(new_n834), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT115), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(new_n906), .C2(new_n796), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1119), .A2(new_n1120), .A3(new_n1144), .ZN(G378));
  NAND3_X1  g0945(.A1(new_n877), .A2(G330), .A3(new_n892), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n348), .A2(new_n350), .A3(new_n854), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT55), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n664), .B2(new_n667), .ZN(new_n1151));
  AOI211_X1 g0951(.A(KEYINPUT55), .B(new_n314), .C1(new_n354), .C2(new_n356), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n348), .A2(new_n350), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT9), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n348), .A2(KEYINPUT9), .A3(new_n350), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n355), .B1(new_n1158), .B2(new_n346), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n356), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n667), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT55), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n664), .A2(new_n1150), .A3(new_n667), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1149), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1146), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1146), .A2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n908), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n906), .A2(new_n907), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n899), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n877), .A2(G330), .A3(new_n892), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1146), .A2(new_n1166), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1172), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1169), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n955), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n834), .A2(new_n202), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n751), .A2(G125), .ZN(new_n1181));
  INV_X1    g0981(.A(G132), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n754), .C1(new_n791), .C2(new_n1138), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G150), .B2(new_n822), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n1130), .B2(new_n762), .C1(new_n934), .C2(new_n774), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n772), .A2(G124), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G33), .B(G41), .C1(new_n1034), .C2(G159), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n287), .A2(new_n378), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n774), .A2(new_n333), .B1(new_n754), .B2(new_n534), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n763), .B2(G107), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n252), .A2(new_n768), .B1(new_n771), .B2(new_n769), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n791), .A2(new_n240), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1195), .A2(new_n937), .A3(new_n1196), .A4(new_n1191), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1194), .B(new_n1197), .C1(new_n216), .C2(new_n785), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1199));
  XNOR2_X1  g0999(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1190), .A2(new_n1192), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n921), .B1(new_n1201), .B2(new_n794), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1180), .B(new_n1202), .C1(new_n1166), .C2(new_n796), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1179), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1103), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1118), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT118), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1172), .A2(new_n1175), .A3(new_n1207), .A4(new_n1176), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1169), .A2(new_n1177), .A3(KEYINPUT118), .ZN(new_n1209));
  AND4_X1   g1009(.A1(KEYINPUT57), .A2(new_n1206), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1118), .A2(new_n1205), .B1(new_n1177), .B2(new_n1169), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n703), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1210), .B2(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n887), .A2(new_n795), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n252), .A2(new_n768), .B1(new_n771), .B2(new_n1130), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n290), .B1(new_n774), .B2(new_n939), .C1(new_n372), .C2(new_n791), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G50), .C2(new_n822), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT120), .Z(new_n1218));
  AOI22_X1  g1018(.A1(new_n763), .A2(G137), .B1(G132), .B2(new_n751), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n754), .C2(new_n1138), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n774), .A2(new_n316), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n772), .A2(G303), .B1(G97), .B2(new_n777), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT119), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n378), .B1(new_n754), .B2(new_n216), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n766), .A2(new_n333), .B1(new_n768), .B2(new_n240), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(G294), .C2(new_n751), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1223), .B(new_n1226), .C1(new_n769), .C2(new_n762), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1220), .B1(new_n1221), .B2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1228), .A2(new_n794), .B1(new_n221), .B2(new_n834), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1214), .A2(new_n808), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1111), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n955), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1111), .A2(new_n1103), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n990), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1115), .ZN(G381));
  NOR4_X1   g1035(.A1(G375), .A2(G384), .A3(G378), .A4(G381), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n990), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n988), .B2(new_n748), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1021), .B(new_n1018), .C1(new_n1238), .C2(new_n955), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n954), .A3(new_n1239), .A4(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n677), .A2(G213), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT121), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OR3_X1    g1044(.A1(G375), .A2(G378), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G407), .A2(G213), .A3(new_n1245), .ZN(G409));
  NAND3_X1  g1046(.A1(new_n1206), .A2(new_n990), .A3(new_n1178), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1209), .A2(new_n955), .A3(new_n1208), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1203), .A3(new_n1248), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1119), .A2(new_n1120), .A3(new_n1144), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT122), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1204), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(KEYINPUT122), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n704), .B1(new_n1233), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1115), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n1257), .C2(new_n1233), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(G384), .A3(new_n1232), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1260), .B2(new_n1232), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1256), .A2(new_n1244), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT125), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1256), .A2(new_n1244), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1243), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1263), .B(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1256), .A2(new_n1244), .A3(new_n1263), .A4(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1267), .A2(new_n1272), .A3(new_n1273), .A4(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1239), .A2(G390), .A3(new_n954), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G390), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1277), .ZN(new_n1282));
  XOR2_X1   g1082(.A(G393), .B(G396), .Z(new_n1283));
  AOI21_X1  g1083(.A(new_n1279), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1281), .A3(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1244), .A4(new_n1263), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1264), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1290), .B(new_n1291), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT126), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(G405));
  AND2_X1   g1100(.A1(new_n1288), .A2(KEYINPUT127), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1287), .B(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1250), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1254), .ZN(new_n1304));
  XOR2_X1   g1104(.A(new_n1304), .B(new_n1263), .Z(new_n1305));
  MUX2_X1   g1105(.A(new_n1301), .B(new_n1302), .S(new_n1305), .Z(G402));
endmodule


