//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(G116), .B(G119), .Z(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(new_n190), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(new_n202), .A3(new_n206), .A4(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n213), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(new_n213), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n208), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n210), .A3(new_n212), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n209), .A3(G143), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n211), .B(G146), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g044(.A(G134), .B(G137), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n206), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n199), .A2(G137), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n201), .A2(G134), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT66), .B(G131), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n229), .A2(new_n232), .A3(new_n207), .A4(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n197), .B1(new_n223), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n225), .A2(new_n210), .A3(new_n212), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(new_n227), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n226), .A2(new_n241), .A3(new_n227), .A4(new_n228), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n232), .A2(new_n207), .A3(new_n235), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n215), .A2(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n243), .A2(new_n244), .B1(new_n245), .B2(new_n208), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n237), .B1(new_n197), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT68), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n244), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n223), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n197), .B1(new_n251), .B2(KEYINPUT69), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n248), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n251), .A2(new_n196), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n256), .B(KEYINPUT28), .C1(new_n257), .C2(new_n237), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n249), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n223), .A2(new_n236), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n250), .A2(KEYINPUT30), .A3(new_n223), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n196), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n246), .A2(new_n197), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n264), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n271), .A2(KEYINPUT31), .A3(new_n272), .A4(new_n264), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n189), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT71), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n259), .A2(new_n265), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  NOR4_X1   g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .A4(new_n189), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n251), .A2(new_n196), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n272), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT28), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n255), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n271), .A2(new_n272), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n264), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n259), .B2(new_n264), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(KEYINPUT29), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT70), .B(new_n282), .C1(new_n280), .C2(new_n189), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n284), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n301), .B(KEYINPUT81), .Z(new_n302));
  INV_X1    g116(.A(KEYINPUT83), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G116), .ZN(new_n306));
  OAI211_X1 g120(.A(G113), .B(new_n306), .C1(new_n194), .C2(new_n304), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n307), .A2(new_n193), .ZN(new_n308));
  INV_X1    g122(.A(G107), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT75), .A3(G104), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n309), .A2(G104), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G101), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(new_n309), .A3(KEYINPUT75), .A4(G104), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n311), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G104), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT76), .A3(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n318), .B2(G107), .ZN(new_n321));
  OAI211_X1 g135(.A(G101), .B(new_n319), .C1(new_n321), .C2(new_n312), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n317), .A2(KEYINPUT77), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT77), .B1(new_n317), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n308), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n311), .A2(new_n313), .A3(new_n316), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n317), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n330), .A3(G101), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n331), .A3(new_n196), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n326), .B1(new_n325), .B2(new_n332), .ZN(new_n334));
  XOR2_X1   g148(.A(G110), .B(G122), .Z(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n332), .A3(new_n336), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT6), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n303), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n229), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n245), .B2(new_n342), .ZN(new_n344));
  INV_X1    g158(.A(G953), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(G224), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n325), .A2(new_n332), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT82), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n325), .A2(new_n332), .A3(new_n326), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n335), .ZN(new_n353));
  INV_X1    g167(.A(new_n339), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT83), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n340), .A2(new_n347), .A3(new_n349), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G210), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n344), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT7), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n346), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT84), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n307), .A2(new_n193), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n317), .A2(new_n322), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n335), .B(KEYINPUT8), .Z(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT85), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n358), .A2(new_n367), .A3(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n344), .B(new_n369), .C1(new_n359), .C2(new_n346), .ZN(new_n370));
  AND4_X1   g184(.A1(new_n361), .A2(new_n366), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n338), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n367), .B1(new_n358), .B2(new_n360), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n356), .A2(new_n357), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n357), .B1(new_n356), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n302), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n342), .A2(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n382), .B(KEYINPUT19), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n209), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT90), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n345), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n211), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n206), .A3(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT16), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G146), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n396), .B(KEYINPUT74), .Z(new_n397));
  INV_X1    g211(.A(KEYINPUT90), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n383), .A2(new_n398), .A3(new_n209), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n385), .A2(new_n393), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n382), .A2(G146), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n380), .A2(new_n381), .A3(new_n209), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(KEYINPUT87), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n382), .A2(new_n404), .A3(G146), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n387), .A2(new_n211), .ZN(new_n409));
  AOI21_X1  g223(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n390), .A2(KEYINPUT86), .A3(new_n408), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n390), .B2(new_n408), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n388), .A2(KEYINPUT88), .A3(new_n389), .A4(new_n407), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT89), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n403), .A2(new_n405), .ZN(new_n422));
  AND4_X1   g236(.A1(KEYINPUT89), .A2(new_n421), .A3(new_n422), .A4(new_n419), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n400), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G113), .B(G122), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(new_n318), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT17), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n429), .B(new_n206), .C1(new_n388), .C2(new_n389), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n396), .A2(KEYINPUT73), .ZN(new_n432));
  AOI21_X1  g246(.A(G146), .B1(new_n394), .B2(new_n395), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n394), .A2(new_n395), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT73), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n209), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n431), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n209), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(KEYINPUT73), .A3(new_n396), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT91), .A3(new_n431), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n415), .A2(KEYINPUT89), .A3(new_n419), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n421), .A2(new_n422), .A3(new_n419), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n453), .A3(new_n426), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n428), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G475), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n188), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT20), .ZN(new_n458));
  AOI21_X1  g272(.A(G475), .B1(new_n428), .B2(new_n454), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n188), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n454), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n426), .B1(new_n448), .B2(new_n453), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n188), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G475), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT92), .B1(new_n224), .B2(G143), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n211), .A3(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n211), .A2(G128), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(KEYINPUT95), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(G134), .A3(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n474), .B(new_n471), .C1(new_n467), .C2(new_n469), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT95), .B1(new_n470), .B2(new_n472), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n199), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G116), .B(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n309), .ZN(new_n483));
  INV_X1    g297(.A(G116), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT14), .A3(G122), .ZN(new_n485));
  INV_X1    g299(.A(new_n482), .ZN(new_n486));
  OAI211_X1 g300(.A(G107), .B(new_n485), .C1(new_n486), .C2(KEYINPUT14), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n481), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n491), .B2(new_n470), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n471), .B1(new_n491), .B2(new_n470), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n490), .A2(KEYINPUT94), .A3(new_n467), .A4(new_n469), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G134), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n486), .A2(G107), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n483), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n480), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT9), .B(G234), .Z(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(G217), .A3(new_n345), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n502), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n488), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n188), .ZN(new_n507));
  INV_X1    g321(.A(G478), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n503), .B2(new_n505), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(KEYINPUT15), .B2(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(G234), .A2(G237), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(G952), .A3(new_n345), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT21), .B(G898), .Z(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(G902), .A3(G953), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n462), .A2(new_n466), .A3(new_n514), .A4(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n378), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n229), .A2(new_n317), .A3(new_n322), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT79), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n341), .A3(new_n363), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n363), .A2(new_n341), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT79), .A3(new_n522), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT80), .ZN(new_n527));
  OR3_X1    g341(.A1(new_n527), .A2(KEYINPUT78), .A3(KEYINPUT12), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n523), .B(new_n525), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n208), .B(new_n529), .C1(new_n530), .C2(new_n527), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT10), .B(new_n243), .C1(new_n323), .C2(new_n324), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n329), .A2(new_n245), .A3(new_n331), .ZN(new_n533));
  INV_X1    g347(.A(new_n208), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT10), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G140), .ZN(new_n538));
  INV_X1    g352(.A(G227), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n538), .B(new_n540), .Z(new_n541));
  NOR2_X1   g355(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n524), .A2(new_n526), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT12), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n531), .A2(new_n537), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n208), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n537), .ZN(new_n548));
  INV_X1    g362(.A(new_n541), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n188), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n188), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n531), .A2(new_n537), .A3(new_n544), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n549), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n547), .A2(new_n537), .A3(new_n541), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(G469), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G221), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n501), .B2(new_n188), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT23), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n305), .B2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n224), .A2(G119), .ZN(new_n568));
  MUX2_X1   g382(.A(new_n566), .B(new_n567), .S(new_n568), .Z(new_n569));
  INV_X1    g383(.A(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(G119), .B(G128), .Z(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT24), .B(G110), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n397), .A2(new_n402), .A3(new_n575), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n569), .A2(new_n570), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n572), .A2(new_n573), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n443), .A4(new_n437), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT22), .B(G137), .ZN(new_n581));
  INV_X1    g395(.A(G234), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n561), .A2(new_n582), .A3(G953), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n581), .B(new_n583), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(new_n579), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n188), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT25), .ZN(new_n589));
  OAI21_X1  g403(.A(G217), .B1(new_n582), .B2(G902), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT72), .Z(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n586), .A2(new_n592), .A3(new_n188), .A4(new_n587), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n586), .A2(new_n587), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n591), .A2(G902), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n300), .A2(new_n521), .A3(new_n565), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NOR2_X1   g415(.A1(new_n511), .A2(G478), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT33), .B1(new_n503), .B2(new_n505), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n505), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n488), .A2(new_n499), .A3(KEYINPUT97), .A4(new_n504), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n488), .A2(new_n499), .A3(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n502), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT96), .B1(new_n488), .B2(new_n499), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT98), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n611), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n502), .A3(new_n609), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n607), .A3(new_n616), .A4(KEYINPUT33), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n603), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n508), .A2(G902), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n602), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n458), .A2(new_n461), .B1(G475), .B2(new_n465), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT99), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n301), .B(new_n519), .C1(new_n376), .C2(new_n377), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n459), .A2(new_n460), .A3(new_n188), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n460), .B1(new_n459), .B2(new_n188), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n466), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n619), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n603), .B(new_n629), .C1(new_n613), .C2(new_n617), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n625), .B(new_n628), .C1(new_n630), .C2(new_n602), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n622), .A2(new_n624), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n278), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n280), .B2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n564), .A2(new_n635), .A3(new_n598), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT91), .B1(new_n444), .B2(new_n431), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n440), .B(new_n430), .C1(new_n443), .C2(new_n437), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n446), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n420), .A2(new_n423), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n427), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n645), .B2(new_n454), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n640), .B1(new_n646), .B2(new_n456), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n465), .A2(KEYINPUT100), .A3(G475), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n462), .A3(new_n513), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n519), .B(KEYINPUT101), .Z(new_n651));
  AND2_X1   g465(.A1(new_n599), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n564), .A2(new_n635), .ZN(new_n654));
  INV_X1    g468(.A(new_n301), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n356), .A2(new_n375), .ZN(new_n656));
  INV_X1    g470(.A(new_n357), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n356), .A2(new_n357), .A3(new_n375), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n580), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n596), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n594), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n521), .A2(new_n654), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AOI21_X1  g489(.A(new_n564), .B1(new_n671), .B2(new_n669), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n300), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n678));
  OR3_X1    g492(.A1(new_n518), .A2(KEYINPUT103), .A3(G900), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT103), .B1(new_n518), .B2(G900), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n516), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n650), .A2(new_n660), .A3(KEYINPUT104), .A4(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n649), .A2(new_n462), .A3(new_n513), .A4(new_n681), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n301), .B1(new_n376), .B2(new_n377), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n677), .A2(new_n678), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n300), .A2(new_n676), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT105), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(G128), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G30));
  NAND2_X1  g507(.A1(new_n291), .A2(new_n264), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n264), .B2(new_n286), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n695), .B2(KEYINPUT107), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(KEYINPUT107), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G472), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n284), .A2(new_n299), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n667), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n681), .B(KEYINPUT39), .Z(new_n702));
  NOR2_X1   g516(.A1(new_n564), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT40), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n658), .A2(new_n659), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT38), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n621), .A2(new_n655), .A3(new_n514), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n701), .A2(new_n704), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  OAI211_X1 g523(.A(new_n628), .B(new_n681), .C1(new_n630), .C2(new_n602), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT108), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n613), .A2(new_n617), .ZN(new_n712));
  INV_X1    g526(.A(new_n603), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n619), .ZN(new_n714));
  INV_X1    g528(.A(new_n602), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n628), .A4(new_n681), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n677), .A3(KEYINPUT109), .A4(new_n660), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n711), .A2(new_n718), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n300), .A2(new_n676), .A3(new_n660), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  AND2_X1   g540(.A1(new_n300), .A2(new_n599), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n551), .A2(new_n188), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n563), .A3(new_n553), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n632), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NOR2_X1   g548(.A1(new_n685), .A2(new_n730), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n300), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n653), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  INV_X1    g552(.A(new_n520), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n739), .A3(new_n672), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  AND2_X1   g555(.A1(new_n707), .A2(new_n705), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n277), .B1(new_n288), .B2(new_n264), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n187), .A3(new_n188), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n634), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n730), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n652), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n668), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n711), .A2(new_n718), .A3(new_n735), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n342), .ZN(G27));
  OR2_X1    g565(.A1(new_n558), .A2(KEYINPUT110), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n558), .A2(KEYINPUT110), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n557), .A2(new_n752), .A3(G469), .A4(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n553), .A3(new_n555), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n563), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n658), .A2(new_n659), .A3(new_n301), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n300), .A2(new_n599), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n719), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n758), .A2(new_n756), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n294), .A2(G472), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n633), .A2(new_n282), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n598), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n711), .A2(new_n718), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT42), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n206), .ZN(G33));
  OR2_X1    g585(.A1(new_n760), .A2(new_n684), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n716), .A2(new_n621), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n635), .A3(new_n667), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n759), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n557), .A2(new_n752), .A3(KEYINPUT45), .A4(new_n753), .ZN(new_n784));
  INV_X1    g598(.A(new_n558), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n556), .B2(new_n549), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n784), .B(G469), .C1(KEYINPUT45), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n555), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n553), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT46), .B1(new_n787), .B2(new_n555), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n563), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(new_n702), .ZN(new_n792));
  OR3_X1    g606(.A1(new_n782), .A2(new_n783), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NAND2_X1  g608(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n796), .B(new_n563), .C1(new_n789), .C2(new_n790), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n300), .A2(new_n599), .A3(new_n758), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n795), .A2(new_n719), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n801));
  NOR2_X1   g615(.A1(G952), .A2(G953), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n719), .A2(new_n749), .A3(new_n764), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n763), .A2(new_n772), .A3(new_n769), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n620), .A2(new_n621), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n302), .B(new_n651), .C1(new_n376), .C2(new_n377), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n636), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n600), .A2(new_n673), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n621), .A2(KEYINPUT113), .A3(new_n513), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n466), .B(new_n513), .C1(new_n626), .C2(new_n627), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n807), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n636), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n809), .A2(new_n740), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n732), .A2(new_n737), .A3(new_n747), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n649), .A2(new_n462), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n676), .A2(new_n822), .A3(new_n681), .A4(new_n759), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n300), .A2(new_n514), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n804), .A2(new_n820), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n699), .A2(new_n668), .A3(new_n681), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n707), .A2(new_n705), .A3(new_n757), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n750), .B(new_n829), .C1(new_n687), .C2(new_n690), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n830), .B2(new_n725), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n750), .B1(new_n687), .B2(new_n690), .ZN(new_n832));
  INV_X1    g646(.A(new_n829), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n725), .A3(KEYINPUT52), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n826), .B(KEYINPUT53), .C1(new_n831), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  INV_X1    g653(.A(new_n750), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n682), .A2(new_n686), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n678), .B1(new_n841), .B2(new_n677), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT105), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n840), .B(new_n833), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n720), .A2(new_n724), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n839), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n834), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(KEYINPUT116), .A3(KEYINPUT53), .A4(new_n826), .ZN(new_n848));
  INV_X1    g662(.A(new_n804), .ZN(new_n849));
  INV_X1    g663(.A(new_n821), .ZN(new_n850));
  INV_X1    g664(.A(new_n820), .ZN(new_n851));
  INV_X1    g665(.A(new_n825), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n691), .A2(new_n840), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n829), .A2(new_n839), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n832), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n855), .A2(new_n725), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n853), .B1(new_n859), .B2(new_n846), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n838), .B(new_n848), .C1(KEYINPUT53), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n847), .B2(new_n826), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(KEYINPUT53), .B2(new_n860), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n861), .A2(KEYINPUT54), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n745), .A2(new_n598), .A3(new_n516), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n779), .A2(new_n731), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n706), .A2(new_n301), .ZN(new_n870));
  OR2_X1    g684(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n868), .A2(new_n301), .A3(new_n706), .ZN(new_n873));
  XOR2_X1   g687(.A(KEYINPUT119), .B(KEYINPUT50), .Z(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n779), .A2(new_n867), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n729), .A2(new_n553), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT118), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n563), .B1(new_n879), .B2(KEYINPUT118), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n795), .A2(new_n797), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n878), .A2(new_n882), .A3(new_n758), .ZN(new_n883));
  INV_X1    g697(.A(new_n749), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n759), .A2(new_n731), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n516), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n777), .A3(new_n778), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n886), .A2(new_n777), .A3(KEYINPUT121), .A4(new_n778), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n885), .A2(new_n699), .A3(new_n598), .A4(new_n516), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n892), .A2(new_n621), .A3(new_n620), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n883), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n875), .B(new_n877), .C1(new_n894), .C2(new_n876), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n622), .A3(new_n631), .ZN(new_n896));
  INV_X1    g710(.A(new_n767), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n889), .B2(new_n890), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT48), .ZN(new_n900));
  OAI211_X1 g714(.A(G952), .B(new_n345), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(KEYINPUT48), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n898), .A2(new_n900), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n872), .B(KEYINPUT120), .C1(new_n873), .C2(new_n874), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT51), .B1(new_n906), .B2(new_n894), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n868), .A2(new_n685), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n802), .B1(new_n866), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n302), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n706), .A2(new_n562), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n774), .A2(new_n598), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n879), .B(KEYINPUT49), .Z(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n700), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT112), .Z(new_n916));
  OAI21_X1  g730(.A(new_n801), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n838), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n848), .B1(new_n860), .B2(KEYINPUT53), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT54), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n865), .A2(new_n863), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n909), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n802), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n916), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(KEYINPUT123), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n917), .A2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n865), .A2(new_n188), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(G210), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n340), .A2(new_n349), .A3(new_n355), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n347), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n345), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  NAND2_X1  g751(.A1(new_n555), .A2(KEYINPUT57), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n555), .A2(KEYINPUT57), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n865), .A2(new_n863), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n859), .A2(new_n846), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(KEYINPUT53), .A3(new_n826), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n826), .B1(new_n831), .B2(new_n835), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT53), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n862), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n551), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n865), .A2(new_n188), .A3(new_n787), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n936), .B1(new_n949), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  INV_X1    g766(.A(new_n455), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n936), .ZN(G60));
  INV_X1    g770(.A(new_n936), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n618), .B(new_n960), .C1(new_n940), .C2(new_n947), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n866), .A2(new_n959), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n957), .B(new_n961), .C1(new_n962), .C2(new_n618), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(G63));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n965), .B1(new_n946), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g783(.A(KEYINPUT124), .B(new_n967), .C1(new_n942), .C2(new_n945), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n665), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT124), .B1(new_n865), .B2(new_n967), .ZN(new_n972));
  INV_X1    g786(.A(new_n595), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n946), .A2(new_n965), .A3(new_n968), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n971), .A2(new_n975), .A3(new_n957), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n971), .A2(new_n975), .A3(KEYINPUT61), .A4(new_n957), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G66));
  AOI21_X1  g794(.A(new_n345), .B1(new_n517), .B2(G224), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n851), .A2(new_n850), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n345), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n931), .B1(G898), .B2(new_n345), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  INV_X1    g801(.A(G900), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n539), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n269), .A2(new_n270), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n383), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n855), .A2(new_n858), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n708), .A3(new_n725), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n993), .A2(KEYINPUT62), .A3(new_n708), .A4(new_n725), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n727), .A2(new_n759), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n814), .A2(new_n805), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n999), .A2(new_n703), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n793), .A2(new_n799), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n998), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n992), .B1(new_n1004), .B2(new_n345), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n993), .A2(new_n725), .ZN(new_n1006));
  INV_X1    g820(.A(new_n742), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n792), .A2(new_n1007), .A3(new_n897), .ZN(new_n1008));
  INV_X1    g822(.A(new_n772), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1008), .A2(new_n770), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1003), .A2(new_n345), .A3(new_n1006), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G900), .A2(G953), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n992), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT127), .B(new_n989), .C1(new_n1005), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1001), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n1016), .B(new_n1002), .C1(new_n996), .C2(new_n997), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n991), .B1(new_n1017), .B2(G953), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1013), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1015), .A2(new_n1021), .ZN(G72));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1004), .B2(new_n982), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1025), .A2(new_n291), .A3(new_n264), .ZN(new_n1026));
  INV_X1    g840(.A(new_n292), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n861), .A2(new_n1027), .A3(new_n694), .A4(new_n1024), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1003), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1024), .B1(new_n1029), .B2(new_n982), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n936), .B1(new_n1030), .B2(new_n292), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1026), .A2(new_n1028), .A3(new_n1031), .ZN(G57));
endmodule


