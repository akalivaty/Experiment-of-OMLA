//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT80), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n196), .A2(new_n201), .A3(KEYINPUT4), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT64), .B1(new_n205), .B2(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n208), .B2(G143), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT65), .A3(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n204), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n216), .A2(KEYINPUT0), .A3(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT68), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(KEYINPUT0), .A3(G128), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n206), .A2(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n204), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n195), .A2(G101), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n203), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n194), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n189), .A2(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n198), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n208), .A2(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n205), .A2(G146), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(G128), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n216), .A2(KEYINPUT66), .A3(new_n233), .A4(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n216), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n230), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n243), .A2(KEYINPUT10), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n210), .A2(new_n214), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n240), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n198), .A4(new_n229), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n226), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G137), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(G137), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT11), .A3(G134), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n226), .A2(new_n258), .A3(new_n244), .A4(new_n248), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G140), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n264), .A2(G227), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n263), .B(new_n265), .Z(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT12), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT82), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n238), .A2(new_n246), .A3(new_n230), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n259), .B(new_n269), .C1(new_n270), .C2(new_n243), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n268), .A2(KEYINPUT82), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n238), .A2(new_n246), .A3(new_n230), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n236), .A2(new_n237), .B1(new_n241), .B2(new_n240), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n230), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n272), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n259), .A3(new_n277), .A4(new_n269), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n261), .A2(new_n266), .A3(new_n273), .A4(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n262), .A2(new_n267), .B1(new_n279), .B2(KEYINPUT84), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n281));
  AOI211_X1 g095(.A(new_n281), .B(new_n266), .C1(new_n260), .C2(new_n261), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n187), .B(new_n188), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n187), .A2(new_n188), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n261), .A2(new_n273), .A3(new_n278), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT83), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n261), .A2(new_n288), .A3(new_n273), .A4(new_n278), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n267), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n260), .A2(new_n261), .A3(new_n266), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n283), .B(new_n285), .C1(new_n187), .C2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  OAI21_X1  g108(.A(G221), .B1(new_n294), .B2(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G110), .B(G122), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n225), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT2), .B(G113), .Z(new_n302));
  XNOR2_X1  g116(.A(G116), .B(G119), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(KEYINPUT67), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(G116), .B(G119), .Z(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n301), .B(new_n309), .C1(new_n200), .C2(new_n202), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G116), .ZN(new_n313));
  OAI211_X1 g127(.A(G113), .B(new_n313), .C1(new_n305), .C2(new_n311), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n305), .B2(new_n306), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n315), .A2(new_n230), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n300), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n309), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n203), .A2(new_n319), .A3(new_n225), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n316), .A3(new_n299), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT85), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT86), .B1(new_n247), .B2(G125), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n220), .B1(new_n221), .B2(new_n204), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n238), .A2(new_n246), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n325), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G224), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G953), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  OAI221_X1 g148(.A(new_n300), .B1(KEYINPUT85), .B2(new_n322), .C1(new_n310), .C2(new_n317), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n299), .B(KEYINPUT8), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n315), .A2(new_n230), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n316), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n331), .B2(new_n333), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n325), .A2(new_n330), .ZN(new_n341));
  INV_X1    g155(.A(new_n333), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n342), .A4(new_n327), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT7), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n331), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(new_n343), .A3(new_n321), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n188), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G210), .B1(G237), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n336), .A2(new_n188), .A3(new_n348), .A4(new_n346), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n298), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n352), .A2(KEYINPUT87), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(KEYINPUT87), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n296), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n329), .A2(G140), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT16), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n358), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT16), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT74), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n361), .B(new_n364), .C1(KEYINPUT16), .C2(new_n357), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(new_n208), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n208), .ZN(new_n367));
  XNOR2_X1  g181(.A(G119), .B(G128), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT24), .B(G110), .Z(new_n369));
  AOI22_X1  g183(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n312), .A2(G128), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n371), .A2(KEYINPUT23), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(KEYINPUT23), .ZN(new_n373));
  INV_X1    g187(.A(G128), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n372), .B(new_n373), .C1(G119), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G110), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n359), .A2(new_n208), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n375), .A2(G110), .B1(new_n368), .B2(new_n369), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n366), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT75), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT22), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G137), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(G137), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n377), .A2(new_n380), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n380), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n376), .B2(new_n370), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n391));
  INV_X1    g205(.A(new_n385), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(new_n386), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(KEYINPUT76), .A3(new_n385), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n388), .B(new_n188), .C1(new_n390), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n377), .A2(new_n380), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n394), .A3(new_n393), .ZN(new_n400));
  INV_X1    g214(.A(new_n397), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n400), .A2(new_n188), .A3(new_n388), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G234), .ZN(new_n404));
  OAI21_X1  g218(.A(G217), .B1(new_n404), .B2(G902), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT73), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n400), .A2(new_n388), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(G902), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n403), .A2(new_n406), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT70), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G237), .ZN(new_n415));
  AOI21_X1  g229(.A(G953), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G210), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT27), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT26), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n420), .A3(G210), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n419), .B1(new_n418), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n197), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(G101), .A3(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n223), .A2(new_n259), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n256), .A2(G131), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n238), .B2(new_n246), .ZN(new_n432));
  INV_X1    g246(.A(new_n253), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n251), .A2(G137), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(new_n309), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT69), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n223), .A2(new_n259), .B1(new_n432), .B2(new_n435), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT69), .A3(new_n309), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n436), .B1(new_n258), .B2(new_n326), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n319), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT28), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT28), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n437), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n429), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n442), .B2(new_n429), .ZN(new_n454));
  AOI211_X1 g268(.A(KEYINPUT71), .B(new_n428), .C1(new_n439), .C2(new_n441), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n443), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n440), .A2(KEYINPUT30), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n319), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT31), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  AND4_X1   g276(.A1(KEYINPUT69), .A2(new_n430), .A3(new_n309), .A4(new_n436), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT69), .B1(new_n440), .B2(new_n309), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n429), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT71), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n442), .A2(new_n453), .A3(new_n429), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n466), .A2(KEYINPUT31), .A3(new_n461), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n452), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(G472), .A2(G902), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT32), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n461), .A3(new_n467), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT31), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n451), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  INV_X1    g291(.A(new_n471), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n461), .A2(new_n442), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n428), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n446), .A2(new_n450), .A3(new_n429), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n440), .A2(new_n309), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n439), .B2(new_n441), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n450), .B1(new_n486), .B2(new_n447), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n429), .A2(KEYINPUT29), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n188), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G472), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n472), .A2(new_n479), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n414), .A2(G237), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n412), .A2(KEYINPUT70), .ZN(new_n494));
  OAI211_X1 g308(.A(G214), .B(new_n264), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT88), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n416), .A2(KEYINPUT88), .A3(G214), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n205), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n416), .A2(G143), .A3(G214), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n498), .A4(new_n205), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G131), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n257), .A3(new_n502), .A4(new_n503), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n366), .A2(new_n367), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(KEYINPUT17), .A3(G131), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n189), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n504), .A2(KEYINPUT18), .A3(G131), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n362), .A2(G146), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n378), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(KEYINPUT18), .A2(G131), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n514), .B(new_n516), .C1(new_n517), .C2(new_n504), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n513), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n504), .A2(KEYINPUT18), .A3(G131), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n516), .B1(new_n504), .B2(new_n517), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n362), .B(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n366), .B1(G146), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n505), .B2(new_n507), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n520), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G475), .A2(G902), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n492), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT20), .B(new_n531), .C1(new_n519), .C2(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n511), .A2(new_n518), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n520), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n534), .B2(new_n519), .ZN(new_n535));
  INV_X1    g349(.A(G475), .ZN(new_n536));
  OAI22_X1  g350(.A1(new_n530), .A2(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G116), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G122), .ZN(new_n539));
  INV_X1    g353(.A(G122), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G116), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n541), .A3(new_n192), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT94), .Z(new_n543));
  OR2_X1    g357(.A1(new_n539), .A2(KEYINPUT14), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(KEYINPUT14), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G107), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n374), .B2(G143), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n205), .A2(KEYINPUT90), .A3(G128), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n205), .B2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n374), .A2(KEYINPUT92), .A3(G143), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n251), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n555), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G134), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n543), .B(new_n547), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n551), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n549), .B(new_n550), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(new_n566), .A3(new_n555), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G134), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n539), .A2(new_n541), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G107), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n542), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n556), .A2(new_n572), .A3(new_n251), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT93), .B1(new_n558), .B2(G134), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n571), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n294), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(G217), .A3(new_n264), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n560), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n560), .B2(new_n575), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n560), .A2(new_n575), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n580), .A3(new_n579), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n586), .A3(new_n188), .ZN(new_n587));
  INV_X1    g401(.A(G478), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT15), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n587), .B(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(G952), .A3(new_n264), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT21), .B(G898), .Z(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n537), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n355), .A2(new_n411), .A3(new_n491), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  OR2_X1    g415(.A1(new_n587), .A2(G478), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n579), .B1(new_n582), .B2(KEYINPUT97), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n560), .A2(new_n575), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n578), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n581), .A2(new_n582), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n604), .A2(new_n580), .A3(new_n578), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n602), .B1(new_n613), .B2(new_n588), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT98), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(new_n602), .C1(new_n613), .C2(new_n588), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n537), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n350), .A2(new_n351), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n297), .ZN(new_n621));
  AOI211_X1 g435(.A(KEYINPUT96), .B(new_n298), .C1(new_n350), .C2(new_n351), .ZN(new_n622));
  NOR4_X1   g436(.A1(new_n618), .A2(new_n621), .A3(new_n622), .A4(new_n598), .ZN(new_n623));
  INV_X1    g437(.A(new_n296), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n477), .B2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n470), .A2(new_n471), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n625), .A2(new_n626), .A3(new_n411), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n623), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n528), .A2(new_n529), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT20), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n531), .B1(new_n519), .B2(new_n527), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n492), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(KEYINPUT99), .A3(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n633), .A2(KEYINPUT99), .A3(new_n492), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n519), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n513), .B1(new_n511), .B2(new_n518), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n188), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n591), .B1(new_n640), .B2(G475), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n635), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  NOR4_X1   g456(.A1(new_n642), .A2(new_n621), .A3(new_n622), .A4(new_n598), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n624), .A3(new_n627), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT100), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT35), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n192), .ZN(G9));
  NAND2_X1  g461(.A1(new_n403), .A2(new_n406), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT36), .B1(new_n393), .B2(new_n394), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n399), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n410), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n625), .A2(new_n626), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT101), .A4(new_n652), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n599), .A3(new_n355), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AND2_X1   g475(.A1(new_n648), .A2(new_n651), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n296), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n621), .A2(new_n622), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n491), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n530), .A2(new_n532), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n636), .B1(new_n666), .B2(KEYINPUT99), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n594), .B(KEYINPUT104), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(G900), .B2(new_n596), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n667), .A2(new_n668), .A3(new_n641), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n635), .A2(new_n637), .A3(new_n641), .A4(new_n671), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT105), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n374), .ZN(G30));
  XNOR2_X1  g491(.A(new_n671), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n624), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT107), .Z(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n486), .A2(new_n429), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n456), .B2(new_n461), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n684), .B2(G902), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n472), .A2(new_n479), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n620), .B(KEYINPUT106), .Z(new_n687));
  INV_X1    g501(.A(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n537), .A2(new_n592), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n689), .A2(new_n297), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n682), .A2(new_n662), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  AND4_X1   g507(.A1(new_n537), .A2(new_n615), .A3(new_n617), .A4(new_n671), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n491), .A2(new_n663), .A3(new_n664), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  OAI21_X1  g510(.A(new_n188), .B1(new_n280), .B2(new_n282), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G469), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n295), .A3(new_n283), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n623), .A2(new_n411), .A3(new_n491), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n643), .A2(new_n411), .A3(new_n491), .A4(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NOR3_X1   g519(.A1(new_n621), .A2(new_n622), .A3(new_n699), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n491), .A3(new_n599), .A4(new_n652), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NAND2_X1  g522(.A1(new_n476), .A2(new_n468), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n487), .A2(new_n428), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n478), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n625), .A3(new_n411), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n621), .A2(new_n622), .A3(new_n598), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n690), .A4(new_n700), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NAND2_X1  g530(.A1(new_n470), .A2(new_n188), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n711), .B1(new_n717), .B2(G472), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n706), .A2(new_n718), .A3(new_n652), .A4(new_n694), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n290), .A2(KEYINPUT109), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n287), .A2(new_n723), .A3(new_n267), .A4(new_n289), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(G469), .A3(new_n291), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n283), .A3(new_n285), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n620), .A2(new_n298), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n726), .A2(new_n727), .A3(new_n295), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n491), .A2(new_n728), .A3(new_n411), .A4(new_n694), .ZN(new_n729));
  NOR2_X1   g543(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n721), .B(new_n731), .C1(new_n733), .C2(new_n730), .ZN(new_n734));
  INV_X1    g548(.A(new_n731), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT111), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n673), .A2(KEYINPUT105), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n673), .A2(KEYINPUT105), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n491), .A2(new_n411), .A3(new_n728), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n672), .A2(new_n674), .A3(KEYINPUT112), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  AND2_X1   g562(.A1(new_n615), .A2(new_n617), .ZN(new_n749));
  INV_X1    g563(.A(new_n666), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n640), .A2(G475), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT43), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n625), .A2(new_n626), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n652), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT114), .ZN(new_n758));
  INV_X1    g572(.A(new_n727), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n755), .B2(new_n756), .ZN(new_n760));
  INV_X1    g574(.A(new_n295), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n291), .A4(new_n724), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n292), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(G469), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n765), .B2(new_n285), .ZN(new_n766));
  INV_X1    g580(.A(new_n283), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n285), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n678), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n758), .A2(new_n760), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n774), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT47), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  INV_X1    g592(.A(new_n694), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n779), .A2(new_n491), .A3(new_n411), .A4(new_n759), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT116), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n777), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(new_n411), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n689), .A2(new_n784), .A3(new_n761), .ZN(new_n785));
  INV_X1    g599(.A(new_n686), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n698), .A2(new_n283), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT117), .Z(new_n789));
  AOI211_X1 g603(.A(new_n298), .B(new_n752), .C1(KEYINPUT49), .C2(new_n787), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n785), .A2(new_n786), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n734), .A2(new_n737), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n701), .A2(new_n704), .A3(new_n707), .A4(new_n715), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n618), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n750), .A2(new_n641), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n537), .A2(new_n615), .A3(KEYINPUT118), .A4(new_n617), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n597), .A3(new_n355), .A4(new_n627), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n657), .A3(new_n600), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n667), .A2(new_n671), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n727), .A2(new_n591), .A3(new_n751), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n491), .A3(new_n663), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n718), .A2(new_n728), .A3(new_n652), .A4(new_n694), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n794), .A2(new_n746), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n792), .B1(new_n793), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n719), .B(new_n695), .C1(new_n675), .C2(new_n665), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n686), .A2(new_n662), .A3(new_n671), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n726), .A2(new_n295), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n664), .A3(new_n690), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT120), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n491), .A2(new_n663), .A3(new_n664), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n672), .A2(new_n674), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n694), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n811), .A2(new_n664), .A3(new_n690), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n662), .A3(new_n671), .A4(new_n686), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n817), .A2(new_n818), .A3(new_n719), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n814), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n814), .B2(new_n821), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n746), .A2(new_n806), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n704), .A2(new_n701), .A3(new_n707), .A4(new_n715), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n800), .A2(new_n657), .A3(new_n600), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(KEYINPUT119), .A3(new_n738), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n808), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n829), .A2(KEYINPUT119), .A3(new_n738), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT119), .B1(new_n829), .B2(new_n738), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n814), .A2(new_n821), .A3(new_n822), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT52), .B1(new_n809), .B2(new_n813), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n832), .B(KEYINPUT54), .C1(new_n836), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n839), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n735), .B2(new_n736), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n807), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n831), .B2(new_n838), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n713), .A2(new_n700), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n664), .A2(new_n753), .A3(new_n669), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n689), .A2(new_n297), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n753), .A3(new_n669), .A4(new_n849), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(KEYINPUT50), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n852), .B2(new_n855), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n686), .A2(new_n594), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n759), .A2(new_n699), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n411), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n858), .A2(new_n537), .A3(new_n860), .A4(new_n749), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n856), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n777), .A2(new_n778), .B1(new_n295), .B2(new_n787), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n753), .A2(new_n669), .A3(new_n713), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n727), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n753), .A2(new_n669), .A3(new_n859), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n652), .A3(new_n718), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n858), .A2(new_n618), .A3(new_n860), .ZN(new_n873));
  INV_X1    g687(.A(G952), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(G953), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n491), .A2(new_n411), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n877), .B2(KEYINPUT48), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n866), .A2(KEYINPUT122), .A3(new_n876), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT48), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n848), .A2(new_n850), .A3(new_n871), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(G952), .A2(G953), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT123), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n791), .B1(new_n884), .B2(new_n886), .ZN(G75));
  NOR2_X1   g701(.A1(new_n845), .A2(new_n188), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(G210), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n324), .A2(new_n335), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n334), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  XOR2_X1   g706(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n893));
  AND3_X1   g707(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n264), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(G51));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n845), .B2(new_n846), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT53), .B1(new_n835), .B2(new_n825), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n901), .B2(new_n844), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n899), .B(KEYINPUT54), .C1(new_n901), .C2(new_n844), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n284), .B(KEYINPUT57), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n280), .A2(new_n282), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n845), .A2(new_n188), .A3(new_n765), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n897), .B1(new_n909), .B2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  INV_X1    g726(.A(new_n528), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n897), .ZN(G60));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n608), .A2(new_n612), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT126), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n904), .A2(new_n903), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n897), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n918), .B1(new_n841), .B2(new_n847), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n921), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n650), .B(new_n929), .C1(new_n901), .C2(new_n844), .ZN(new_n930));
  INV_X1    g744(.A(new_n407), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n845), .B2(new_n928), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n932), .A3(new_n923), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n933), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  AOI21_X1  g753(.A(new_n264), .B1(new_n595), .B2(G224), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n794), .A2(new_n801), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n264), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n890), .B1(G898), .B2(new_n264), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  INV_X1    g758(.A(new_n876), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n771), .A2(new_n945), .A3(new_n664), .A4(new_n690), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n772), .A2(new_n782), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n809), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n738), .A2(new_n746), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n264), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n460), .B(new_n524), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n950), .B(new_n952), .C1(G227), .C2(new_n264), .ZN(new_n953));
  OAI21_X1  g767(.A(G900), .B1(new_n952), .B2(G227), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n692), .A2(new_n948), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n692), .A2(KEYINPUT62), .A3(new_n948), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n945), .A2(new_n799), .ZN(new_n961));
  OR3_X1    g775(.A1(new_n680), .A2(new_n759), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n960), .A2(new_n782), .A3(new_n772), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n264), .A3(new_n951), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n953), .A2(new_n955), .A3(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n963), .B2(new_n941), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n429), .A3(new_n480), .ZN(new_n969));
  INV_X1    g783(.A(new_n480), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n947), .A2(new_n941), .A3(new_n949), .ZN(new_n971));
  INV_X1    g785(.A(new_n967), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n428), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n481), .B2(new_n474), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n832), .B(new_n974), .C1(new_n836), .C2(new_n840), .ZN(new_n975));
  AND4_X1   g789(.A1(new_n923), .A2(new_n969), .A3(new_n973), .A4(new_n975), .ZN(G57));
endmodule


