//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT66), .A2(G137), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT11), .A2(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT11), .B1(new_n189), .B2(G134), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  AOI21_X1  g010(.A(G131), .B1(new_n196), .B2(G137), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT66), .A2(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT66), .A2(G137), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n189), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n199), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT69), .B1(new_n198), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(G143), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n206), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT68), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT68), .A2(G128), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(G146), .ZN(new_n219));
  INV_X1    g033(.A(new_n210), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n226));
  INV_X1    g040(.A(new_n203), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n190), .A2(new_n191), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n196), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n225), .B(new_n226), .C1(new_n229), .C2(new_n199), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n205), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n196), .A2(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n193), .A2(new_n195), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT0), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(new_n221), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(KEYINPUT0), .B2(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n221), .A3(KEYINPUT64), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n210), .B1(new_n208), .B2(G146), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n209), .A2(new_n241), .B1(new_n242), .B2(new_n237), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(G116), .B(G119), .Z(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n231), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n231), .A2(new_n244), .A3(new_n251), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n231), .A2(new_n244), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n247), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n256), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n253), .A2(new_n255), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT74), .B(G902), .Z(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n198), .B2(new_n204), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n225), .B(KEYINPUT67), .C1(new_n229), .C2(new_n199), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n224), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n244), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n235), .B2(new_n243), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n248), .B1(new_n276), .B2(new_n231), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n249), .ZN(new_n279));
  INV_X1    g093(.A(new_n262), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT29), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n250), .A2(new_n252), .B1(new_n247), .B2(new_n273), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n262), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n268), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n187), .B1(new_n266), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n249), .A2(new_n262), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n278), .A2(new_n288), .A3(KEYINPUT31), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT31), .B1(new_n278), .B2(new_n288), .ZN(new_n290));
  OAI22_X1  g104(.A1(new_n289), .A2(new_n290), .B1(new_n282), .B2(new_n262), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n205), .A2(new_n224), .A3(new_n230), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n200), .A2(new_n201), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n194), .B1(new_n296), .B2(new_n192), .ZN(new_n297));
  AOI22_X1  g111(.A1(G131), .A2(new_n233), .B1(new_n297), .B2(new_n197), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n209), .A2(new_n241), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n219), .A2(new_n220), .A3(new_n237), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT30), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n247), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT30), .B1(new_n272), .B2(new_n244), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n249), .A2(new_n262), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n294), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n278), .A2(new_n288), .A3(KEYINPUT31), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n273), .A2(new_n247), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n253), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n280), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(KEYINPUT71), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n287), .B1(new_n293), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n285), .B1(new_n314), .B2(KEYINPUT32), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n314), .B2(KEYINPUT32), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n309), .A2(KEYINPUT71), .A3(new_n312), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT71), .B1(new_n309), .B2(new_n312), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n286), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT32), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n315), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(KEYINPUT68), .A2(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(KEYINPUT68), .A2(G128), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(KEYINPUT76), .A3(G119), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G119), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n212), .A2(new_n213), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n221), .B2(G119), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT16), .ZN(new_n338));
  INV_X1    g152(.A(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n340), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  INV_X1    g159(.A(G146), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(G146), .B(new_n340), .C1(new_n344), .C2(new_n338), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n327), .B2(G128), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT23), .B1(new_n221), .B2(G119), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n221), .A2(KEYINPUT79), .A3(G119), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n324), .A2(KEYINPUT23), .A3(G119), .A4(new_n325), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n212), .A2(new_n213), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n358), .A2(KEYINPUT78), .A3(KEYINPUT23), .A4(G119), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n354), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G110), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n349), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n331), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n360), .A2(new_n361), .B1(new_n363), .B2(new_n333), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n346), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n348), .A2(new_n366), .ZN(new_n367));
  OAI22_X1  g181(.A1(new_n337), .A2(new_n362), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT22), .B(G137), .ZN(new_n369));
  INV_X1    g183(.A(G221), .ZN(new_n370));
  INV_X1    g184(.A(G234), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n370), .A2(new_n371), .A3(G953), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n369), .B(new_n372), .Z(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  OAI221_X1 g189(.A(new_n349), .B1(new_n361), .B2(new_n360), .C1(new_n335), .C2(new_n336), .ZN(new_n376));
  AOI211_X1 g190(.A(G110), .B(new_n354), .C1(new_n357), .C2(new_n359), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n331), .A2(new_n334), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n366), .B(new_n348), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n379), .A3(new_n373), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n267), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n381), .A2(KEYINPUT25), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT25), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n375), .A2(new_n380), .A3(new_n383), .A4(new_n267), .ZN(new_n384));
  OAI21_X1  g198(.A(G217), .B1(new_n268), .B2(new_n371), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT75), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT80), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n375), .A2(new_n380), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n387), .A2(G902), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(KEYINPUT25), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n387), .A4(new_n384), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n389), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n323), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(KEYINPUT83), .A2(G107), .ZN(new_n401));
  NOR2_X1   g215(.A1(KEYINPUT83), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(G116), .B(G122), .Z(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n405), .A2(KEYINPUT14), .ZN(new_n407));
  INV_X1    g221(.A(G107), .ZN(new_n408));
  INV_X1    g222(.A(G122), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(G116), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n410), .B2(KEYINPUT14), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n358), .A2(G143), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n208), .A2(G128), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n417), .A2(new_n196), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT96), .ZN(new_n421));
  AOI21_X1  g235(.A(G134), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n412), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n196), .B1(new_n417), .B2(new_n418), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT97), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(KEYINPUT97), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n404), .B(new_n405), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT13), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n413), .B1(new_n414), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n414), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT95), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n414), .A2(new_n434), .A3(new_n430), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n429), .B1(new_n436), .B2(new_n196), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n423), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT9), .B(G234), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(G217), .A3(new_n258), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n436), .A2(new_n196), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(new_n426), .A3(new_n429), .A4(new_n427), .ZN(new_n444));
  INV_X1    g258(.A(new_n441), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n423), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n400), .B1(new_n447), .B2(new_n267), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n268), .B(new_n399), .C1(new_n442), .C2(new_n446), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n257), .A2(new_n258), .A3(G214), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n452), .A2(new_n206), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n208), .A2(new_n452), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(G131), .ZN(new_n456));
  AND2_X1   g270(.A1(KEYINPUT94), .A2(KEYINPUT19), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n344), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n344), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n346), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n348), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(KEYINPUT18), .A2(G131), .ZN(new_n463));
  OR3_X1    g277(.A1(new_n455), .A2(KEYINPUT93), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n344), .A2(G146), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n366), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n463), .B1(new_n455), .B2(KEYINPUT93), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G113), .B(G122), .ZN(new_n470));
  INV_X1    g284(.A(G104), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n456), .A2(KEYINPUT17), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n455), .A2(KEYINPUT17), .A3(G131), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n347), .A3(new_n348), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n472), .B(new_n468), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G475), .A2(G902), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n451), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n480), .ZN(new_n482));
  AOI211_X1 g296(.A(KEYINPUT20), .B(new_n482), .C1(new_n474), .C2(new_n478), .ZN(new_n483));
  INV_X1    g297(.A(G475), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n468), .B1(new_n475), .B2(new_n477), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n473), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n481), .A2(new_n483), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n258), .A2(G952), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(G234), .B2(G237), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n258), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G898), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n450), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n397), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G214), .B1(G237), .B2(G902), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT86), .Z(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT91), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  OR2_X1    g317(.A1(KEYINPUT82), .A2(G104), .ZN(new_n504));
  NAND2_X1  g318(.A1(KEYINPUT82), .A2(G104), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(G107), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n507));
  OR2_X1    g321(.A1(KEYINPUT83), .A2(G107), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT83), .A2(G107), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n506), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G101), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n515), .A2(new_n247), .ZN(new_n516));
  AND2_X1   g330(.A1(KEYINPUT82), .A2(G104), .ZN(new_n517));
  NOR2_X1   g331(.A1(KEYINPUT82), .A2(G104), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n408), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n519), .A2(KEYINPUT3), .B1(new_n403), .B2(new_n507), .ZN(new_n520));
  INV_X1    g334(.A(G101), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n506), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n514), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n513), .A2(G101), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT84), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n516), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G113), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n327), .A2(G116), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n245), .B2(new_n529), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n245), .A2(new_n246), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(G104), .B1(new_n508), .B2(new_n509), .ZN(new_n535));
  OAI21_X1  g349(.A(G101), .B1(new_n511), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n506), .A2(new_n521), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n527), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G110), .B(G122), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n503), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT84), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT4), .B1(new_n537), .B2(new_n538), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n521), .B1(new_n520), .B2(new_n506), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n524), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n540), .B1(new_n551), .B2(new_n516), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT88), .B1(new_n552), .B2(new_n543), .ZN(new_n553));
  AND4_X1   g367(.A1(KEYINPUT88), .A2(new_n527), .A3(new_n541), .A4(new_n543), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n545), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n542), .A2(new_n503), .A3(new_n544), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n224), .A2(new_n342), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n342), .B2(new_n301), .ZN(new_n558));
  INV_X1    g372(.A(G224), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G953), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT89), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n558), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n555), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n542), .B2(new_n544), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n543), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n543), .B(KEYINPUT8), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n519), .B1(new_n403), .B2(G104), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n520), .A2(new_n522), .B1(new_n569), .B2(G101), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n534), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT5), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n531), .B1(new_n572), .B2(new_n245), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n539), .B1(new_n533), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n558), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT7), .A3(new_n561), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n561), .A2(KEYINPUT7), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n558), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n567), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n502), .B1(new_n563), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI211_X1 g399(.A(KEYINPUT92), .B(new_n502), .C1(new_n563), .C2(new_n582), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n563), .A2(new_n582), .A3(new_n502), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n499), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G902), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n370), .B1(new_n440), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n590), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n242), .B1(G128), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n570), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n539), .A2(new_n215), .A3(new_n223), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n235), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT85), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n515), .A2(new_n243), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n549), .B2(new_n550), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n215), .B2(new_n223), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n570), .ZN(new_n608));
  INV_X1    g422(.A(new_n242), .ZN(new_n609));
  AOI21_X1  g423(.A(G146), .B1(new_n216), .B2(new_n218), .ZN(new_n610));
  OAI21_X1  g424(.A(G128), .B1(new_n610), .B2(new_n211), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n594), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n539), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n608), .B1(new_n613), .B2(KEYINPUT10), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n603), .B1(new_n615), .B2(new_n298), .ZN(new_n616));
  INV_X1    g430(.A(new_n604), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n525), .B2(new_n526), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n597), .A2(new_n606), .B1(new_n570), .B2(new_n607), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n603), .A4(new_n298), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n602), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(G110), .B(G140), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT81), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n258), .A2(G227), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n618), .A2(new_n619), .A3(new_n298), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT85), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n629), .B2(new_n620), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n235), .B1(new_n605), .B2(new_n614), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n622), .A2(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n593), .B1(new_n632), .B2(G469), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n620), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n634), .A2(new_n626), .A3(new_n602), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n626), .B1(new_n634), .B2(new_n631), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n592), .B(new_n267), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n591), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n589), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n497), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n521), .ZN(G3));
  AOI21_X1  g455(.A(new_n268), .B1(new_n293), .B2(new_n313), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n319), .B1(new_n642), .B2(new_n187), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n644), .A2(new_n638), .A3(new_n396), .ZN(new_n645));
  INV_X1    g459(.A(new_n499), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n563), .A2(new_n582), .A3(new_n502), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(new_n583), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n268), .A2(new_n398), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n447), .A2(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n447), .A2(KEYINPUT33), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(G478), .B1(new_n447), .B2(new_n267), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n488), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n648), .A2(new_n655), .A3(new_n494), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n645), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  NOR4_X1   g473(.A1(new_n648), .A2(new_n450), .A3(new_n488), .A4(new_n494), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n374), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n368), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n391), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n389), .A2(new_n395), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n389), .A2(KEYINPUT98), .A3(new_n395), .A4(new_n666), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n496), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n589), .A2(new_n638), .A3(new_n644), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR2_X1   g489(.A1(new_n648), .A2(new_n671), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n491), .B1(new_n492), .B2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n450), .A2(new_n488), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n676), .A2(new_n323), .A3(new_n638), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  NAND2_X1  g495(.A1(new_n587), .A2(new_n588), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n678), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n638), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n255), .A2(new_n249), .A3(new_n280), .ZN(new_n690));
  INV_X1    g504(.A(new_n249), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n275), .B2(new_n277), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n692), .B2(new_n280), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n693), .B2(KEYINPUT100), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n187), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n314), .B2(KEYINPUT32), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n316), .A2(new_n697), .A3(new_n322), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n488), .B1(new_n448), .B2(new_n449), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n699), .A2(new_n667), .A3(new_n499), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n684), .A2(new_n688), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n208), .ZN(G45));
  INV_X1    g517(.A(new_n652), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n447), .A2(KEYINPUT33), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n649), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n654), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n678), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n488), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n676), .A2(new_n323), .A3(new_n638), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NOR2_X1   g527(.A1(new_n635), .A2(new_n636), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(new_n268), .ZN(new_n715));
  INV_X1    g529(.A(new_n591), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n637), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n656), .A2(new_n323), .A3(new_n396), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n660), .A2(new_n323), .A3(new_n396), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NOR2_X1   g537(.A1(new_n717), .A2(new_n648), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n323), .A3(new_n672), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n323), .A3(new_n672), .A4(KEYINPUT102), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NAND2_X1  g544(.A1(new_n563), .A2(new_n582), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n501), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n499), .B(new_n699), .C1(new_n732), .C2(new_n588), .ZN(new_n733));
  INV_X1    g547(.A(new_n309), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n262), .B1(new_n253), .B2(new_n255), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n286), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n396), .B(new_n736), .C1(new_n642), .C2(new_n187), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n718), .A2(new_n733), .A3(new_n738), .A4(new_n495), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  OAI211_X1 g554(.A(new_n667), .B(new_n736), .C1(new_n642), .C2(new_n187), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n710), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n588), .A2(new_n646), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n585), .A2(new_n586), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n323), .A2(new_n747), .A3(new_n638), .A4(new_n396), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n748), .B2(new_n710), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(KEYINPUT103), .B(new_n745), .C1(new_n748), .C2(new_n710), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n315), .B1(KEYINPUT32), .B2(new_n314), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n754), .A2(KEYINPUT104), .A3(new_n396), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT104), .B1(new_n754), .B2(new_n396), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n747), .A2(new_n638), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n711), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  XOR2_X1   g576(.A(new_n679), .B(KEYINPUT105), .Z(new_n763));
  OR2_X1    g577(.A1(new_n748), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n622), .A2(new_n627), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n630), .A2(new_n631), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n592), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n632), .A2(KEYINPUT45), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n593), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n593), .B1(new_n770), .B2(new_n771), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n637), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n716), .B(new_n686), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n488), .B1(new_n706), .B2(new_n707), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(KEYINPUT107), .B2(KEYINPUT43), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n667), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n783), .B1(new_n788), .B2(new_n644), .ZN(new_n789));
  INV_X1    g603(.A(new_n747), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n644), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(KEYINPUT44), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n781), .A2(new_n782), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  OAI21_X1  g608(.A(new_n716), .B1(new_n776), .B2(new_n778), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n797), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  OR4_X1    g615(.A1(new_n323), .A2(new_n790), .A3(new_n396), .A4(new_n710), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n798), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND3_X1  g618(.A1(new_n784), .A2(new_n646), .A3(new_n716), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n715), .A2(new_n637), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n806), .B(new_n396), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n807), .B2(new_n809), .ZN(new_n811));
  INV_X1    g625(.A(new_n698), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n684), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n718), .A2(new_n747), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n491), .A2(new_n815), .A3(new_n396), .A4(new_n812), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n489), .A3(new_n707), .A4(new_n706), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n815), .A2(new_n491), .A3(new_n787), .ZN(new_n818));
  INV_X1    g632(.A(new_n741), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n787), .A2(new_n491), .A3(new_n738), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n646), .A3(new_n717), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n684), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n823), .A2(KEYINPUT50), .A3(new_n684), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(KEYINPUT118), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(KEYINPUT118), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n821), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n809), .A2(new_n591), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n798), .B2(new_n801), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n822), .A2(new_n790), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n818), .B1(new_n756), .B2(new_n755), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT48), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n490), .B(KEYINPUT119), .Z(new_n842));
  INV_X1    g656(.A(new_n724), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n822), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n655), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n844), .B1(new_n816), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT120), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n847), .A2(KEYINPUT120), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n839), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n680), .A2(new_n712), .A3(new_n743), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n389), .A2(new_n395), .A3(new_n666), .A4(new_n709), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n591), .B(new_n855), .C1(new_n633), .C2(new_n637), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n698), .A2(new_n856), .A3(new_n733), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n698), .A2(new_n856), .A3(new_n733), .A4(KEYINPUT111), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n853), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n854), .B1(new_n853), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n852), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n680), .A2(new_n712), .A3(new_n743), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT52), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n719), .A2(new_n739), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n729), .A2(new_n722), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n760), .B2(new_n753), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n448), .ZN(new_n874));
  INV_X1    g688(.A(new_n449), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT109), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT109), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n448), .B2(new_n449), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n488), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n845), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n494), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n589), .A3(new_n645), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n673), .C1(new_n497), .C2(new_n639), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n488), .A2(new_n678), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n876), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n638), .A2(new_n885), .A3(new_n669), .A4(new_n670), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(KEYINPUT110), .A3(new_n323), .A4(new_n747), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n323), .A2(new_n747), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n758), .A2(new_n742), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n764), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n883), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(KEYINPUT53), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n871), .A2(new_n872), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n868), .A2(new_n873), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT112), .B1(new_n865), .B2(new_n866), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n853), .A2(new_n854), .A3(new_n861), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT52), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n864), .A2(new_n871), .A3(new_n901), .A4(new_n895), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n902), .A2(KEYINPUT114), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT114), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n851), .B(new_n898), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n871), .A2(new_n895), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n868), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n902), .A2(new_n903), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT54), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n835), .B(KEYINPUT116), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n798), .B2(new_n801), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n837), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT51), .B1(new_n834), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n850), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n813), .B1(new_n916), .B2(new_n917), .ZN(G75));
  OAI21_X1  g732(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n501), .A3(new_n268), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n555), .A2(new_n556), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n562), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT55), .Z(new_n924));
  AND3_X1   g738(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n920), .B2(new_n921), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n258), .A2(G952), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n593), .B(KEYINPUT57), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n902), .A2(new_n903), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT114), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n902), .A2(KEYINPUT114), .A3(new_n903), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n851), .B1(new_n934), .B2(new_n898), .ZN(new_n935));
  INV_X1    g749(.A(new_n906), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n714), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n919), .A2(new_n268), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(new_n772), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n927), .B1(new_n939), .B2(new_n941), .ZN(G54));
  NAND2_X1  g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n479), .ZN(new_n945));
  INV_X1    g759(.A(new_n927), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n478), .B(new_n474), .C1(new_n940), .C2(new_n943), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G60));
  NAND2_X1  g762(.A1(G478), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT59), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n911), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n704), .A2(new_n705), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n952), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n950), .C1(new_n935), .C2(new_n936), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n953), .A2(new_n946), .A3(new_n955), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT121), .Z(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n919), .A2(new_n665), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n959), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n934), .B2(new_n898), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n960), .B(new_n946), .C1(new_n962), .C2(new_n390), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n919), .A2(new_n959), .ZN(new_n966));
  INV_X1    g780(.A(new_n390), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n927), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n960), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n969), .ZN(G66));
  NOR2_X1   g784(.A1(new_n870), .A2(new_n883), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(G953), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n493), .B2(new_n559), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(G898), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n922), .B1(new_n976), .B2(G953), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n975), .B(new_n977), .Z(G69));
  AND2_X1   g792(.A1(new_n793), .A2(new_n803), .ZN(new_n979));
  NOR4_X1   g793(.A1(new_n397), .A2(new_n790), .A3(new_n880), .A4(new_n687), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  OR3_X1    g795(.A1(new_n702), .A2(new_n981), .A3(new_n866), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n702), .B2(new_n866), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(G953), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n304), .B1(new_n231), .B2(new_n276), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(new_n460), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n986), .B1(new_n985), .B2(new_n988), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n258), .B1(G227), .B2(G900), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n989), .A2(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n757), .A2(new_n648), .A3(new_n699), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n781), .A2(new_n782), .A3(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n761), .A2(new_n764), .A3(new_n853), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n979), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n979), .A2(new_n996), .A3(new_n999), .A4(new_n995), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n258), .A2(G900), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n988), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n992), .A2(new_n991), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n993), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1005), .B1(new_n993), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1006), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  NAND2_X1  g824(.A1(new_n979), .A2(new_n984), .ZN(new_n1011));
  INV_X1    g825(.A(new_n971), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1015), .B(new_n1010), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1014), .A2(new_n262), .A3(new_n279), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n908), .A2(new_n909), .ZN(new_n1018));
  OAI22_X1  g832(.A1(new_n692), .A2(new_n262), .B1(new_n305), .B2(new_n306), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n1010), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1017), .B(new_n946), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n278), .A2(new_n249), .A3(new_n280), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n998), .A2(new_n1000), .A3(new_n971), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1023), .B2(new_n1010), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1021), .A2(new_n1024), .ZN(G57));
endmodule


