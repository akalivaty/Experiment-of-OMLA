//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n458), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n463), .A2(G136), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT66), .Z(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT67), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(new_n475), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT68), .Z(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n459), .A2(new_n461), .A3(G126), .A4(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n459), .A2(new_n461), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n486), .A2(new_n487), .A3(G138), .A4(new_n475), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n459), .A2(new_n461), .A3(G138), .A4(new_n475), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n488), .B2(new_n490), .ZN(G164));
  XNOR2_X1  g066(.A(KEYINPUT6), .B(G651), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G543), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G50), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT69), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n499), .A2(G88), .B1(new_n507), .B2(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n496), .A2(new_n508), .ZN(G166));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n510));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  INV_X1    g088(.A(G89), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n498), .ZN(new_n515));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n503), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT70), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n502), .A2(new_n504), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n492), .A2(G51), .A3(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT71), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n516), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n502), .A2(new_n504), .A3(new_n520), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n520), .B1(new_n502), .B2(new_n504), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n492), .A2(G51), .A3(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n515), .B1(new_n524), .B2(new_n531), .ZN(G168));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n498), .A2(new_n533), .B1(new_n493), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n519), .A2(new_n521), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n539), .B2(G651), .ZN(G171));
  XOR2_X1   g115(.A(KEYINPUT74), .B(G81), .Z(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n498), .A2(new_n541), .B1(new_n493), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  OAI21_X1  g120(.A(G56), .B1(new_n526), .B2(new_n527), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n519), .B2(new_n521), .ZN(new_n552));
  INV_X1    g127(.A(new_n547), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n492), .A2(G53), .A3(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n492), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n505), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n499), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(new_n535), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n536), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n545), .ZN(G301));
  INV_X1    g151(.A(new_n515), .ZN(new_n577));
  NOR3_X1   g152(.A1(new_n522), .A2(KEYINPUT71), .A3(new_n523), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(G286));
  NAND2_X1  g155(.A1(new_n496), .A2(new_n508), .ZN(G303));
  NAND2_X1  g156(.A1(new_n494), .A2(G49), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n582), .A2(new_n583), .B1(G87), .B2(new_n499), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n494), .A2(KEYINPUT75), .A3(G49), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  INV_X1    g163(.A(G73), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT76), .B1(new_n589), .B2(new_n501), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(G73), .A3(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n590), .B(new_n592), .C1(new_n505), .C2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(G86), .A2(new_n499), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n492), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n545), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n498), .A2(new_n602), .B1(new_n493), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n499), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n498), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n505), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(G54), .A2(new_n494), .B1(new_n615), .B2(G651), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(G868), .B2(new_n617), .ZN(G284));
  OAI21_X1  g193(.A(new_n607), .B1(G868), .B2(new_n617), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G299), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G168), .B2(new_n620), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(G168), .B2(new_n620), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n612), .A2(new_n616), .ZN(new_n626));
  OAI21_X1  g201(.A(G868), .B1(new_n626), .B2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n556), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n486), .A2(new_n464), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n478), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n463), .A2(G135), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(G2100), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT16), .B(G1341), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(G14), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n647), .A2(new_n653), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT17), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT78), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n660), .B2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2096), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT79), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n672), .A3(new_n673), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT81), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n672), .A2(new_n673), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n682), .A2(new_n674), .A3(new_n676), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT82), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n693), .A3(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G29), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G162), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT29), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G2090), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n617), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G4), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT87), .B(G1348), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G26), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n478), .A2(G128), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n463), .A2(G140), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(new_n707), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G2067), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n704), .B2(new_n705), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n702), .A2(G20), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT23), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G299), .B2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n721), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(G1956), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n706), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G1956), .B2(new_n724), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n702), .A2(G19), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n556), .B2(new_n702), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1341), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n701), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G168), .A2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT93), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G21), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n638), .A2(new_n707), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT94), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G160), .B2(new_n707), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G2084), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(G29), .A2(G32), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G105), .B2(new_n464), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n478), .A2(G129), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n463), .A2(G141), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(new_n707), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT31), .B(G11), .Z(new_n757));
  INV_X1    g332(.A(G28), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT30), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n758), .B2(KEYINPUT30), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n707), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n707), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n746), .A2(new_n756), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G171), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1961), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n737), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G33), .ZN(new_n771));
  NAND2_X1  g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  INV_X1    g347(.A(G127), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n462), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT89), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n464), .A2(G103), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n463), .A2(G139), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n771), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G2072), .Z(new_n786));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n744), .A2(G2084), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT91), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n754), .B2(new_n755), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n787), .B1(new_n786), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n770), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(new_n770), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n732), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G23), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n586), .A2(new_n587), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n702), .A2(G6), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n595), .A2(new_n598), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n702), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT84), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n702), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n702), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(G1971), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(G1971), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n809), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n798), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n803), .A2(new_n814), .A3(new_n798), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n702), .A2(G24), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n605), .B2(new_n702), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n707), .A2(G25), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G119), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n463), .A2(G131), .ZN(new_n824));
  OR2_X1    g399(.A1(G95), .A2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n822), .B1(new_n828), .B2(new_n707), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  NOR2_X1   g406(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n818), .A2(KEYINPUT85), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT85), .B1(new_n818), .B2(new_n832), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n815), .B(new_n817), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n815), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n836), .A2(new_n816), .A3(KEYINPUT36), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n797), .B1(new_n835), .B2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n835), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n839), .A2(new_n794), .A3(new_n796), .A4(new_n732), .ZN(G150));
  AOI22_X1  g415(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n492), .A2(new_n497), .A3(G93), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n492), .A2(G55), .A3(G543), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT96), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT96), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n841), .A2(new_n545), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NOR2_X1   g423(.A1(new_n626), .A2(new_n624), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n536), .A2(G67), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n845), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT96), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n854), .A2(G651), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n550), .B2(new_n555), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n543), .B1(new_n554), .B2(KEYINPUT73), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n548), .A2(new_n549), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n846), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n851), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n851), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n848), .B1(new_n863), .B2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n753), .B(new_n715), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G164), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n784), .ZN(new_n869));
  INV_X1    g444(.A(new_n782), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n463), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n475), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G130), .B2(new_n478), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n631), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n827), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n470), .B(new_n638), .ZN(new_n882));
  XNOR2_X1  g457(.A(G162), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n871), .A2(new_n878), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n880), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n879), .A2(new_n883), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g466(.A1(G290), .A2(new_n587), .A3(new_n586), .ZN(new_n892));
  NAND2_X1  g467(.A1(G288), .A2(new_n605), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(G305), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT98), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT42), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n626), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G299), .B1(new_n612), .B2(new_n616), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n617), .A2(G299), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n626), .A2(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n626), .A2(G559), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n862), .B(new_n912), .ZN(new_n913));
  MUX2_X1   g488(.A(new_n910), .B(new_n911), .S(new_n913), .Z(new_n914));
  OR2_X1    g489(.A1(new_n901), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n620), .B1(new_n901), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n915), .A2(new_n916), .B1(new_n620), .B2(new_n846), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(new_n918), .ZN(G295));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n918), .ZN(G331));
  AND3_X1   g497(.A1(new_n859), .A2(new_n860), .A3(new_n846), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n924));
  NOR2_X1   g499(.A1(G286), .A2(G171), .ZN(new_n925));
  NOR2_X1   g500(.A1(G168), .A2(G301), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G286), .A2(G171), .ZN(new_n928));
  NAND2_X1  g503(.A1(G168), .A2(G301), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n858), .A2(new_n928), .A3(new_n861), .A4(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n911), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT103), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n927), .A2(new_n933), .A3(new_n930), .A4(new_n911), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n935));
  AOI221_X4 g510(.A(new_n935), .B1(new_n906), .B2(new_n909), .C1(new_n927), .C2(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n927), .A2(new_n930), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT102), .B1(new_n937), .B2(new_n910), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n932), .B(new_n934), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n899), .A2(new_n898), .ZN(new_n940));
  INV_X1    g515(.A(new_n897), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n910), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n935), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n937), .A2(KEYINPUT102), .A3(new_n910), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n932), .A2(new_n934), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n900), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n939), .A2(new_n942), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n943), .A2(new_n944), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT101), .B(KEYINPUT43), .Z(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n949), .A3(new_n900), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(KEYINPUT104), .ZN(new_n957));
  INV_X1    g532(.A(new_n954), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n945), .A2(new_n931), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n942), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n957), .A2(new_n958), .A3(new_n951), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n943), .A2(new_n944), .A3(new_n951), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT105), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n953), .A2(new_n954), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n966), .A2(KEYINPUT105), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G397));
  AND3_X1   g546(.A1(new_n465), .A2(G40), .A3(new_n469), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(G164), .B2(G1384), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(G290), .A2(G1986), .ZN(new_n977));
  NAND2_X1  g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n753), .B(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G2067), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n715), .B(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n828), .A2(new_n830), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n828), .A2(new_n830), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n981), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n976), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT114), .B(G1956), .Z(new_n988));
  NOR2_X1   g563(.A1(G164), .A2(G1384), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n972), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n975), .A2(new_n972), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT56), .B(G2072), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n903), .A2(KEYINPUT115), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n999), .A2(KEYINPUT115), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(KEYINPUT115), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G299), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n994), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n994), .B2(new_n998), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT119), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT61), .ZN(new_n1008));
  NOR2_X1   g583(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n996), .A2(new_n980), .A3(new_n972), .A4(new_n975), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n989), .A2(new_n972), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT58), .B(G1341), .Z(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1014), .B2(new_n556), .ZN(new_n1015));
  NAND2_X1  g590(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT118), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1017), .ZN(new_n1019));
  AOI211_X1 g594(.A(new_n1009), .B(new_n1019), .C1(new_n1014), .C2(new_n556), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT61), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT119), .B(new_n1022), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1008), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT120), .ZN(new_n1025));
  OR3_X1    g600(.A1(new_n1011), .A2(KEYINPUT116), .A3(G2067), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n1011), .B2(G2067), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n488), .A2(new_n490), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n485), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n972), .A3(new_n991), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1026), .B(new_n1027), .C1(new_n1033), .C2(G1348), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1034), .A2(KEYINPUT60), .A3(new_n626), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1034), .B(new_n617), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(KEYINPUT60), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1008), .A2(new_n1021), .A3(new_n1038), .A4(new_n1023), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1025), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1034), .A2(new_n617), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1005), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1006), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1030), .A2(new_n974), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n975), .A2(new_n972), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1050), .A2(G1971), .B1(new_n1032), .B2(G2090), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1047), .A2(new_n1051), .A3(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1047), .B1(G8), .B2(new_n1051), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n586), .A2(G1976), .A3(new_n587), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT106), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1011), .B2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  AOI211_X1 g633(.A(KEYINPUT106), .B(new_n1058), .C1(new_n989), .C2(new_n972), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(KEYINPUT107), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1055), .B(new_n1062), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1065));
  NOR2_X1   g640(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G288), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n805), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G305), .A2(G1981), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT49), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1057), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1011), .A2(new_n1056), .A3(G8), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1073), .A2(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT110), .B1(new_n1068), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1060), .A2(new_n1063), .B1(G288), .B2(new_n1066), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1082), .B2(new_n1065), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT110), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1054), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n995), .A2(new_n764), .A3(new_n996), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1050), .A2(KEYINPUT53), .A3(new_n764), .ZN(new_n1090));
  INV_X1    g665(.A(G1961), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1032), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1086), .B1(new_n1093), .B2(G171), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1087), .A2(new_n1088), .B1(new_n1032), .B2(new_n1091), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(G301), .A3(new_n1090), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1096), .B2(new_n1090), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1094), .A2(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(new_n1086), .A3(KEYINPUT54), .A4(new_n1097), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n736), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT111), .B(G2084), .Z(new_n1106));
  NAND4_X1  g681(.A1(new_n1031), .A2(new_n972), .A3(new_n991), .A4(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g684(.A(G168), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1058), .B1(KEYINPUT122), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(KEYINPUT122), .B2(new_n1111), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT51), .B1(new_n1116), .B2(G8), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(G286), .B(new_n1114), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G168), .A2(new_n1058), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1115), .A2(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1085), .A2(new_n1103), .A3(KEYINPUT124), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1117), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1100), .B(new_n1102), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1068), .A2(KEYINPUT110), .A3(new_n1079), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1080), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1124), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1044), .A2(new_n1123), .A3(new_n1131), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1058), .B(G286), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT112), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1128), .B(new_n1134), .C1(new_n1129), .C2(new_n1080), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1128), .A2(new_n1134), .A3(KEYINPUT63), .A4(new_n1083), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1052), .A2(new_n1053), .A3(new_n1136), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1141), .A2(KEYINPUT113), .A3(new_n1083), .A4(new_n1134), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1128), .B(new_n1099), .C1(new_n1129), .C2(new_n1080), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT125), .B1(new_n1121), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(KEYINPUT62), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1121), .A2(new_n1146), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1083), .A2(new_n1052), .ZN(new_n1152));
  OR2_X1    g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1070), .B1(new_n1078), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT108), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT109), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1143), .A2(new_n1151), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n987), .B1(new_n1132), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT46), .ZN(new_n1163));
  INV_X1    g738(.A(new_n976), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(G1996), .ZN(new_n1165));
  INV_X1    g740(.A(new_n983), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n976), .B1(new_n1166), .B2(new_n753), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n976), .A2(KEYINPUT46), .A3(new_n980), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT47), .Z(new_n1170));
  NOR2_X1   g745(.A1(new_n977), .A2(new_n1164), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT126), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(KEYINPUT48), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1172), .A2(KEYINPUT48), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1173), .B(new_n1174), .C1(new_n976), .C2(new_n986), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n981), .A2(new_n983), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1176), .A2(new_n985), .B1(G2067), .B2(new_n715), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1170), .B(new_n1175), .C1(new_n976), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1162), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g754(.A(G319), .B1(new_n654), .B2(new_n655), .ZN(new_n1181));
  NOR2_X1   g755(.A1(G227), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n695), .A2(new_n696), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n1183), .B1(new_n887), .B2(new_n889), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n962), .A2(new_n1184), .ZN(G225));
  NAND2_X1  g759(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1186));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n1187), .A3(new_n1184), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1188), .ZN(G308));
endmodule


