//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n541, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  INV_X1    g037(.A(G101), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n458), .A2(G2104), .ZN(new_n464));
  OAI22_X1  g039(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n459), .A2(new_n460), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OR3_X1    g042(.A1(new_n466), .A2(KEYINPUT65), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT65), .B1(new_n466), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n471), .B2(G2105), .ZN(G160));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n458), .ZN(new_n473));
  MUX2_X1   g048(.A(G100), .B(G112), .S(G2105), .Z(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G124), .B1(G2104), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT66), .Z(G162));
  INV_X1    g053(.A(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G138), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G114), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(G126), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n466), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT4), .A2(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n466), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n458), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n482), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  XNOR2_X1  g067(.A(KEYINPUT5), .B(G543), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n493), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n495), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n502), .A2(new_n503), .A3(new_n493), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n502), .B2(new_n493), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT69), .B(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n502), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n496), .B1(new_n512), .B2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n516));
  AND3_X1   g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n493), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n502), .A2(G543), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(G89), .B2(new_n506), .ZN(G168));
  NAND2_X1  g098(.A1(new_n506), .A2(G90), .ZN(new_n524));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT5), .B(G543), .Z(new_n526));
  INV_X1    g101(.A(G64), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n510), .A2(G52), .B1(new_n528), .B2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  NAND2_X1  g106(.A1(new_n506), .A2(G81), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(G43), .ZN(new_n533));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G56), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n510), .A2(new_n533), .B1(new_n536), .B2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G188));
  INV_X1    g120(.A(new_n497), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n495), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT67), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n493), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT68), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n502), .A2(new_n503), .A3(new_n493), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(G91), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n553), .B(new_n554), .C1(new_n521), .C2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n493), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n495), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n552), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n510), .A2(KEYINPUT73), .A3(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n553), .B1(new_n521), .B2(new_n555), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n506), .A2(G89), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n510), .A2(G51), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n564), .A2(new_n565), .A3(new_n519), .A4(new_n518), .ZN(G286));
  NAND2_X1  g141(.A1(new_n506), .A2(G87), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n493), .A2(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n510), .A2(G49), .B1(G651), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n526), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n510), .A2(G48), .B1(new_n573), .B2(G651), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n550), .A2(new_n551), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n493), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n495), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n506), .A2(G85), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n510), .A2(G47), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G301), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n550), .A2(G92), .A3(new_n551), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n550), .A2(KEYINPUT10), .A3(G92), .A4(new_n551), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n521), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n502), .A2(KEYINPUT75), .A3(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n526), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n594), .A2(G54), .B1(G651), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n585), .B1(new_n600), .B2(new_n584), .ZN(G284));
  AOI21_X1  g176(.A(new_n585), .B1(new_n600), .B2(new_n584), .ZN(G321));
  MUX2_X1   g177(.A(G286), .B(G299), .S(new_n584), .Z(G297));
  MUX2_X1   g178(.A(G286), .B(G299), .S(new_n584), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n600), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n605), .A3(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n539), .A2(new_n584), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT11), .Z(G282));
  INV_X1    g185(.A(new_n609), .ZN(G323));
  NAND2_X1  g186(.A1(new_n479), .A2(G2104), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n613), .B(new_n615), .ZN(new_n616));
  MUX2_X1   g191(.A(G99), .B(G111), .S(G2105), .Z(new_n617));
  AOI22_X1  g192(.A1(new_n473), .A2(G123), .B1(G2104), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G135), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n461), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT15), .B(G2435), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2427), .ZN(new_n627));
  INV_X1    g202(.A(G2430), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT77), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n630), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT78), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT79), .Z(G401));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT17), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2084), .B(G2090), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n646), .B2(new_n644), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT80), .Z(new_n652));
  INV_X1    g227(.A(new_n649), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n653), .A2(new_n646), .A3(new_n644), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n646), .A2(new_n649), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n655), .B1(new_n645), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n621), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G229));
  NOR2_X1   g252(.A1(G16), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT84), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n685), .B2(G22), .ZN(new_n686));
  AND3_X1   g261(.A1(new_n685), .A2(KEYINPUT85), .A3(G22), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n686), .B(new_n687), .C1(G303), .C2(G16), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G6), .A2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G305), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT32), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n688), .A2(new_n689), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n684), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n684), .A2(new_n696), .A3(new_n697), .A4(new_n699), .ZN(new_n702));
  OR2_X1    g277(.A1(G16), .A2(G24), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G290), .B2(new_n685), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT81), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n473), .A2(G119), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n479), .A2(G131), .ZN(new_n712));
  MUX2_X1   g287(.A(G95), .B(G107), .S(G2105), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2104), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(new_n708), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AND4_X1   g294(.A1(KEYINPUT86), .A2(new_n706), .A3(new_n707), .A4(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n701), .A2(new_n702), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT29), .Z(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT97), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT24), .A2(G34), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(G29), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G160), .B2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2084), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n727), .B2(new_n728), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n708), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  MUX2_X1   g314(.A(G104), .B(G116), .S(G2105), .Z(new_n740));
  AOI22_X1  g315(.A1(new_n473), .A2(G128), .B1(G2104), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G140), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n461), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT87), .Z(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n744), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(G2067), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n708), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n473), .A2(G129), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT93), .Z(new_n750));
  XOR2_X1   g325(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n479), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  INV_X1    g330(.A(new_n464), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G105), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n748), .B1(new_n759), .B2(new_n708), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n685), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n685), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G27), .A2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G164), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n762), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n737), .A2(new_n747), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G4), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n600), .B2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G1348), .Z(new_n775));
  NOR2_X1   g350(.A1(new_n734), .A2(G2084), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G19), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n539), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1341), .ZN(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G127), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n466), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n458), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n479), .A2(KEYINPUT88), .A3(G139), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n788));
  INV_X1    g363(.A(G139), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n461), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT25), .ZN(new_n791));
  INV_X1    g366(.A(G103), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n464), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n756), .A2(KEYINPUT25), .A3(G103), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n787), .A2(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT90), .Z(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  AOI211_X1 g373(.A(new_n777), .B(new_n780), .C1(new_n798), .C2(G2072), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n730), .A2(new_n772), .A3(new_n775), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(G2072), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT91), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n685), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  INV_X1    g379(.A(G299), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n685), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1956), .Z(new_n807));
  NOR2_X1   g382(.A1(new_n764), .A2(new_n765), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT31), .B(G11), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT30), .B(G28), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n708), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n620), .B2(new_n708), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n685), .A2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G168), .B2(new_n685), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1966), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n808), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n802), .A2(new_n807), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n800), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n723), .A2(new_n724), .A3(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  NAND2_X1  g398(.A1(new_n600), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n493), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(new_n495), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT98), .B(G93), .Z(new_n828));
  NAND3_X1  g403(.A1(new_n550), .A2(new_n551), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n510), .A2(G55), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n829), .A2(KEYINPUT99), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT99), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n538), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n539), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n825), .B(new_n839), .Z(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n834), .A2(new_n836), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n849), .ZN(G145));
  MUX2_X1   g425(.A(G106), .B(G118), .S(G2105), .Z(new_n851));
  AOI22_X1  g426(.A1(new_n473), .A2(G130), .B1(G2104), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n461), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n613), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n715), .B(KEYINPUT103), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n797), .B(new_n759), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n744), .B(G164), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  OAI211_X1 g437(.A(KEYINPUT104), .B(new_n857), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n864), .A2(new_n860), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(G162), .B(G160), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n620), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n868), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(G395));
  NOR2_X1   g450(.A1(new_n846), .A2(G868), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n679), .B(G290), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  NAND2_X1  g453(.A1(G303), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(KEYINPUT107), .B(new_n496), .C1(new_n512), .C2(new_n513), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(G305), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G305), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n877), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n600), .A2(new_n605), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n839), .B(new_n890), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n599), .A2(G299), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n590), .A2(new_n559), .A3(new_n598), .A4(new_n562), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n839), .B(new_n890), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n900), .A3(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT41), .B1(new_n893), .B2(new_n895), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI211_X1 g480(.A(KEYINPUT106), .B(new_n900), .C1(new_n892), .C2(new_n894), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  AND4_X1   g484(.A1(new_n889), .A2(new_n897), .A3(new_n898), .A4(new_n909), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n889), .A2(new_n898), .B1(new_n897), .B2(new_n909), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n910), .A2(new_n911), .B1(KEYINPUT108), .B2(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n897), .A2(new_n909), .ZN(new_n913));
  INV_X1    g488(.A(new_n898), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n888), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n889), .A2(new_n897), .A3(new_n898), .A4(new_n909), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n876), .B1(new_n919), .B2(G868), .ZN(G295));
  AOI21_X1  g495(.A(new_n876), .B1(new_n919), .B2(G868), .ZN(G331));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND3_X1  g497(.A1(G286), .A2(KEYINPUT110), .A3(G301), .ZN(new_n923));
  NAND2_X1  g498(.A1(G301), .A2(KEYINPUT110), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(G168), .B1(G301), .B2(KEYINPUT110), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n837), .A2(new_n838), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n837), .B2(new_n838), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n904), .B2(new_n901), .ZN(new_n931));
  INV_X1    g506(.A(new_n927), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n839), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n837), .A2(new_n838), .A3(new_n927), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n896), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n889), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n930), .A2(KEYINPUT112), .A3(new_n896), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n906), .B1(new_n904), .B2(new_n903), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n930), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n934), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT111), .B1(new_n944), .B2(new_n908), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n939), .B(new_n940), .C1(new_n943), .C2(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n922), .B(new_n937), .C1(new_n946), .C2(new_n889), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n889), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n941), .B1(new_n930), .B2(new_n942), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(new_n908), .A3(KEYINPUT111), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(new_n888), .A3(new_n939), .A4(new_n940), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n949), .A2(new_n950), .A3(new_n922), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n947), .A2(new_n950), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n922), .A4(new_n954), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(G397));
  XNOR2_X1  g536(.A(new_n744), .B(new_n746), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n759), .B(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G160), .A2(G40), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n480), .A2(new_n481), .B1(new_n489), .B2(new_n458), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n966), .B2(new_n486), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT114), .Z(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n715), .B(new_n718), .Z(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(G290), .A2(G1986), .ZN(new_n977));
  AND2_X1   g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT115), .Z(new_n980));
  AND2_X1   g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT124), .ZN(new_n982));
  AND2_X1   g557(.A1(G160), .A2(G40), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n967), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT119), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n967), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n491), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(KEYINPUT119), .A3(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1348), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n965), .A2(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n746), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n982), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n986), .B1(new_n990), .B2(new_n993), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT124), .B(new_n997), .C1(new_n1000), .C2(G1348), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n599), .B1(new_n1002), .B2(KEYINPUT60), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT60), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1004), .B(new_n600), .C1(new_n999), .C2(new_n1001), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n1003), .A2(new_n1005), .B1(KEYINPUT60), .B2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT61), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n984), .B1(new_n491), .B2(new_n991), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1008), .A2(new_n965), .A3(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(G1956), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G299), .B(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n969), .B1(new_n491), .B2(new_n991), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n965), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n967), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT117), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1013), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1013), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1007), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1022), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n1020), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT58), .B(G1341), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1026), .A2(G1996), .B1(new_n996), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT126), .A3(new_n539), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT59), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1028), .A2(KEYINPUT126), .A3(new_n1031), .A4(new_n539), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1023), .A2(new_n1025), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT125), .B1(new_n1002), .B2(new_n599), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT125), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n999), .A2(new_n1001), .A3(new_n1036), .A4(new_n600), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1024), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1006), .A2(new_n1034), .B1(new_n1038), .B2(new_n1020), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1015), .B(new_n769), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1000), .A2(G1961), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT127), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT127), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1046), .A3(new_n1042), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(G301), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n983), .B(KEYINPUT122), .C1(KEYINPUT45), .C2(new_n967), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(new_n965), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n967), .A2(new_n969), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1055), .A2(new_n1042), .A3(G2078), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1000), .A2(G1961), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1040), .B1(new_n1049), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  XNOR2_X1  g637(.A(G305), .B(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(KEYINPUT49), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n965), .B2(new_n992), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n692), .A2(new_n1062), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G305), .A2(G1981), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1065), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n679), .B2(G1976), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n1076));
  INV_X1    g651(.A(G1976), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G288), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1066), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1067), .A2(new_n1074), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1072), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G303), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1026), .A2(new_n689), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n987), .A2(new_n728), .A3(new_n994), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(G8), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1026), .A2(new_n689), .B1(new_n1010), .B2(new_n728), .ZN(new_n1093));
  INV_X1    g668(.A(G8), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1086), .B(new_n1087), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1083), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1055), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G2084), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1000), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1100), .A3(G168), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT51), .ZN(new_n1103));
  AOI21_X1  g678(.A(G168), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  OAI211_X1 g680(.A(G8), .B(new_n1101), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1096), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1058), .A2(G301), .A3(new_n1059), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(KEYINPUT54), .C1(G301), .C2(new_n1048), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1061), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1039), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1060), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n1096), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT62), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1103), .A2(new_n1106), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G288), .A2(G1976), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1070), .B1(new_n1072), .B2(new_n1119), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1092), .A2(new_n1082), .B1(new_n1120), .B2(new_n1066), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(G8), .A3(G168), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1091), .A2(G8), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1125), .A2(new_n1092), .A3(new_n1083), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1124), .B1(new_n1096), .B2(new_n1123), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1121), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1118), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n981), .B1(new_n1111), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G1996), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n971), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT46), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(KEYINPUT46), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n962), .A2(new_n759), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1135), .A2(new_n1136), .B1(new_n1137), .B2(new_n971), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT47), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n971), .A2(new_n977), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT48), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n976), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n716), .A2(new_n718), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n974), .A2(new_n1143), .B1(G2067), .B2(new_n744), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1144), .A2(new_n971), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1139), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1132), .A2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g722(.A(new_n642), .ZN(new_n1149));
  INV_X1    g723(.A(G319), .ZN(new_n1150));
  NOR4_X1   g724(.A1(new_n1149), .A2(new_n1150), .A3(G227), .A4(G229), .ZN(new_n1151));
  NAND4_X1  g725(.A1(new_n957), .A2(new_n1151), .A3(new_n873), .A4(new_n958), .ZN(G225));
  INV_X1    g726(.A(G225), .ZN(G308));
endmodule


