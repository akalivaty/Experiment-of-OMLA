

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  NOR2_X1 U381 ( .A1(n615), .A2(n711), .ZN(n617) );
  XNOR2_X1 U382 ( .A(n399), .B(n398), .ZN(n740) );
  XNOR2_X1 U383 ( .A(n384), .B(n358), .ZN(n531) );
  INV_X1 U384 ( .A(KEYINPUT64), .ZN(n411) );
  NOR2_X1 U385 ( .A1(n682), .A2(n537), .ZN(n540) );
  INV_X2 U386 ( .A(G146), .ZN(n431) );
  OR2_X1 U387 ( .A1(n578), .A2(n572), .ZN(n580) );
  XNOR2_X2 U388 ( .A(n410), .B(n409), .ZN(n495) );
  NOR2_X2 U389 ( .A1(G902), .A2(n709), .ZN(n454) );
  XNOR2_X2 U390 ( .A(n431), .B(G125), .ZN(n468) );
  XNOR2_X2 U391 ( .A(n499), .B(n421), .ZN(n727) );
  XNOR2_X2 U392 ( .A(n467), .B(G134), .ZN(n499) );
  XOR2_X2 U393 ( .A(G122), .B(G104), .Z(n484) );
  NOR2_X2 U394 ( .A1(n532), .A2(n506), .ZN(n412) );
  INV_X1 U395 ( .A(KEYINPUT48), .ZN(n419) );
  AND2_X1 U396 ( .A1(n371), .A2(n362), .ZN(n592) );
  XNOR2_X1 U397 ( .A(n372), .B(n419), .ZN(n371) );
  AND2_X1 U398 ( .A1(n553), .A2(n692), .ZN(n374) );
  OR2_X1 U399 ( .A1(n578), .A2(n400), .ZN(n399) );
  XNOR2_X1 U400 ( .A(n543), .B(n542), .ZN(n560) );
  NOR2_X1 U401 ( .A1(n460), .A2(G902), .ZN(n462) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n493) );
  XNOR2_X2 U403 ( .A(KEYINPUT101), .B(n519), .ZN(n650) );
  XNOR2_X2 U404 ( .A(n479), .B(n478), .ZN(n712) );
  XNOR2_X2 U405 ( .A(n420), .B(KEYINPUT39), .ZN(n517) );
  XNOR2_X2 U406 ( .A(n388), .B(KEYINPUT96), .ZN(n573) );
  XNOR2_X2 U407 ( .A(n462), .B(n461), .ZN(n388) );
  AND2_X1 U408 ( .A1(n397), .A2(n395), .ZN(n579) );
  INV_X1 U409 ( .A(n740), .ZN(n397) );
  NOR2_X1 U410 ( .A1(n509), .A2(n630), .ZN(n521) );
  XNOR2_X1 U411 ( .A(n504), .B(G469), .ZN(n523) );
  XNOR2_X1 U412 ( .A(n394), .B(n364), .ZN(n415) );
  NAND2_X1 U413 ( .A1(n560), .A2(n559), .ZN(n394) );
  AND2_X1 U414 ( .A1(n380), .A2(n378), .ZN(n377) );
  NOR2_X1 U415 ( .A1(n379), .A2(KEYINPUT79), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n393), .B(n425), .ZN(n392) );
  NAND2_X1 U417 ( .A1(n493), .A2(G210), .ZN(n393) );
  XNOR2_X1 U418 ( .A(n426), .B(n390), .ZN(n389) );
  XNOR2_X1 U419 ( .A(n391), .B(KEYINPUT73), .ZN(n390) );
  INV_X1 U420 ( .A(KEYINPUT90), .ZN(n391) );
  XNOR2_X1 U421 ( .A(G113), .B(KEYINPUT3), .ZN(n423) );
  XNOR2_X1 U422 ( .A(n417), .B(n416), .ZN(n403) );
  XOR2_X1 U423 ( .A(G116), .B(G107), .Z(n498) );
  XNOR2_X1 U424 ( .A(n448), .B(n430), .ZN(n433) );
  XNOR2_X1 U425 ( .A(G131), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X1 U426 ( .A(KEYINPUT33), .B(n563), .ZN(n655) );
  AND2_X1 U427 ( .A1(n581), .A2(n584), .ZN(n563) );
  OR2_X1 U428 ( .A1(n698), .A2(G902), .ZN(n384) );
  INV_X1 U429 ( .A(G472), .ZN(n461) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT12), .ZN(n485) );
  XOR2_X1 U431 ( .A(KEYINPUT93), .B(G143), .Z(n492) );
  NOR2_X1 U432 ( .A1(n655), .A2(n570), .ZN(n564) );
  XNOR2_X1 U433 ( .A(n523), .B(n505), .ZN(n628) );
  NAND2_X1 U434 ( .A1(n415), .A2(n414), .ZN(n571) );
  NOR2_X1 U435 ( .A1(n648), .A2(n630), .ZN(n414) );
  BUF_X1 U436 ( .A(n388), .Z(n369) );
  XNOR2_X1 U437 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U438 ( .A(KEYINPUT25), .ZN(n451) );
  AND2_X2 U439 ( .A1(n407), .A2(n406), .ZN(n707) );
  AND2_X1 U440 ( .A1(n595), .A2(n622), .ZN(n406) );
  NAND2_X1 U441 ( .A1(n404), .A2(n408), .ZN(n407) );
  INV_X1 U442 ( .A(KEYINPUT2), .ZN(n408) );
  NOR2_X1 U443 ( .A1(n729), .A2(G952), .ZN(n711) );
  XNOR2_X1 U444 ( .A(n518), .B(KEYINPUT40), .ZN(n741) );
  NAND2_X1 U445 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U446 ( .A1(n376), .A2(n375), .ZN(n546) );
  XNOR2_X1 U447 ( .A(n425), .B(G140), .ZN(n448) );
  INV_X1 U448 ( .A(KEYINPUT81), .ZN(n554) );
  XOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT92), .Z(n486) );
  XNOR2_X1 U450 ( .A(n467), .B(n468), .ZN(n470) );
  XOR2_X1 U451 ( .A(KEYINPUT17), .B(KEYINPUT75), .Z(n472) );
  XNOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n471) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n456) );
  XNOR2_X1 U454 ( .A(n392), .B(n389), .ZN(n427) );
  XNOR2_X1 U455 ( .A(n591), .B(KEYINPUT66), .ZN(n401) );
  INV_X1 U456 ( .A(KEYINPUT8), .ZN(n409) );
  XNOR2_X1 U457 ( .A(G119), .B(G128), .ZN(n442) );
  XOR2_X1 U458 ( .A(G122), .B(KEYINPUT94), .Z(n497) );
  XNOR2_X1 U459 ( .A(n365), .B(n359), .ZN(n604) );
  XNOR2_X1 U460 ( .A(n434), .B(n727), .ZN(n365) );
  XOR2_X1 U461 ( .A(G110), .B(G101), .Z(n436) );
  INV_X1 U462 ( .A(G953), .ZN(n716) );
  AND2_X1 U463 ( .A1(n368), .A2(n367), .ZN(n544) );
  INV_X1 U464 ( .A(n523), .ZN(n367) );
  XNOR2_X1 U465 ( .A(n522), .B(KEYINPUT28), .ZN(n368) );
  XNOR2_X1 U466 ( .A(n385), .B(n361), .ZN(n698) );
  XNOR2_X1 U467 ( .A(n489), .B(n490), .ZN(n385) );
  NOR2_X1 U468 ( .A1(n527), .A2(n535), .ZN(n528) );
  XNOR2_X1 U469 ( .A(n568), .B(KEYINPUT35), .ZN(n739) );
  INV_X1 U470 ( .A(KEYINPUT32), .ZN(n398) );
  NAND2_X1 U471 ( .A1(n396), .A2(n575), .ZN(n395) );
  XNOR2_X1 U472 ( .A(n580), .B(KEYINPUT97), .ZN(n396) );
  NAND2_X1 U473 ( .A1(n360), .A2(n386), .ZN(n586) );
  XNOR2_X1 U474 ( .A(n613), .B(n614), .ZN(n615) );
  XOR2_X1 U475 ( .A(KEYINPUT13), .B(G475), .Z(n358) );
  XOR2_X1 U476 ( .A(n436), .B(n435), .Z(n359) );
  AND2_X1 U477 ( .A1(n455), .A2(n562), .ZN(n360) );
  XOR2_X1 U478 ( .A(n494), .B(n422), .Z(n361) );
  INV_X1 U479 ( .A(G104), .ZN(n430) );
  INV_X1 U480 ( .A(G137), .ZN(n425) );
  AND2_X1 U481 ( .A1(n695), .A2(n697), .ZN(n362) );
  NAND2_X1 U482 ( .A1(n588), .A2(KEYINPUT71), .ZN(n363) );
  XOR2_X1 U483 ( .A(n561), .B(KEYINPUT0), .Z(n364) );
  NAND2_X1 U484 ( .A1(n495), .A2(G217), .ZN(n496) );
  OR2_X2 U485 ( .A1(n704), .A2(G902), .ZN(n413) );
  XNOR2_X1 U486 ( .A(n449), .B(n726), .ZN(n709) );
  XNOR2_X1 U487 ( .A(n490), .B(n448), .ZN(n726) );
  NAND2_X1 U488 ( .A1(n513), .A2(n644), .ZN(n527) );
  NAND2_X1 U489 ( .A1(n521), .A2(n557), .ZN(n510) );
  NAND2_X1 U490 ( .A1(n403), .A2(n590), .ZN(n402) );
  NAND2_X1 U491 ( .A1(n418), .A2(n366), .ZN(n417) );
  INV_X1 U492 ( .A(n739), .ZN(n366) );
  NAND2_X1 U493 ( .A1(n373), .A2(n374), .ZN(n372) );
  XNOR2_X1 U494 ( .A(n712), .B(n480), .ZN(n610) );
  XNOR2_X2 U495 ( .A(n524), .B(KEYINPUT42), .ZN(n737) );
  NAND2_X1 U496 ( .A1(n645), .A2(n644), .ZN(n519) );
  XNOR2_X2 U497 ( .A(n535), .B(KEYINPUT38), .ZN(n645) );
  XNOR2_X2 U498 ( .A(n370), .B(KEYINPUT41), .ZN(n642) );
  NAND2_X1 U499 ( .A1(n650), .A2(n569), .ZN(n370) );
  XNOR2_X1 U500 ( .A(n526), .B(n525), .ZN(n373) );
  INV_X1 U501 ( .A(n683), .ZN(n375) );
  NAND2_X1 U502 ( .A1(n377), .A2(n363), .ZN(n376) );
  AND2_X1 U503 ( .A1(n545), .A2(KEYINPUT71), .ZN(n379) );
  NOR2_X1 U504 ( .A1(n545), .A2(KEYINPUT71), .ZN(n381) );
  INV_X1 U505 ( .A(n588), .ZN(n382) );
  INV_X1 U506 ( .A(KEYINPUT79), .ZN(n383) );
  INV_X1 U507 ( .A(n369), .ZN(n386) );
  XNOR2_X1 U508 ( .A(n388), .B(n387), .ZN(n581) );
  INV_X1 U509 ( .A(KEYINPUT6), .ZN(n387) );
  NOR2_X1 U510 ( .A1(n634), .A2(n369), .ZN(n635) );
  NAND2_X1 U511 ( .A1(n584), .A2(n369), .ZN(n638) );
  INV_X2 U512 ( .A(n541), .ZN(n535) );
  XNOR2_X2 U513 ( .A(n592), .B(n554), .ZN(n618) );
  NAND2_X1 U514 ( .A1(n729), .A2(G234), .ZN(n410) );
  XNOR2_X2 U515 ( .A(n411), .B(G953), .ZN(n729) );
  INV_X1 U516 ( .A(n415), .ZN(n570) );
  INV_X1 U517 ( .A(n395), .ZN(n678) );
  OR2_X1 U518 ( .A1(n577), .A2(n628), .ZN(n400) );
  XNOR2_X2 U519 ( .A(n402), .B(n401), .ZN(n717) );
  NAND2_X1 U520 ( .A1(n405), .A2(n717), .ZN(n404) );
  XNOR2_X1 U521 ( .A(n618), .B(KEYINPUT74), .ZN(n405) );
  XNOR2_X2 U522 ( .A(n412), .B(n507), .ZN(n686) );
  XNOR2_X2 U523 ( .A(n413), .B(G478), .ZN(n532) );
  XNOR2_X2 U524 ( .A(G143), .B(G128), .ZN(n467) );
  INV_X1 U525 ( .A(KEYINPUT44), .ZN(n416) );
  XNOR2_X1 U526 ( .A(n579), .B(KEYINPUT86), .ZN(n418) );
  NAND2_X1 U527 ( .A1(n517), .A2(n686), .ZN(n518) );
  NAND2_X1 U528 ( .A1(n530), .A2(n645), .ZN(n420) );
  NOR2_X2 U529 ( .A1(n465), .A2(n466), .ZN(n530) );
  INV_X1 U530 ( .A(n477), .ZN(n478) );
  AND2_X1 U531 ( .A1(G214), .A2(n493), .ZN(n422) );
  XNOR2_X1 U532 ( .A(n431), .B(G107), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n480) );
  INV_X1 U535 ( .A(G469), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U537 ( .A(KEYINPUT63), .ZN(n599) );
  XNOR2_X1 U538 ( .A(n669), .B(n668), .ZN(G75) );
  XNOR2_X1 U539 ( .A(n727), .B(G146), .ZN(n429) );
  XOR2_X1 U540 ( .A(G101), .B(G119), .Z(n424) );
  XNOR2_X1 U541 ( .A(n424), .B(n423), .ZN(n477) );
  XNOR2_X1 U542 ( .A(G116), .B(KEYINPUT5), .ZN(n426) );
  XNOR2_X1 U543 ( .A(n477), .B(n427), .ZN(n428) );
  XNOR2_X1 U544 ( .A(n429), .B(n428), .ZN(n460) );
  XNOR2_X1 U545 ( .A(n460), .B(KEYINPUT62), .ZN(n597) );
  NAND2_X1 U546 ( .A1(G227), .A2(n729), .ZN(n435) );
  NOR2_X1 U547 ( .A1(G902), .A2(n604), .ZN(n504) );
  XNOR2_X1 U548 ( .A(n504), .B(n437), .ZN(n455) );
  XOR2_X1 U549 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n440) );
  XOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .Z(n595) );
  INV_X1 U551 ( .A(n595), .ZN(n438) );
  NAND2_X1 U552 ( .A1(G234), .A2(n438), .ZN(n439) );
  XNOR2_X1 U553 ( .A(n440), .B(n439), .ZN(n450) );
  NAND2_X1 U554 ( .A1(n450), .A2(G221), .ZN(n441) );
  XNOR2_X1 U555 ( .A(n441), .B(KEYINPUT21), .ZN(n630) );
  NAND2_X1 U556 ( .A1(G221), .A2(n495), .ZN(n447) );
  XOR2_X1 U557 ( .A(KEYINPUT88), .B(G110), .Z(n443) );
  XOR2_X1 U558 ( .A(n443), .B(n442), .Z(n445) );
  XOR2_X1 U559 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n444) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U561 ( .A(KEYINPUT10), .B(n468), .Z(n490) );
  NAND2_X1 U562 ( .A1(n450), .A2(G217), .ZN(n452) );
  XNOR2_X2 U563 ( .A(n454), .B(n453), .ZN(n631) );
  NOR2_X1 U564 ( .A1(n630), .A2(n631), .ZN(n562) );
  XOR2_X1 U565 ( .A(KEYINPUT14), .B(n456), .Z(n661) );
  INV_X1 U566 ( .A(n661), .ZN(n557) );
  NOR2_X1 U567 ( .A1(n729), .A2(G900), .ZN(n457) );
  NAND2_X1 U568 ( .A1(G902), .A2(n457), .ZN(n458) );
  NAND2_X1 U569 ( .A1(G952), .A2(n716), .ZN(n555) );
  NAND2_X1 U570 ( .A1(n458), .A2(n555), .ZN(n508) );
  AND2_X1 U571 ( .A1(n557), .A2(n508), .ZN(n459) );
  NAND2_X1 U572 ( .A1(n360), .A2(n459), .ZN(n466) );
  NOR2_X1 U573 ( .A1(G237), .A2(G902), .ZN(n463) );
  XOR2_X1 U574 ( .A(KEYINPUT72), .B(n463), .Z(n481) );
  NAND2_X1 U575 ( .A1(n481), .A2(G214), .ZN(n644) );
  NAND2_X1 U576 ( .A1(n573), .A2(n644), .ZN(n464) );
  XNOR2_X1 U577 ( .A(n464), .B(KEYINPUT30), .ZN(n465) );
  NAND2_X1 U578 ( .A1(G224), .A2(n729), .ZN(n469) );
  XNOR2_X1 U579 ( .A(n470), .B(n469), .ZN(n474) );
  XNOR2_X1 U580 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U581 ( .A(G110), .B(KEYINPUT16), .Z(n475) );
  XNOR2_X1 U582 ( .A(n484), .B(n475), .ZN(n476) );
  XNOR2_X1 U583 ( .A(n476), .B(n498), .ZN(n479) );
  NOR2_X1 U584 ( .A1(n595), .A2(n610), .ZN(n483) );
  NAND2_X1 U585 ( .A1(G210), .A2(n481), .ZN(n482) );
  XNOR2_X1 U586 ( .A(n483), .B(n482), .ZN(n541) );
  XNOR2_X1 U587 ( .A(n484), .B(KEYINPUT91), .ZN(n488) );
  XNOR2_X1 U588 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U589 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U590 ( .A(G113), .B(G131), .ZN(n491) );
  XNOR2_X1 U591 ( .A(n492), .B(n491), .ZN(n494) );
  INV_X1 U592 ( .A(n531), .ZN(n506) );
  XNOR2_X1 U593 ( .A(n497), .B(n496), .ZN(n503) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n501) );
  XNOR2_X1 U595 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U596 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U597 ( .A(n503), .B(n502), .Z(n704) );
  NAND2_X1 U598 ( .A1(n506), .A2(n532), .ZN(n679) );
  INV_X1 U599 ( .A(n679), .ZN(n688) );
  NAND2_X1 U600 ( .A1(n517), .A2(n688), .ZN(n695) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(KEYINPUT67), .Z(n505) );
  INV_X1 U602 ( .A(n628), .ZN(n572) );
  INV_X1 U603 ( .A(KEYINPUT95), .ZN(n507) );
  INV_X1 U604 ( .A(n581), .ZN(n576) );
  NAND2_X1 U605 ( .A1(n631), .A2(n508), .ZN(n509) );
  NOR2_X1 U606 ( .A1(n576), .A2(n510), .ZN(n511) );
  NAND2_X1 U607 ( .A1(n686), .A2(n511), .ZN(n512) );
  XNOR2_X1 U608 ( .A(n512), .B(KEYINPUT99), .ZN(n513) );
  NOR2_X1 U609 ( .A1(n572), .A2(n527), .ZN(n515) );
  XOR2_X1 U610 ( .A(KEYINPUT43), .B(KEYINPUT100), .Z(n514) );
  XNOR2_X1 U611 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U612 ( .A1(n535), .A2(n516), .ZN(n697) );
  NOR2_X1 U613 ( .A1(n532), .A2(n531), .ZN(n569) );
  AND2_X1 U614 ( .A1(n573), .A2(n557), .ZN(n520) );
  AND2_X1 U615 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U616 ( .A1(n642), .A2(n544), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n741), .A2(n737), .ZN(n526) );
  XNOR2_X1 U618 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n528), .B(KEYINPUT36), .ZN(n529) );
  NAND2_X1 U620 ( .A1(n529), .A2(n572), .ZN(n692) );
  NAND2_X1 U621 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U622 ( .A(KEYINPUT98), .B(n533), .Z(n565) );
  NAND2_X1 U623 ( .A1(n530), .A2(n565), .ZN(n534) );
  NOR2_X1 U624 ( .A1(n535), .A2(n534), .ZN(n682) );
  NOR2_X2 U625 ( .A1(n688), .A2(n686), .ZN(n588) );
  INV_X1 U626 ( .A(KEYINPUT47), .ZN(n538) );
  NOR2_X1 U627 ( .A1(n382), .A2(n538), .ZN(n536) );
  NOR2_X1 U628 ( .A1(KEYINPUT80), .A2(n536), .ZN(n537) );
  NAND2_X1 U629 ( .A1(KEYINPUT79), .A2(n538), .ZN(n539) );
  NAND2_X1 U630 ( .A1(n540), .A2(n539), .ZN(n547) );
  NAND2_X1 U631 ( .A1(n541), .A2(n644), .ZN(n543) );
  XNOR2_X1 U632 ( .A(KEYINPUT19), .B(KEYINPUT68), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n544), .A2(n560), .ZN(n683) );
  XNOR2_X1 U634 ( .A(KEYINPUT70), .B(KEYINPUT47), .ZN(n545) );
  NOR2_X1 U635 ( .A1(n547), .A2(n546), .ZN(n552) );
  NAND2_X1 U636 ( .A1(n588), .A2(KEYINPUT80), .ZN(n549) );
  NAND2_X1 U637 ( .A1(n683), .A2(n383), .ZN(n548) );
  NAND2_X1 U638 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U639 ( .A1(KEYINPUT47), .A2(n550), .ZN(n551) );
  AND2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U641 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n591) );
  NOR2_X1 U642 ( .A1(G898), .A2(n716), .ZN(n714) );
  NAND2_X1 U643 ( .A1(n714), .A2(G902), .ZN(n556) );
  NAND2_X1 U644 ( .A1(n556), .A2(n555), .ZN(n558) );
  AND2_X1 U645 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U646 ( .A(KEYINPUT69), .B(KEYINPUT87), .ZN(n561) );
  INV_X1 U647 ( .A(n562), .ZN(n627) );
  NOR2_X1 U648 ( .A1(n627), .A2(n628), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n564), .B(KEYINPUT34), .ZN(n567) );
  XNOR2_X1 U650 ( .A(n565), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U651 ( .A1(n567), .A2(n566), .ZN(n568) );
  INV_X1 U652 ( .A(n569), .ZN(n648) );
  XNOR2_X1 U653 ( .A(n571), .B(KEYINPUT22), .ZN(n578) );
  INV_X1 U654 ( .A(n573), .ZN(n574) );
  AND2_X1 U655 ( .A1(n631), .A2(n574), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n576), .A2(n631), .ZN(n577) );
  NOR2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n582), .B(KEYINPUT85), .ZN(n583) );
  NOR2_X1 U659 ( .A1(n631), .A2(n583), .ZN(n670) );
  NOR2_X1 U660 ( .A1(n570), .A2(n638), .ZN(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT31), .B(n585), .Z(n689) );
  NOR2_X1 U662 ( .A1(n570), .A2(n586), .ZN(n675) );
  NOR2_X1 U663 ( .A1(n689), .A2(n675), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U665 ( .A1(n670), .A2(n589), .ZN(n590) );
  NAND2_X1 U666 ( .A1(KEYINPUT2), .A2(n592), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT83), .B(n593), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n594), .A2(n717), .ZN(n622) );
  NAND2_X1 U669 ( .A1(n707), .A2(G472), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n597), .B(n596), .ZN(n598) );
  NOR2_X2 U671 ( .A1(n598), .A2(n711), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(n599), .ZN(G57) );
  XOR2_X1 U673 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n602) );
  XNOR2_X1 U674 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(n603) );
  XOR2_X1 U676 ( .A(n604), .B(n603), .Z(n606) );
  NAND2_X1 U677 ( .A1(n707), .A2(G469), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X2 U679 ( .A1(n607), .A2(n711), .ZN(n609) );
  INV_X1 U680 ( .A(KEYINPUT119), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n609), .B(n608), .ZN(G54) );
  XOR2_X1 U682 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n612) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT78), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n707), .A2(G210), .ZN(n613) );
  XNOR2_X1 U686 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(G51) );
  INV_X1 U688 ( .A(n618), .ZN(n728) );
  INV_X1 U689 ( .A(n717), .ZN(n619) );
  NOR2_X1 U690 ( .A1(n728), .A2(n619), .ZN(n620) );
  NOR2_X1 U691 ( .A1(KEYINPUT2), .A2(n620), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT77), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n624), .A2(n716), .ZN(n667) );
  INV_X1 U695 ( .A(n655), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n642), .A2(n625), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT114), .ZN(n664) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U699 ( .A(KEYINPUT50), .B(n629), .ZN(n636) );
  XOR2_X1 U700 ( .A(KEYINPUT49), .B(KEYINPUT107), .Z(n633) );
  NAND2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n640) );
  XOR2_X1 U705 ( .A(KEYINPUT51), .B(KEYINPUT108), .Z(n639) );
  XNOR2_X1 U706 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U708 ( .A(n643), .B(KEYINPUT109), .ZN(n657) );
  NOR2_X1 U709 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U710 ( .A(n646), .B(KEYINPUT110), .ZN(n647) );
  NOR2_X1 U711 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U712 ( .A(n649), .B(KEYINPUT111), .ZN(n652) );
  NAND2_X1 U713 ( .A1(n650), .A2(n382), .ZN(n651) );
  NAND2_X1 U714 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U715 ( .A(KEYINPUT112), .B(n653), .Z(n654) );
  NOR2_X1 U716 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U717 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U718 ( .A(n658), .B(KEYINPUT113), .Z(n659) );
  XNOR2_X1 U719 ( .A(KEYINPUT52), .B(n659), .ZN(n660) );
  NOR2_X1 U720 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U721 ( .A1(n662), .A2(G952), .ZN(n663) );
  NAND2_X1 U722 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U723 ( .A(n665), .B(KEYINPUT115), .Z(n666) );
  NOR2_X1 U724 ( .A1(n667), .A2(n666), .ZN(n669) );
  XNOR2_X1 U725 ( .A(KEYINPUT53), .B(KEYINPUT116), .ZN(n668) );
  XOR2_X1 U726 ( .A(G101), .B(n670), .Z(G3) );
  NAND2_X1 U727 ( .A1(n675), .A2(n686), .ZN(n671) );
  XNOR2_X1 U728 ( .A(n671), .B(G104), .ZN(G6) );
  XOR2_X1 U729 ( .A(KEYINPUT27), .B(KEYINPUT103), .Z(n673) );
  XNOR2_X1 U730 ( .A(G107), .B(KEYINPUT102), .ZN(n672) );
  XNOR2_X1 U731 ( .A(n673), .B(n672), .ZN(n674) );
  XOR2_X1 U732 ( .A(KEYINPUT26), .B(n674), .Z(n677) );
  NAND2_X1 U733 ( .A1(n675), .A2(n688), .ZN(n676) );
  XNOR2_X1 U734 ( .A(n677), .B(n676), .ZN(G9) );
  XOR2_X1 U735 ( .A(G110), .B(n678), .Z(G12) );
  NOR2_X1 U736 ( .A1(n679), .A2(n683), .ZN(n681) );
  XNOR2_X1 U737 ( .A(G128), .B(KEYINPUT29), .ZN(n680) );
  XNOR2_X1 U738 ( .A(n681), .B(n680), .ZN(G30) );
  XOR2_X1 U739 ( .A(G143), .B(n682), .Z(G45) );
  INV_X1 U740 ( .A(n686), .ZN(n684) );
  NOR2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U742 ( .A(G146), .B(n685), .Z(G48) );
  NAND2_X1 U743 ( .A1(n689), .A2(n686), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n687), .B(G113), .ZN(G15) );
  NAND2_X1 U745 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U746 ( .A(n690), .B(KEYINPUT104), .ZN(n691) );
  XNOR2_X1 U747 ( .A(G116), .B(n691), .ZN(G18) );
  XNOR2_X1 U748 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n693) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U750 ( .A(G125), .B(n694), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G134), .B(KEYINPUT106), .ZN(n696) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(G36) );
  XNOR2_X1 U753 ( .A(G140), .B(n697), .ZN(G42) );
  XOR2_X1 U754 ( .A(n698), .B(KEYINPUT59), .Z(n700) );
  NAND2_X1 U755 ( .A1(n707), .A2(G475), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X2 U757 ( .A1(n701), .A2(n711), .ZN(n702) );
  XNOR2_X1 U758 ( .A(n702), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U759 ( .A1(n707), .A2(G478), .ZN(n703) );
  XNOR2_X1 U760 ( .A(n703), .B(KEYINPUT120), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n711), .A2(n706), .ZN(G63) );
  NAND2_X1 U763 ( .A1(G217), .A2(n707), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(G66) );
  XNOR2_X1 U766 ( .A(KEYINPUT123), .B(n712), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U768 ( .A(KEYINPUT124), .B(n715), .ZN(n725) );
  NAND2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT122), .ZN(n723) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n720) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n725), .B(n724), .ZN(G69) );
  XNOR2_X1 U777 ( .A(n727), .B(n726), .ZN(n731) );
  XNOR2_X1 U778 ( .A(n728), .B(n731), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(n729), .ZN(n736) );
  XNOR2_X1 U780 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n732), .A2(G900), .ZN(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT125), .B(n733), .Z(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(G72) );
  XNOR2_X1 U785 ( .A(G137), .B(n737), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n738), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U787 ( .A(G122), .B(n739), .Z(G24) );
  XOR2_X1 U788 ( .A(G119), .B(n740), .Z(G21) );
  XOR2_X1 U789 ( .A(G131), .B(n741), .Z(n742) );
  XNOR2_X1 U790 ( .A(KEYINPUT127), .B(n742), .ZN(G33) );
endmodule

