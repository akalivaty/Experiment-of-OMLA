

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792;

  INV_X1 U371 ( .A(n789), .ZN(n351) );
  INV_X1 U372 ( .A(n613), .ZN(n350) );
  AND2_X1 U373 ( .A1(n378), .A2(n376), .ZN(n375) );
  AND2_X1 U374 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U375 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U376 ( .A(n412), .B(n543), .ZN(n766) );
  XNOR2_X1 U377 ( .A(n544), .B(n542), .ZN(n412) );
  XNOR2_X2 U378 ( .A(n669), .B(KEYINPUT92), .ZN(n751) );
  XOR2_X2 U379 ( .A(n675), .B(KEYINPUT62), .Z(n676) );
  XNOR2_X2 U380 ( .A(n731), .B(KEYINPUT6), .ZN(n621) );
  AND2_X2 U381 ( .A1(n480), .A2(n479), .ZN(n478) );
  NOR2_X2 U382 ( .A1(n791), .A2(n792), .ZN(n642) );
  NAND2_X1 U383 ( .A1(n351), .A2(n350), .ZN(n411) );
  AND2_X2 U384 ( .A1(n408), .A2(n407), .ZN(n406) );
  NOR2_X2 U385 ( .A1(n374), .A2(n602), .ZN(n373) );
  XNOR2_X2 U386 ( .A(n494), .B(n493), .ZN(n658) );
  NAND2_X2 U387 ( .A1(n406), .A2(n409), .ZN(n405) );
  XNOR2_X2 U388 ( .A(n588), .B(KEYINPUT22), .ZN(n589) );
  INV_X1 U389 ( .A(n724), .ZN(n392) );
  XNOR2_X2 U390 ( .A(n630), .B(n524), .ZN(n724) );
  XNOR2_X1 U391 ( .A(G134), .B(G107), .ZN(n570) );
  AND2_X2 U392 ( .A1(n465), .A2(n657), .ZN(n472) );
  XNOR2_X2 U393 ( .A(n523), .B(n522), .ZN(n630) );
  OR2_X1 U394 ( .A1(n789), .A2(KEYINPUT44), .ZN(n371) );
  NAND2_X1 U395 ( .A1(n728), .A2(n585), .ZN(n725) );
  NOR2_X1 U396 ( .A1(n601), .A2(n600), .ZN(n640) );
  XNOR2_X1 U397 ( .A(n593), .B(n592), .ZN(n674) );
  AND2_X1 U398 ( .A1(n434), .A2(n431), .ZN(n430) );
  XNOR2_X1 U399 ( .A(n481), .B(n435), .ZN(n434) );
  NAND2_X2 U400 ( .A1(n478), .A2(n474), .ZN(n731) );
  XNOR2_X1 U401 ( .A(n569), .B(G475), .ZN(n600) );
  XNOR2_X1 U402 ( .A(n536), .B(KEYINPUT10), .ZN(n780) );
  NOR2_X1 U403 ( .A1(G237), .A2(G953), .ZN(n526) );
  NAND2_X1 U404 ( .A1(n477), .A2(n476), .ZN(n475) );
  INV_X1 U405 ( .A(n620), .ZN(n728) );
  NOR2_X1 U406 ( .A1(n646), .A2(n636), .ZN(n395) );
  NOR2_X1 U407 ( .A1(n604), .A2(n432), .ZN(n431) );
  NOR2_X1 U408 ( .A1(n621), .A2(n386), .ZN(n381) );
  NAND2_X1 U409 ( .A1(n422), .A2(n386), .ZN(n385) );
  XNOR2_X1 U410 ( .A(n511), .B(n512), .ZN(n620) );
  OR2_X1 U411 ( .A1(n762), .A2(G902), .ZN(n511) );
  INV_X1 U412 ( .A(G953), .ZN(n451) );
  INV_X1 U413 ( .A(KEYINPUT15), .ZN(n493) );
  XNOR2_X1 U414 ( .A(G902), .B(KEYINPUT93), .ZN(n494) );
  XNOR2_X1 U415 ( .A(n497), .B(n496), .ZN(n727) );
  XNOR2_X1 U416 ( .A(n554), .B(n441), .ZN(n440) );
  XNOR2_X1 U417 ( .A(n442), .B(G137), .ZN(n441) );
  INV_X1 U418 ( .A(G134), .ZN(n442) );
  INV_X1 U419 ( .A(KEYINPUT30), .ZN(n435) );
  XNOR2_X1 U420 ( .A(n490), .B(n489), .ZN(n601) );
  XNOR2_X1 U421 ( .A(n579), .B(KEYINPUT109), .ZN(n489) );
  OR2_X1 U422 ( .A1(n758), .A2(G902), .ZN(n490) );
  INV_X1 U423 ( .A(KEYINPUT86), .ZN(n389) );
  NAND2_X1 U424 ( .A1(n656), .A2(n492), .ZN(n368) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n436) );
  NAND2_X1 U426 ( .A1(n400), .A2(n352), .ZN(n398) );
  XNOR2_X1 U427 ( .A(n780), .B(n447), .ZN(n446) );
  XNOR2_X1 U428 ( .A(n504), .B(n448), .ZN(n447) );
  INV_X1 U429 ( .A(KEYINPUT23), .ZN(n504) );
  INV_X1 U430 ( .A(KEYINPUT24), .ZN(n448) );
  XNOR2_X1 U431 ( .A(n487), .B(n486), .ZN(n571) );
  XNOR2_X1 U432 ( .A(G116), .B(G122), .ZN(n486) );
  XNOR2_X1 U433 ( .A(n488), .B(KEYINPUT9), .ZN(n487) );
  XNOR2_X1 U434 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n488) );
  INV_X1 U435 ( .A(KEYINPUT7), .ZN(n573) );
  XNOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n508) );
  XNOR2_X1 U437 ( .A(n483), .B(n482), .ZN(n743) );
  XNOR2_X1 U438 ( .A(KEYINPUT117), .B(KEYINPUT41), .ZN(n482) );
  NAND2_X1 U439 ( .A1(n485), .A2(n484), .ZN(n483) );
  INV_X1 U440 ( .A(n717), .ZN(n485) );
  NAND2_X1 U441 ( .A1(n377), .A2(n387), .ZN(n376) );
  INV_X1 U442 ( .A(n455), .ZN(n456) );
  XNOR2_X1 U443 ( .A(n632), .B(KEYINPUT116), .ZN(n636) );
  XNOR2_X1 U444 ( .A(n629), .B(n413), .ZN(n631) );
  XNOR2_X1 U445 ( .A(KEYINPUT115), .B(KEYINPUT28), .ZN(n413) );
  OR2_X1 U446 ( .A1(n415), .A2(KEYINPUT87), .ZN(n461) );
  NOR2_X1 U447 ( .A1(KEYINPUT47), .A2(n648), .ZN(n650) );
  XNOR2_X1 U448 ( .A(n364), .B(KEYINPUT88), .ZN(n611) );
  NAND2_X1 U449 ( .A1(n599), .A2(n674), .ZN(n364) );
  XNOR2_X1 U450 ( .A(n443), .B(G131), .ZN(n554) );
  INV_X1 U451 ( .A(KEYINPUT70), .ZN(n443) );
  XNOR2_X1 U452 ( .A(n495), .B(n423), .ZN(n499) );
  XNOR2_X1 U453 ( .A(KEYINPUT20), .B(KEYINPUT98), .ZN(n423) );
  XNOR2_X1 U454 ( .A(G122), .B(KEYINPUT12), .ZN(n560) );
  XOR2_X1 U455 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n561) );
  XNOR2_X1 U456 ( .A(n780), .B(n554), .ZN(n558) );
  XNOR2_X1 U457 ( .A(G143), .B(G113), .ZN(n556) );
  XOR2_X1 U458 ( .A(G140), .B(G104), .Z(n555) );
  XOR2_X1 U459 ( .A(KEYINPUT71), .B(G140), .Z(n516) );
  NOR2_X1 U460 ( .A1(n368), .A2(n658), .ZN(n467) );
  NAND2_X1 U461 ( .A1(n451), .A2(G224), .ZN(n450) );
  XNOR2_X1 U462 ( .A(n396), .B(KEYINPUT18), .ZN(n534) );
  INV_X1 U463 ( .A(KEYINPUT90), .ZN(n396) );
  XNOR2_X1 U464 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n514) );
  NAND2_X1 U465 ( .A1(G234), .A2(G237), .ZN(n548) );
  XNOR2_X1 U466 ( .A(n456), .B(KEYINPUT38), .ZN(n715) );
  AND2_X1 U467 ( .A1(n620), .A2(n619), .ZN(n628) );
  INV_X1 U468 ( .A(G237), .ZN(n545) );
  INV_X1 U469 ( .A(n718), .ZN(n484) );
  INV_X1 U470 ( .A(n725), .ZN(n391) );
  INV_X1 U471 ( .A(KEYINPUT33), .ZN(n386) );
  INV_X1 U472 ( .A(n383), .ZN(n379) );
  INV_X1 U473 ( .A(n604), .ZN(n428) );
  NOR2_X1 U474 ( .A1(n753), .A2(G902), .ZN(n523) );
  XNOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT102), .ZN(n525) );
  INV_X1 U476 ( .A(n368), .ZN(n367) );
  XNOR2_X1 U477 ( .A(n639), .B(n491), .ZN(n651) );
  INV_X1 U478 ( .A(n433), .ZN(n429) );
  NOR2_X1 U479 ( .A1(n415), .A2(n728), .ZN(n590) );
  INV_X1 U480 ( .A(G953), .ZN(n782) );
  XNOR2_X1 U481 ( .A(n368), .B(n784), .ZN(n783) );
  XNOR2_X1 U482 ( .A(n445), .B(n444), .ZN(n762) );
  XNOR2_X1 U483 ( .A(n505), .B(n510), .ZN(n444) );
  XNOR2_X1 U484 ( .A(n446), .B(n507), .ZN(n445) );
  XNOR2_X1 U485 ( .A(n578), .B(n357), .ZN(n758) );
  XNOR2_X1 U486 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U487 ( .A1(n636), .A2(n743), .ZN(n637) );
  NAND2_X1 U488 ( .A1(n375), .A2(n372), .ZN(n582) );
  XNOR2_X1 U489 ( .A(n370), .B(KEYINPUT114), .ZN(n790) );
  AND2_X1 U490 ( .A1(n473), .A2(n420), .ZN(n419) );
  INV_X1 U491 ( .A(n456), .ZN(n420) );
  BUF_X1 U492 ( .A(n705), .Z(n421) );
  NAND2_X1 U493 ( .A1(n459), .A2(n458), .ZN(n457) );
  INV_X1 U494 ( .A(KEYINPUT87), .ZN(n458) );
  INV_X1 U495 ( .A(n658), .ZN(n471) );
  BUF_X1 U496 ( .A(n724), .Z(n415) );
  AND2_X1 U497 ( .A1(n410), .A2(n399), .ZN(n352) );
  OR2_X1 U498 ( .A1(n618), .A2(n617), .ZN(n353) );
  INV_X1 U499 ( .A(n388), .ZN(n660) );
  OR2_X1 U500 ( .A1(KEYINPUT80), .A2(n719), .ZN(n354) );
  AND2_X1 U501 ( .A1(n585), .A2(n353), .ZN(n355) );
  NAND2_X1 U502 ( .A1(n369), .A2(n354), .ZN(n356) );
  XOR2_X1 U503 ( .A(n581), .B(KEYINPUT112), .Z(n649) );
  NAND2_X1 U504 ( .A1(n392), .A2(n391), .ZN(n422) );
  AND2_X1 U505 ( .A1(n577), .A2(G217), .ZN(n357) );
  AND2_X1 U506 ( .A1(n546), .A2(G210), .ZN(n358) );
  AND2_X1 U507 ( .A1(n590), .A2(n621), .ZN(n359) );
  AND2_X1 U508 ( .A1(n635), .A2(KEYINPUT47), .ZN(n360) );
  INV_X1 U509 ( .A(G902), .ZN(n476) );
  AND2_X1 U510 ( .A1(n461), .A2(n728), .ZN(n361) );
  AND2_X1 U511 ( .A1(n614), .A2(KEYINPUT66), .ZN(n362) );
  INV_X1 U512 ( .A(KEYINPUT34), .ZN(n387) );
  NAND2_X1 U513 ( .A1(KEYINPUT84), .A2(n471), .ZN(n363) );
  NAND2_X1 U514 ( .A1(n367), .A2(n365), .ZN(n388) );
  NAND2_X1 U515 ( .A1(n365), .A2(n782), .ZN(n774) );
  NAND2_X1 U516 ( .A1(n467), .A2(n365), .ZN(n470) );
  NAND2_X1 U517 ( .A1(n466), .A2(n365), .ZN(n465) );
  NAND2_X2 U518 ( .A1(n401), .A2(n398), .ZN(n365) );
  XNOR2_X2 U519 ( .A(n366), .B(n532), .ZN(n675) );
  XNOR2_X1 U520 ( .A(n366), .B(n520), .ZN(n753) );
  XNOR2_X2 U521 ( .A(n779), .B(n515), .ZN(n366) );
  NOR2_X1 U522 ( .A1(n368), .A2(n363), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n790), .B(KEYINPUT82), .ZN(n369) );
  NAND2_X1 U524 ( .A1(n419), .A2(n649), .ZN(n370) );
  NAND2_X1 U525 ( .A1(n371), .A2(KEYINPUT66), .ZN(n394) );
  XNOR2_X2 U526 ( .A(n583), .B(KEYINPUT35), .ZN(n789) );
  NAND2_X1 U527 ( .A1(n383), .A2(n380), .ZN(n722) );
  NAND2_X1 U528 ( .A1(n373), .A2(n383), .ZN(n372) );
  NAND2_X1 U529 ( .A1(n380), .A2(KEYINPUT34), .ZN(n374) );
  NAND2_X1 U530 ( .A1(n397), .A2(n380), .ZN(n377) );
  NAND2_X1 U531 ( .A1(n379), .A2(n387), .ZN(n378) );
  INV_X1 U532 ( .A(n422), .ZN(n382) );
  NAND2_X1 U533 ( .A1(n621), .A2(n386), .ZN(n384) );
  NAND2_X1 U534 ( .A1(n595), .A2(n621), .ZN(n390) );
  NAND2_X1 U535 ( .A1(n595), .A2(n359), .ZN(n593) );
  XNOR2_X1 U536 ( .A(n390), .B(n389), .ZN(n464) );
  NAND2_X1 U537 ( .A1(n411), .A2(n614), .ZN(n407) );
  NAND2_X1 U538 ( .A1(n394), .A2(n393), .ZN(n409) );
  INV_X1 U539 ( .A(n611), .ZN(n393) );
  XNOR2_X1 U540 ( .A(n535), .B(n536), .ZN(n537) );
  XNOR2_X2 U541 ( .A(n425), .B(G101), .ZN(n535) );
  XNOR2_X1 U542 ( .A(n437), .B(n436), .ZN(n656) );
  NOR2_X1 U543 ( .A1(n650), .A2(n360), .ZN(n418) );
  NOR2_X1 U544 ( .A1(n356), .A2(n417), .ZN(n439) );
  NOR2_X1 U545 ( .A1(n395), .A2(n647), .ZN(n648) );
  NAND2_X1 U546 ( .A1(n403), .A2(KEYINPUT45), .ZN(n402) );
  INV_X1 U547 ( .A(n397), .ZN(n602) );
  NAND2_X1 U548 ( .A1(n587), .A2(n397), .ZN(n416) );
  XNOR2_X2 U549 ( .A(n424), .B(KEYINPUT0), .ZN(n397) );
  NAND2_X1 U550 ( .A1(n397), .A2(n606), .ZN(n693) );
  INV_X1 U551 ( .A(KEYINPUT45), .ZN(n399) );
  INV_X1 U552 ( .A(n405), .ZN(n400) );
  AND2_X2 U553 ( .A1(n404), .A2(n402), .ZN(n401) );
  INV_X1 U554 ( .A(n410), .ZN(n403) );
  NAND2_X1 U555 ( .A1(n405), .A2(KEYINPUT45), .ZN(n404) );
  NAND2_X1 U556 ( .A1(n611), .A2(n362), .ZN(n408) );
  XNOR2_X2 U557 ( .A(n610), .B(KEYINPUT111), .ZN(n410) );
  NOR2_X2 U558 ( .A1(G953), .A2(KEYINPUT17), .ZN(n449) );
  INV_X2 U559 ( .A(KEYINPUT69), .ZN(n425) );
  NAND2_X1 U560 ( .A1(n452), .A2(n453), .ZN(n454) );
  NAND2_X1 U561 ( .A1(n450), .A2(KEYINPUT17), .ZN(n453) );
  XNOR2_X2 U562 ( .A(n517), .B(G104), .ZN(n544) );
  NAND2_X1 U563 ( .A1(n449), .A2(G224), .ZN(n452) );
  NAND2_X1 U564 ( .A1(n598), .A2(n620), .ZN(n599) );
  XNOR2_X1 U565 ( .A(n414), .B(n766), .ZN(n665) );
  XNOR2_X1 U566 ( .A(n539), .B(n540), .ZN(n414) );
  INV_X1 U567 ( .A(n599), .ZN(n696) );
  NAND2_X1 U568 ( .A1(n651), .A2(n640), .ZN(n641) );
  NAND2_X1 U569 ( .A1(n430), .A2(n429), .ZN(n639) );
  NOR2_X1 U570 ( .A1(n681), .A2(G902), .ZN(n568) );
  XNOR2_X1 U571 ( .A(n565), .B(n566), .ZN(n681) );
  XNOR2_X2 U572 ( .A(n416), .B(n589), .ZN(n595) );
  NAND2_X1 U573 ( .A1(n455), .A2(n714), .ZN(n623) );
  NAND2_X1 U574 ( .A1(n418), .A2(n712), .ZN(n417) );
  NOR2_X2 U575 ( .A1(n702), .A2(n553), .ZN(n424) );
  XNOR2_X2 U576 ( .A(n426), .B(n358), .ZN(n455) );
  NAND2_X1 U577 ( .A1(n665), .A2(n658), .ZN(n426) );
  NOR2_X1 U578 ( .A1(n427), .A2(n433), .ZN(n473) );
  NAND2_X1 U579 ( .A1(n434), .A2(n428), .ZN(n427) );
  INV_X1 U580 ( .A(n715), .ZN(n432) );
  NOR2_X1 U581 ( .A1(n604), .A2(n725), .ZN(n638) );
  NAND2_X1 U582 ( .A1(n355), .A2(n728), .ZN(n433) );
  NAND2_X1 U583 ( .A1(n439), .A2(n438), .ZN(n437) );
  XNOR2_X1 U584 ( .A(n642), .B(KEYINPUT46), .ZN(n438) );
  XNOR2_X2 U585 ( .A(n539), .B(n440), .ZN(n779) );
  XNOR2_X1 U586 ( .A(n454), .B(n534), .ZN(n538) );
  NAND2_X1 U587 ( .A1(n655), .A2(n456), .ZN(n673) );
  NAND2_X2 U588 ( .A1(n460), .A2(n457), .ZN(n687) );
  INV_X1 U589 ( .A(n464), .ZN(n459) );
  AND2_X2 U590 ( .A1(n462), .A2(n361), .ZN(n460) );
  NAND2_X1 U591 ( .A1(n464), .A2(n463), .ZN(n462) );
  AND2_X1 U592 ( .A1(n415), .A2(KEYINPUT87), .ZN(n463) );
  NAND2_X1 U593 ( .A1(n472), .A2(n468), .ZN(n659) );
  NAND2_X1 U594 ( .A1(n470), .A2(n469), .ZN(n468) );
  INV_X1 U595 ( .A(KEYINPUT84), .ZN(n469) );
  OR2_X1 U596 ( .A1(n675), .A2(n475), .ZN(n474) );
  INV_X1 U597 ( .A(n533), .ZN(n477) );
  NAND2_X1 U598 ( .A1(n533), .A2(G902), .ZN(n479) );
  NAND2_X1 U599 ( .A1(n675), .A2(n533), .ZN(n480) );
  NAND2_X1 U600 ( .A1(n731), .A2(n714), .ZN(n481) );
  XNOR2_X2 U601 ( .A(n572), .B(n514), .ZN(n539) );
  XNOR2_X2 U602 ( .A(G146), .B(G125), .ZN(n536) );
  XOR2_X1 U603 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n491) );
  AND2_X1 U604 ( .A1(n713), .A2(n673), .ZN(n492) );
  AND2_X1 U605 ( .A1(n727), .A2(n353), .ZN(n619) );
  XNOR2_X1 U606 ( .A(n535), .B(G146), .ZN(n515) );
  XNOR2_X1 U607 ( .A(n521), .B(G469), .ZN(n522) );
  XNOR2_X1 U608 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U609 ( .A(n576), .B(n575), .ZN(n578) );
  XNOR2_X1 U610 ( .A(n753), .B(n754), .ZN(n755) );
  XNOR2_X1 U611 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U612 ( .A1(n658), .A2(G234), .ZN(n495) );
  NAND2_X1 U613 ( .A1(G221), .A2(n499), .ZN(n497) );
  XOR2_X1 U614 ( .A(KEYINPUT100), .B(KEYINPUT21), .Z(n496) );
  INV_X1 U615 ( .A(KEYINPUT101), .ZN(n498) );
  XNOR2_X1 U616 ( .A(n727), .B(n498), .ZN(n585) );
  XOR2_X1 U617 ( .A(KEYINPUT25), .B(KEYINPUT99), .Z(n501) );
  NAND2_X1 U618 ( .A1(G217), .A2(n499), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n501), .B(n500), .ZN(n512) );
  XOR2_X1 U620 ( .A(G110), .B(G119), .Z(n503) );
  XNOR2_X1 U621 ( .A(G137), .B(G128), .ZN(n502) );
  XNOR2_X1 U622 ( .A(n503), .B(n502), .ZN(n505) );
  INV_X1 U623 ( .A(n516), .ZN(n506) );
  XOR2_X1 U624 ( .A(n506), .B(KEYINPUT97), .Z(n507) );
  NAND2_X1 U625 ( .A1(n782), .A2(G234), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n509), .B(n508), .ZN(n577) );
  NAND2_X1 U627 ( .A1(n577), .A2(G221), .ZN(n510) );
  XNOR2_X2 U628 ( .A(G128), .B(KEYINPUT79), .ZN(n513) );
  XNOR2_X2 U629 ( .A(n513), .B(G143), .ZN(n572) );
  XOR2_X1 U630 ( .A(KEYINPUT96), .B(n516), .Z(n778) );
  NAND2_X1 U631 ( .A1(G227), .A2(n782), .ZN(n518) );
  XNOR2_X2 U632 ( .A(G110), .B(G107), .ZN(n517) );
  XOR2_X1 U633 ( .A(n518), .B(n544), .Z(n519) );
  XNOR2_X1 U634 ( .A(n778), .B(n519), .ZN(n520) );
  INV_X1 U635 ( .A(KEYINPUT72), .ZN(n521) );
  INV_X1 U636 ( .A(KEYINPUT1), .ZN(n524) );
  XNOR2_X1 U637 ( .A(n525), .B(KEYINPUT77), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n526), .B(KEYINPUT78), .ZN(n559) );
  NAND2_X1 U639 ( .A1(G210), .A2(n559), .ZN(n527) );
  XNOR2_X1 U640 ( .A(n528), .B(n527), .ZN(n531) );
  XNOR2_X1 U641 ( .A(G116), .B(G113), .ZN(n530) );
  XNOR2_X1 U642 ( .A(KEYINPUT3), .B(G119), .ZN(n529) );
  XNOR2_X1 U643 ( .A(n530), .B(n529), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n543), .B(n531), .ZN(n532) );
  XOR2_X1 U645 ( .A(G472), .B(KEYINPUT73), .Z(n533) );
  XNOR2_X1 U646 ( .A(n537), .B(n538), .ZN(n540) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n541) );
  XNOR2_X1 U648 ( .A(n541), .B(G122), .ZN(n542) );
  NAND2_X1 U649 ( .A1(n476), .A2(n545), .ZN(n546) );
  NAND2_X1 U650 ( .A1(n546), .A2(G214), .ZN(n714) );
  INV_X1 U651 ( .A(KEYINPUT19), .ZN(n547) );
  XNOR2_X2 U652 ( .A(n623), .B(n547), .ZN(n702) );
  XNOR2_X1 U653 ( .A(n548), .B(KEYINPUT14), .ZN(n549) );
  XNOR2_X1 U654 ( .A(KEYINPUT76), .B(n549), .ZN(n550) );
  NAND2_X1 U655 ( .A1(G952), .A2(n550), .ZN(n742) );
  NOR2_X1 U656 ( .A1(G953), .A2(n742), .ZN(n618) );
  NAND2_X1 U657 ( .A1(n550), .A2(G902), .ZN(n615) );
  XOR2_X1 U658 ( .A(KEYINPUT94), .B(G898), .Z(n771) );
  NAND2_X1 U659 ( .A1(G953), .A2(n771), .ZN(n767) );
  NOR2_X1 U660 ( .A1(n615), .A2(n767), .ZN(n551) );
  OR2_X1 U661 ( .A1(n618), .A2(n551), .ZN(n552) );
  XNOR2_X1 U662 ( .A(n552), .B(KEYINPUT95), .ZN(n553) );
  XNOR2_X1 U663 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U664 ( .A(n558), .B(n557), .ZN(n566) );
  NAND2_X1 U665 ( .A1(n559), .A2(G214), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U667 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U668 ( .A(n564), .B(KEYINPUT11), .Z(n565) );
  XNOR2_X1 U669 ( .A(KEYINPUT13), .B(KEYINPUT105), .ZN(n567) );
  XNOR2_X1 U670 ( .A(n568), .B(n567), .ZN(n569) );
  INV_X1 U671 ( .A(n600), .ZN(n580) );
  XNOR2_X1 U672 ( .A(n571), .B(n570), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n572), .B(KEYINPUT108), .ZN(n574) );
  INV_X1 U674 ( .A(G478), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n580), .A2(n601), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n582), .A2(n649), .ZN(n583) );
  INV_X1 U677 ( .A(n601), .ZN(n584) );
  NAND2_X1 U678 ( .A1(n584), .A2(n600), .ZN(n717) );
  INV_X1 U679 ( .A(n585), .ZN(n586) );
  NOR2_X1 U680 ( .A1(n717), .A2(n586), .ZN(n587) );
  INV_X1 U681 ( .A(KEYINPUT74), .ZN(n588) );
  INV_X1 U682 ( .A(KEYINPUT67), .ZN(n591) );
  XNOR2_X1 U683 ( .A(n591), .B(KEYINPUT32), .ZN(n592) );
  INV_X1 U684 ( .A(n731), .ZN(n605) );
  AND2_X1 U685 ( .A1(n415), .A2(n605), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U687 ( .A(KEYINPUT68), .ZN(n596) );
  XNOR2_X1 U688 ( .A(n597), .B(n596), .ZN(n598) );
  AND2_X1 U689 ( .A1(n601), .A2(n600), .ZN(n692) );
  NOR2_X1 U690 ( .A1(n692), .A2(n640), .ZN(n719) );
  XNOR2_X1 U691 ( .A(n719), .B(KEYINPUT81), .ZN(n645) );
  NAND2_X1 U692 ( .A1(n382), .A2(n731), .ZN(n734) );
  NOR2_X1 U693 ( .A1(n734), .A2(n602), .ZN(n603) );
  XNOR2_X1 U694 ( .A(n603), .B(KEYINPUT31), .ZN(n707) );
  INV_X1 U695 ( .A(n630), .ZN(n604) );
  AND2_X1 U696 ( .A1(n638), .A2(n605), .ZN(n606) );
  NAND2_X1 U697 ( .A1(n707), .A2(n693), .ZN(n607) );
  NAND2_X1 U698 ( .A1(n645), .A2(n607), .ZN(n608) );
  XNOR2_X1 U699 ( .A(n608), .B(KEYINPUT110), .ZN(n609) );
  NAND2_X1 U700 ( .A1(n687), .A2(n609), .ZN(n610) );
  INV_X1 U701 ( .A(KEYINPUT44), .ZN(n613) );
  NAND2_X1 U702 ( .A1(n613), .A2(KEYINPUT66), .ZN(n614) );
  OR2_X1 U703 ( .A1(n782), .A2(n615), .ZN(n616) );
  NOR2_X1 U704 ( .A1(G900), .A2(n616), .ZN(n617) );
  XNOR2_X1 U705 ( .A(n640), .B(KEYINPUT113), .ZN(n705) );
  NOR2_X1 U706 ( .A1(n621), .A2(n705), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n628), .A2(n622), .ZN(n652) );
  XNOR2_X1 U708 ( .A(KEYINPUT118), .B(n652), .ZN(n624) );
  NOR2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n626) );
  XOR2_X1 U710 ( .A(KEYINPUT36), .B(KEYINPUT89), .Z(n625) );
  XNOR2_X1 U711 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n627), .A2(n392), .ZN(n712) );
  NAND2_X1 U713 ( .A1(n628), .A2(n731), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n631), .A2(n428), .ZN(n632) );
  INV_X1 U715 ( .A(n636), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n719), .A2(KEYINPUT80), .ZN(n633) );
  INV_X1 U717 ( .A(n702), .ZN(n644) );
  AND2_X1 U718 ( .A1(n633), .A2(n644), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n643), .A2(n634), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n715), .A2(n714), .ZN(n718) );
  XNOR2_X1 U721 ( .A(n637), .B(KEYINPUT42), .ZN(n792) );
  XOR2_X1 U722 ( .A(KEYINPUT40), .B(n641), .Z(n791) );
  INV_X1 U723 ( .A(KEYINPUT80), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n651), .A2(n692), .ZN(n713) );
  NOR2_X1 U726 ( .A1(n392), .A2(n652), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n653), .A2(n714), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT43), .ZN(n655) );
  INV_X1 U729 ( .A(KEYINPUT2), .ZN(n661) );
  OR2_X1 U730 ( .A1(n658), .A2(n661), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT65), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n388), .A2(n661), .ZN(n662) );
  NOR2_X2 U733 ( .A1(n663), .A2(n662), .ZN(n752) );
  NAND2_X1 U734 ( .A1(n752), .A2(G210), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n664) );
  XNOR2_X1 U736 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(n670) );
  INV_X1 U738 ( .A(G952), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n668), .A2(G953), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n670), .A2(n751), .ZN(n672) );
  INV_X1 U741 ( .A(KEYINPUT56), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G51) );
  XNOR2_X1 U743 ( .A(n673), .B(G140), .ZN(G42) );
  XNOR2_X1 U744 ( .A(n674), .B(G119), .ZN(G21) );
  NAND2_X1 U745 ( .A1(n752), .A2(G472), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n678), .A2(n751), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n679), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U749 ( .A1(n752), .A2(G475), .ZN(n683) );
  XOR2_X1 U750 ( .A(KEYINPUT91), .B(KEYINPUT59), .Z(n680) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n684), .A2(n751), .ZN(n686) );
  XNOR2_X1 U753 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n685) );
  XNOR2_X1 U754 ( .A(n686), .B(n685), .ZN(G60) );
  XNOR2_X1 U755 ( .A(n687), .B(G101), .ZN(G3) );
  NOR2_X1 U756 ( .A1(n421), .A2(n693), .ZN(n689) );
  XNOR2_X1 U757 ( .A(G104), .B(KEYINPUT119), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n689), .B(n688), .ZN(G6) );
  XOR2_X1 U759 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n691) );
  XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT120), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n691), .B(n690), .ZN(n695) );
  INV_X1 U762 ( .A(n692), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n708), .A2(n693), .ZN(n694) );
  XOR2_X1 U764 ( .A(n695), .B(n694), .Z(G9) );
  XNOR2_X1 U765 ( .A(n696), .B(G110), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(KEYINPUT121), .ZN(G12) );
  XOR2_X1 U767 ( .A(KEYINPUT29), .B(KEYINPUT122), .Z(n700) );
  NOR2_X1 U768 ( .A1(n708), .A2(n702), .ZN(n698) );
  NAND2_X1 U769 ( .A1(n643), .A2(n698), .ZN(n699) );
  XNOR2_X1 U770 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U771 ( .A(G128), .B(n701), .ZN(G30) );
  NOR2_X1 U772 ( .A1(n421), .A2(n702), .ZN(n703) );
  AND2_X1 U773 ( .A1(n643), .A2(n703), .ZN(n704) );
  XOR2_X1 U774 ( .A(G146), .B(n704), .Z(G48) );
  NOR2_X1 U775 ( .A1(n421), .A2(n707), .ZN(n706) );
  XOR2_X1 U776 ( .A(G113), .B(n706), .Z(G15) );
  NOR2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U778 ( .A(G116), .B(KEYINPUT123), .ZN(n709) );
  XNOR2_X1 U779 ( .A(n710), .B(n709), .ZN(G18) );
  XOR2_X1 U780 ( .A(G125), .B(KEYINPUT37), .Z(n711) );
  XNOR2_X1 U781 ( .A(n712), .B(n711), .ZN(G27) );
  XNOR2_X1 U782 ( .A(G134), .B(n713), .ZN(G36) );
  XNOR2_X1 U783 ( .A(n660), .B(KEYINPUT2), .ZN(n748) );
  NOR2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n739) );
  NAND2_X1 U789 ( .A1(n725), .A2(n415), .ZN(n726) );
  XNOR2_X1 U790 ( .A(n726), .B(KEYINPUT50), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U792 ( .A(KEYINPUT49), .B(n729), .Z(n730) );
  NOR2_X1 U793 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U794 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U795 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U796 ( .A(KEYINPUT51), .B(n736), .ZN(n737) );
  NOR2_X1 U797 ( .A1(n737), .A2(n743), .ZN(n738) );
  NOR2_X1 U798 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U799 ( .A(n740), .B(KEYINPUT52), .ZN(n741) );
  NOR2_X1 U800 ( .A1(n742), .A2(n741), .ZN(n746) );
  NOR2_X1 U801 ( .A1(n722), .A2(n743), .ZN(n744) );
  XNOR2_X1 U802 ( .A(KEYINPUT124), .B(n744), .ZN(n745) );
  NOR2_X1 U803 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U804 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U805 ( .A1(n749), .A2(G953), .ZN(n750) );
  XNOR2_X1 U806 ( .A(n750), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U807 ( .A(n751), .ZN(n765) );
  BUF_X2 U808 ( .A(n752), .Z(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(G469), .ZN(n756) );
  XOR2_X1 U810 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n754) );
  NOR2_X1 U811 ( .A1(n765), .A2(n757), .ZN(G54) );
  NAND2_X1 U812 ( .A1(n761), .A2(G478), .ZN(n759) );
  XNOR2_X1 U813 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n765), .A2(n760), .ZN(G63) );
  NAND2_X1 U815 ( .A1(n761), .A2(G217), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U817 ( .A1(n765), .A2(n764), .ZN(G66) );
  XNOR2_X1 U818 ( .A(n766), .B(G101), .ZN(n768) );
  NAND2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n777) );
  NAND2_X1 U820 ( .A1(G953), .A2(G224), .ZN(n769) );
  XOR2_X1 U821 ( .A(KEYINPUT61), .B(n769), .Z(n770) );
  NOR2_X1 U822 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U823 ( .A(KEYINPUT126), .B(n772), .Z(n773) );
  NAND2_X1 U824 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U825 ( .A(n775), .B(KEYINPUT127), .ZN(n776) );
  XNOR2_X1 U826 ( .A(n777), .B(n776), .ZN(G69) );
  XNOR2_X1 U827 ( .A(n779), .B(n778), .ZN(n781) );
  XOR2_X1 U828 ( .A(n780), .B(n781), .Z(n784) );
  NAND2_X1 U829 ( .A1(n783), .A2(n782), .ZN(n788) );
  XNOR2_X1 U830 ( .A(G227), .B(n784), .ZN(n785) );
  NAND2_X1 U831 ( .A1(n785), .A2(G900), .ZN(n786) );
  NAND2_X1 U832 ( .A1(G953), .A2(n786), .ZN(n787) );
  NAND2_X1 U833 ( .A1(n788), .A2(n787), .ZN(G72) );
  XOR2_X1 U834 ( .A(n789), .B(G122), .Z(G24) );
  XNOR2_X1 U835 ( .A(G143), .B(n790), .ZN(G45) );
  XOR2_X1 U836 ( .A(G131), .B(n791), .Z(G33) );
  XOR2_X1 U837 ( .A(G137), .B(n792), .Z(G39) );
endmodule

