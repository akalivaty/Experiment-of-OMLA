//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT67), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n209), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G50), .A2(G226), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n207), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n207), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT0), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n227), .A2(G1), .A3(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n222), .A2(new_n223), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n224), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n220), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(G270), .Z(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G226), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n240), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G107), .ZN(new_n253));
  INV_X1    g0053(.A(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n251), .B(new_n255), .Z(G351));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n258), .A2(KEYINPUT77), .B1(new_n260), .B2(G77), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n261), .B1(KEYINPUT77), .B2(new_n258), .C1(new_n230), .C2(G68), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n207), .A2(new_n259), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n229), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(KEYINPUT11), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n226), .B2(new_n228), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G20), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G68), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT71), .B(G1), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n277), .A2(new_n278), .A3(new_n230), .ZN(new_n279));
  INV_X1    g0079(.A(G68), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT12), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n262), .A2(new_n265), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n276), .B(new_n282), .C1(KEYINPUT11), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G232), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G226), .B2(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n287), .A2(new_n291), .B1(new_n259), .B2(new_n212), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n259), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n229), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n225), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(G45), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n272), .A2(G41), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(G238), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n293), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT70), .A2(G41), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n268), .B(G274), .C1(new_n305), .C2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n296), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT13), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n296), .A2(new_n301), .A3(new_n309), .A4(new_n306), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n308), .A2(G190), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n308), .B2(new_n310), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n284), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n274), .A2(G77), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n257), .A2(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n257), .A2(KEYINPUT74), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT75), .ZN(new_n323));
  OR2_X1    g0123(.A1(KEYINPUT15), .A2(G87), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g0125(.A1(KEYINPUT15), .A2(G87), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n260), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G20), .B2(G77), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n315), .B1(G77), .B2(new_n316), .C1(new_n331), .C2(new_n267), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT3), .B(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G238), .A3(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G107), .ZN(new_n335));
  INV_X1    g0135(.A(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n334), .B1(new_n335), .B2(new_n333), .C1(new_n337), .C2(new_n285), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n295), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G244), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n306), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n332), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n308), .B2(new_n310), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n351), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n308), .A2(G179), .A3(new_n310), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n352), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n314), .B(new_n349), .C1(new_n357), .C2(new_n284), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n274), .A2(G50), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  INV_X1    g0160(.A(new_n257), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n317), .A2(new_n329), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(G20), .B2(new_n203), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n359), .B1(G50), .B2(new_n316), .C1(new_n363), .C2(new_n267), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT9), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n340), .A2(G226), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT72), .A2(G223), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT72), .A2(G223), .ZN(new_n369));
  OAI21_X1  g0169(.A(G1698), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n336), .A2(G222), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n333), .A3(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n295), .C1(G77), .C2(new_n333), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n306), .A3(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n364), .A2(new_n365), .B1(new_n374), .B2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n374), .A2(KEYINPUT76), .A3(new_n376), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n366), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(new_n346), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n374), .A2(G179), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n386), .A2(KEYINPUT73), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(KEYINPUT73), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n364), .B(new_n385), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n332), .B1(G200), .B2(new_n342), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n343), .A2(G190), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND4_X1   g0192(.A1(new_n383), .A2(new_n384), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n340), .A2(G232), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n333), .A2(G226), .A3(G1698), .ZN(new_n395));
  INV_X1    g0195(.A(G223), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n337), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n259), .A2(new_n210), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n295), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n399), .A3(new_n306), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n346), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n400), .A2(G179), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n230), .B1(new_n232), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n333), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n404), .B1(new_n408), .B2(G68), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n361), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT16), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n280), .B1(new_n406), .B2(new_n407), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n414), .A2(new_n415), .A3(new_n411), .A4(new_n404), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n413), .A2(new_n416), .A3(new_n267), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n273), .A2(new_n318), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT79), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n279), .A2(new_n265), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n420), .A2(new_n421), .B1(new_n279), .B2(new_n317), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n401), .B(new_n402), .C1(new_n417), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n333), .A2(new_n405), .A3(G20), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT7), .B1(new_n291), .B2(new_n230), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n404), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n412), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n415), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n409), .A2(KEYINPUT16), .A3(new_n412), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n265), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n422), .B1(new_n346), .B2(new_n400), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT18), .B1(new_n435), .B2(new_n402), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n400), .A2(G200), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n394), .A2(new_n399), .A3(G190), .A4(new_n306), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n434), .A2(new_n422), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(KEYINPUT17), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(KEYINPUT17), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n426), .A2(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT80), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n424), .A2(new_n425), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n402), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n434), .A2(new_n422), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n437), .A4(new_n438), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(KEYINPUT17), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n445), .A2(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT80), .ZN(new_n452));
  AND4_X1   g0252(.A1(new_n358), .A2(new_n393), .A3(new_n444), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n303), .A2(new_n455), .A3(new_n304), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n272), .A3(G45), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G264), .A3(new_n298), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n288), .A2(new_n290), .A3(G257), .A4(G1698), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n288), .A2(new_n290), .A3(G250), .A4(new_n336), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G294), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n295), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n269), .B2(new_n271), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(new_n456), .A3(G274), .A4(new_n457), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n297), .ZN(new_n469));
  OAI21_X1  g0269(.A(G169), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n459), .A2(KEYINPUT87), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n468), .A2(new_n297), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT87), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n458), .A2(new_n473), .A3(G264), .A4(new_n298), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n464), .A4(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n470), .B1(new_n475), .B2(new_n344), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n470), .B(KEYINPUT88), .C1(new_n475), .C2(new_n344), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n333), .A2(new_n230), .A3(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n333), .A2(new_n483), .A3(new_n230), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n260), .A2(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n230), .A2(G107), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT23), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n485), .A2(new_n491), .A3(new_n486), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n265), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n272), .A2(G33), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n316), .A2(new_n267), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n316), .A2(G107), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n480), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n475), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n472), .A2(new_n459), .A3(new_n464), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n503), .A2(G200), .B1(G190), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n498), .A3(new_n494), .A4(new_n500), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n288), .A2(new_n290), .A3(G244), .A4(new_n336), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n333), .A2(G250), .A3(G1698), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n333), .A2(G244), .A3(new_n336), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n510), .A2(new_n511), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(new_n295), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n458), .A2(G257), .A3(new_n298), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n297), .B2(new_n468), .ZN(new_n518));
  OAI21_X1  g0318(.A(G200), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n316), .A2(G97), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n408), .A2(G107), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT81), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT6), .A2(G97), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(G107), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n335), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(G97), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n212), .A2(new_n335), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G20), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n361), .A2(new_n250), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n521), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n520), .B1(new_n535), .B2(new_n265), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n497), .A2(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n515), .A2(new_n295), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(G190), .A3(new_n472), .A4(new_n517), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n519), .A2(new_n536), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n520), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n335), .B1(new_n406), .B2(new_n407), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n230), .B1(new_n526), .B2(new_n530), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n542), .A2(new_n543), .A3(new_n533), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n541), .B(new_n537), .C1(new_n544), .C2(new_n267), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n346), .B1(new_n516), .B2(new_n518), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n538), .A2(new_n344), .A3(new_n472), .A4(new_n517), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n502), .A2(new_n506), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT84), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n323), .A2(new_n327), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n421), .A2(new_n551), .A3(new_n552), .A4(new_n495), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT84), .B1(new_n496), .B2(new_n328), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n328), .A2(new_n279), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n333), .A2(new_n230), .A3(G68), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n260), .A2(G97), .ZN(new_n557));
  OR2_X1    g0357(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n558));
  NAND2_X1  g0358(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(G33), .A3(G97), .A4(new_n559), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n230), .B1(new_n210), .B2(new_n529), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n265), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n288), .A2(new_n290), .A3(G244), .A4(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n288), .A2(new_n290), .A3(G238), .A4(new_n336), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G116), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n295), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n211), .B1(new_n277), .B2(new_n466), .ZN(new_n572));
  INV_X1    g0372(.A(G274), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n272), .A2(G45), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n298), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n344), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n566), .B(new_n578), .C1(G169), .C2(new_n577), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n316), .A2(new_n267), .A3(new_n495), .A4(G87), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n565), .A2(new_n555), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(G200), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(new_n376), .C2(new_n576), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n458), .A2(G270), .A3(new_n298), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT85), .B1(new_n585), .B2(new_n469), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n333), .B(new_n587), .C1(new_n213), .C2(G1698), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n295), .C1(G303), .C2(new_n333), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n458), .A2(G270), .A3(new_n298), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT85), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n297), .C2(new_n468), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT86), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT86), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n586), .A2(new_n595), .A3(new_n589), .A4(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n514), .A2(new_n230), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n259), .B2(G97), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n267), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n230), .A2(G116), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  NOR4_X1   g0405(.A1(new_n267), .A2(new_n600), .A3(new_n605), .A4(new_n602), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n316), .A2(G116), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n496), .B2(new_n254), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n594), .A2(G190), .A3(new_n596), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n598), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(G169), .B1(new_n607), .B2(new_n610), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n586), .A2(G179), .A3(new_n589), .A4(new_n592), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n611), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n597), .A2(KEYINPUT21), .A3(new_n615), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n613), .A2(new_n618), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NOR4_X1   g0423(.A1(new_n454), .A2(new_n550), .A3(new_n584), .A4(new_n623), .ZN(G372));
  AOI21_X1  g0424(.A(KEYINPUT89), .B1(new_n576), .B2(new_n346), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n626), .B(G169), .C1(new_n571), .C2(new_n575), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n566), .B(new_n578), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n628), .A2(new_n583), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n628), .B2(new_n583), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n549), .B(new_n506), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT21), .B1(new_n597), .B2(new_n615), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n617), .B(new_n614), .C1(new_n594), .C2(new_n596), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n633), .A2(new_n634), .A3(new_n620), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n501), .A2(new_n476), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  INV_X1    g0438(.A(new_n548), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n638), .B(new_n639), .C1(new_n630), .C2(new_n631), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n584), .B2(new_n548), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n628), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n453), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n381), .B(KEYINPUT10), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n449), .A2(new_n450), .ZN(new_n645));
  INV_X1    g0445(.A(new_n314), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n357), .A2(new_n284), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n348), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n445), .A2(new_n446), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n644), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n389), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n643), .A2(new_n653), .ZN(G369));
  NOR2_X1   g0454(.A1(new_n278), .A2(G20), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT27), .B1(new_n277), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n272), .A2(new_n658), .A3(new_n655), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n657), .A2(new_n659), .A3(G213), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G343), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT91), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n502), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n502), .A2(new_n506), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n501), .A2(new_n662), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT92), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n635), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n663), .A2(new_n611), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n623), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n636), .A2(new_n662), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n635), .A2(new_n662), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n668), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n221), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n305), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n529), .A2(new_n210), .A3(new_n254), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(G1), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n232), .A2(G50), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n683), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n689));
  XNOR2_X1  g0489(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  INV_X1    g0491(.A(new_n632), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n618), .A2(new_n502), .A3(new_n621), .A4(new_n622), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT26), .B(new_n639), .C1(new_n630), .C2(new_n631), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n638), .B1(new_n584), .B2(new_n548), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT95), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n698), .B(new_n638), .C1(new_n584), .C2(new_n548), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n694), .A2(new_n628), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n691), .B1(new_n701), .B2(new_n663), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n618), .A2(new_n621), .A3(new_n622), .A4(new_n636), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n692), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n640), .A2(new_n628), .A3(new_n641), .ZN(new_n705));
  AOI211_X1 g0505(.A(KEYINPUT29), .B(new_n662), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n516), .A2(new_n518), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n471), .A2(new_n464), .A3(new_n474), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n577), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n709), .B1(new_n712), .B2(new_n619), .ZN(new_n713));
  AND4_X1   g0513(.A1(G179), .A2(new_n586), .A3(new_n589), .A4(new_n592), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n516), .A2(new_n518), .A3(new_n576), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n344), .B(new_n576), .C1(new_n516), .C2(new_n518), .ZN(new_n718));
  AOI211_X1 g0518(.A(new_n503), .B(new_n718), .C1(new_n594), .C2(new_n596), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n662), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(KEYINPUT31), .B(new_n662), .C1(new_n717), .C2(new_n719), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(KEYINPUT94), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT94), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n725), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n623), .ZN(new_n728));
  INV_X1    g0528(.A(new_n550), .ZN(new_n729));
  INV_X1    g0529(.A(new_n584), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n663), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n708), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n707), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT96), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n690), .B1(new_n735), .B2(G1), .ZN(G364));
  NOR2_X1   g0536(.A1(new_n673), .A2(G330), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n268), .B1(new_n655), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n682), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n674), .A3(new_n742), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n346), .A2(KEYINPUT99), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n346), .A2(KEYINPUT99), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(G20), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(new_n226), .A3(new_n228), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n251), .A2(G45), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n681), .A2(new_n333), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(G45), .C2(new_n687), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n333), .A2(G355), .A3(new_n221), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G116), .B2(new_n221), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT98), .Z(new_n759));
  AOI21_X1  g0559(.A(new_n753), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n230), .A2(new_n344), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n312), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n291), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n230), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n763), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n767), .A2(G322), .B1(new_n770), .B2(G283), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n376), .A2(G179), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n230), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n771), .B1(new_n772), .B2(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT101), .Z(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n765), .B(new_n777), .C1(G329), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n766), .A2(new_n312), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT100), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G326), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n762), .A2(new_n778), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n782), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT102), .Z(new_n789));
  INV_X1    g0589(.A(new_n767), .ZN(new_n790));
  INV_X1    g0590(.A(G58), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n769), .A2(new_n335), .ZN(new_n793));
  INV_X1    g0593(.A(new_n779), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(KEYINPUT32), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n793), .B(new_n796), .C1(G50), .C2(new_n783), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n333), .B1(new_n764), .B2(new_n280), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(G77), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n776), .A2(new_n210), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n774), .A2(new_n212), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(KEYINPUT32), .C2(new_n795), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n797), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n789), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n742), .B1(new_n805), .B2(new_n748), .ZN(new_n806));
  INV_X1    g0606(.A(new_n751), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n673), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n743), .B1(new_n760), .B2(new_n808), .ZN(G396));
  NAND4_X1  g0609(.A1(new_n332), .A2(new_n345), .A3(new_n347), .A4(new_n662), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT105), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n348), .A2(KEYINPUT104), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT104), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n332), .A2(new_n345), .A3(new_n813), .A4(new_n347), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n332), .A2(new_n662), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n392), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n811), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n663), .B(new_n818), .C1(new_n637), .C2(new_n642), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT106), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n662), .B1(new_n704), .B2(new_n705), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT106), .B1(new_n822), .B2(new_n818), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n821), .A2(new_n823), .B1(new_n822), .B2(new_n818), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(new_n732), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n742), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n780), .A2(new_n827), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n333), .B1(new_n776), .B2(new_n202), .C1(new_n774), .C2(new_n791), .ZN(new_n829));
  INV_X1    g0629(.A(new_n764), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n783), .A2(G137), .B1(new_n830), .B2(G150), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n832), .B2(new_n790), .C1(new_n410), .C2(new_n787), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n828), .B(new_n829), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .C1(new_n280), .C2(new_n769), .ZN(new_n836));
  INV_X1    g0636(.A(G283), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n764), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n770), .A2(G87), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n790), .B2(new_n772), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G303), .B2(new_n783), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n291), .B1(new_n787), .B2(new_n254), .ZN(new_n842));
  INV_X1    g0642(.A(new_n776), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n802), .C1(G107), .C2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(new_n786), .C2(new_n780), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n836), .B1(new_n838), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n747), .A2(new_n750), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT103), .Z(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n846), .A2(new_n748), .B1(new_n250), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n741), .C1(new_n818), .C2(new_n750), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n826), .A2(new_n851), .ZN(G384));
  INV_X1    g0652(.A(KEYINPUT40), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n284), .A2(new_n662), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n648), .A2(new_n646), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n284), .B(new_n662), .C1(new_n357), .C2(new_n314), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n857), .A2(new_n818), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n623), .A2(new_n550), .A3(new_n584), .A4(new_n662), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n722), .A2(new_n723), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n434), .A2(new_n422), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n660), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n424), .A2(new_n863), .A3(new_n439), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n863), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n442), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n863), .B1(new_n650), .B2(new_n645), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n435), .A2(new_n402), .B1(new_n862), .B2(new_n660), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT37), .B1(new_n873), .B2(new_n439), .ZN(new_n874));
  NOR4_X1   g0674(.A1(new_n871), .A2(new_n872), .A3(new_n874), .A4(new_n866), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n853), .B1(new_n861), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n866), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n869), .C1(new_n451), .C2(new_n863), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n872), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n731), .A2(new_n722), .A3(new_n723), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n883), .A4(new_n858), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT110), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n453), .A2(new_n883), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(G330), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n815), .A2(new_n663), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT108), .Z(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n821), .B2(new_n823), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n882), .A3(new_n857), .ZN(new_n894));
  INV_X1    g0694(.A(new_n660), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n651), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT109), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n898), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n900), .B(new_n901), .C1(new_n870), .C2(new_n875), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n648), .A2(new_n662), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT109), .A4(KEYINPUT39), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n894), .A2(new_n896), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n453), .B1(new_n702), .B2(new_n706), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n653), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n906), .B(new_n908), .Z(new_n909));
  XNOR2_X1  g0709(.A(new_n889), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n272), .B2(new_n655), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n403), .A2(G77), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n687), .A2(new_n912), .B1(G50), .B2(new_n280), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n278), .A3(new_n277), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n254), .B1(new_n531), .B2(KEYINPUT35), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(new_n231), .C1(KEYINPUT35), .C2(new_n531), .ZN(new_n916));
  XOR2_X1   g0716(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n911), .A2(new_n914), .A3(new_n918), .ZN(G367));
  NOR2_X1   g0719(.A1(new_n769), .A2(new_n250), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n774), .A2(new_n280), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n920), .B(new_n921), .C1(G150), .C2(new_n767), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n333), .B1(new_n787), .B2(new_n202), .C1(new_n410), .C2(new_n764), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G137), .B2(new_n794), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n784), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n925), .B1(new_n791), .B2(new_n776), .C1(new_n832), .C2(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n790), .A2(new_n775), .B1(new_n212), .B2(new_n769), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n774), .A2(new_n335), .ZN(new_n929));
  INV_X1    g0729(.A(G317), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n291), .B1(new_n779), .B2(new_n930), .C1(new_n772), .C2(new_n764), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT46), .B1(new_n843), .B2(G116), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n837), .B2(new_n787), .C1(new_n786), .C2(new_n926), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n843), .A2(KEYINPUT46), .A3(G116), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT115), .Z(new_n936));
  OAI21_X1  g0736(.A(new_n927), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT47), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n742), .B1(new_n938), .B2(new_n748), .ZN(new_n939));
  INV_X1    g0739(.A(new_n755), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n752), .B1(new_n221), .B2(new_n328), .C1(new_n240), .C2(new_n940), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n630), .A2(new_n631), .B1(new_n581), .B2(new_n663), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n663), .A2(new_n628), .A3(new_n581), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n939), .B(new_n941), .C1(new_n807), .C2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n739), .B(KEYINPUT114), .Z(new_n946));
  INV_X1    g0746(.A(new_n679), .ZN(new_n947));
  INV_X1    g0747(.A(new_n545), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n549), .B1(new_n948), .B2(new_n663), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n639), .A2(new_n662), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT44), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT44), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n679), .A2(new_n954), .A3(new_n951), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT45), .B1(new_n679), .B2(new_n951), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n953), .A2(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n675), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n676), .B1(new_n956), .B2(new_n957), .C1(new_n953), .C2(new_n955), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n678), .B1(new_n673), .B2(G330), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n668), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n735), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n735), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n682), .B(KEYINPUT41), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n946), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n676), .A2(KEYINPUT112), .A3(new_n952), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT112), .B1(new_n676), .B2(new_n952), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n944), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n967), .A2(new_n970), .A3(new_n971), .A4(new_n968), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n668), .A2(new_n678), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n976), .A2(KEYINPUT42), .A3(new_n952), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n548), .B1(new_n949), .B2(new_n502), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n663), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT42), .B1(new_n976), .B2(new_n952), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT113), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n973), .A2(new_n983), .A3(new_n981), .A4(new_n974), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n945), .B1(new_n966), .B2(new_n987), .ZN(G387));
  OR2_X1    g0788(.A1(new_n735), .A2(new_n962), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n735), .A2(new_n962), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n682), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n962), .A2(new_n946), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n317), .A2(KEYINPUT50), .A3(G50), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n684), .B1(G68), .B2(G77), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT50), .B1(new_n317), .B2(G50), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n466), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n940), .B1(new_n245), .B2(G45), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n685), .A2(new_n681), .A3(new_n291), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n681), .A2(new_n335), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n753), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n784), .A2(G322), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n767), .A2(G317), .B1(new_n799), .B2(G303), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n786), .C2(new_n764), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n837), .B2(new_n774), .C1(new_n772), .C2(new_n776), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n794), .A2(G326), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n333), .B1(new_n770), .B2(G116), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n764), .A2(new_n317), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n776), .A2(new_n250), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G97), .B2(new_n770), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n202), .B2(new_n790), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G159), .B2(new_n783), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n774), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n552), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n333), .B1(new_n779), .B2(new_n360), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G68), .B2(new_n799), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1012), .B1(new_n1013), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1001), .B1(new_n1023), .B2(new_n748), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n741), .C1(new_n668), .C2(new_n807), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT116), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n991), .A2(new_n992), .A3(new_n1026), .ZN(G393));
  NAND2_X1  g0827(.A1(new_n959), .A2(new_n960), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n990), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n682), .A3(new_n963), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n959), .A2(new_n960), .A3(new_n946), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G150), .A2(new_n783), .B1(new_n767), .B2(G159), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT51), .Z(new_n1033));
  NOR2_X1   g0833(.A1(new_n774), .A2(new_n250), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n787), .A2(new_n317), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n333), .B1(new_n779), .B2(new_n832), .C1(new_n202), .C2(new_n764), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G68), .C2(new_n843), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1033), .A2(new_n839), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G311), .A2(new_n767), .B1(new_n783), .B2(G317), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT52), .Z(new_n1041));
  OAI22_X1  g0841(.A1(new_n774), .A2(new_n254), .B1(new_n787), .B2(new_n772), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n333), .B1(new_n794), .B2(G322), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n335), .B2(new_n769), .C1(new_n837), .C2(new_n776), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT118), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1041), .B(new_n1046), .C1(new_n1045), .C2(new_n1044), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n764), .A2(new_n775), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1039), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT119), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n742), .B1(new_n1050), .B2(new_n748), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n752), .B1(new_n212), .B2(new_n221), .C1(new_n255), .C2(new_n940), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT117), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n807), .C2(new_n951), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1030), .A2(new_n1031), .A3(new_n1054), .ZN(G390));
  NAND3_X1  g0855(.A1(new_n453), .A2(new_n883), .A3(G330), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT120), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n907), .A2(new_n1056), .A3(new_n1057), .A4(new_n653), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n907), .A2(new_n1056), .A3(new_n653), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT120), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n819), .A2(new_n820), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n822), .A2(KEYINPUT106), .A3(new_n818), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n891), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n727), .A2(new_n731), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(G330), .A3(new_n818), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n857), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n883), .A2(G330), .A3(new_n858), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(G330), .A3(new_n818), .A4(new_n857), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n700), .A2(new_n628), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n662), .B1(new_n1071), .B2(new_n694), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1072), .A2(new_n818), .B1(new_n663), .B2(new_n815), .ZN(new_n1073));
  OAI211_X1 g0873(.A(G330), .B(new_n818), .C1(new_n859), .C2(new_n860), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1066), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1058), .B(new_n1060), .C1(new_n1069), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(KEYINPUT121), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n857), .B1(new_n732), .B2(new_n818), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n883), .A2(G330), .A3(new_n858), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n893), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT121), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n882), .B1(new_n648), .B2(new_n662), .C1(new_n1073), .C2(new_n1066), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n903), .B1(new_n893), .B2(new_n857), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n902), .A2(new_n904), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1068), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1070), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1087), .B(new_n1092), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n683), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n946), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n333), .B1(new_n1100), .B2(new_n787), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G159), .A2(new_n1018), .B1(new_n783), .B2(G128), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n202), .B2(new_n769), .C1(new_n827), .C2(new_n790), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G125), .C2(new_n781), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n830), .A2(G137), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n776), .A2(new_n360), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT122), .Z(new_n1109));
  NOR2_X1   g0909(.A1(new_n787), .A2(new_n212), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1035), .B1(new_n254), .B2(new_n790), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G283), .B2(new_n783), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n291), .B1(new_n764), .B2(new_n335), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n801), .B(new_n1113), .C1(G68), .C2(new_n770), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(new_n772), .C2(new_n780), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n742), .B1(new_n1116), .B2(new_n748), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n318), .B2(new_n848), .C1(new_n1089), .C2(new_n750), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1097), .A2(new_n1098), .A3(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(KEYINPUT57), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT124), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1060), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1058), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1060), .A2(KEYINPUT124), .A3(new_n1058), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n877), .A2(G330), .A3(new_n884), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n906), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT56), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n644), .A2(new_n389), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n364), .A2(new_n660), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT55), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1131), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1138), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(KEYINPUT56), .A3(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1128), .A2(new_n894), .A3(new_n896), .A4(new_n905), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1130), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1130), .B2(new_n1144), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1120), .B1(new_n1127), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n882), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1128), .B1(new_n1151), .B2(new_n896), .ZN(new_n1152));
  AND4_X1   g0952(.A1(new_n896), .A2(new_n1128), .A3(new_n894), .A4(new_n905), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1142), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1130), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1078), .A2(new_n1085), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(KEYINPUT57), .C1(new_n1157), .C2(new_n1126), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1148), .A2(new_n682), .A3(new_n1158), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n305), .C2(new_n333), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n333), .B(new_n305), .C1(new_n830), .C2(G97), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n328), .B2(new_n787), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n921), .B(new_n1162), .C1(G283), .C2(new_n781), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n769), .A2(new_n791), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1164), .B(new_n1014), .C1(G116), .C2(new_n783), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(new_n335), .C2(new_n790), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT123), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1167), .A2(KEYINPUT58), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(KEYINPUT58), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n767), .A2(G128), .B1(new_n799), .B2(G137), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n783), .A2(G125), .B1(new_n843), .B2(new_n1099), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1018), .A2(G150), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n830), .A2(G132), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n794), .A2(G124), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n770), .C2(G159), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AND4_X1   g0979(.A1(new_n1160), .A2(new_n1168), .A3(new_n1169), .A4(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1180), .A2(new_n747), .B1(G50), .B2(new_n848), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n742), .B(new_n1181), .C1(new_n1143), .C2(new_n749), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1156), .B2(new_n946), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1159), .A2(new_n1183), .ZN(G375));
  NAND2_X1  g0984(.A1(new_n1083), .A2(new_n946), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n781), .A2(G128), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n333), .B1(new_n787), .B2(new_n360), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1164), .B(new_n1187), .C1(G132), .C2(new_n783), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n830), .A2(new_n1099), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n774), .A2(new_n202), .B1(new_n776), .B2(new_n410), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G137), .B2(new_n767), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n333), .B1(new_n830), .B2(G116), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n799), .A2(G107), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1019), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n920), .B(new_n1195), .C1(G294), .C2(new_n783), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n781), .A2(G303), .B1(G97), .B2(new_n843), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT125), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(KEYINPUT125), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n790), .A2(new_n837), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1192), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1202), .A2(new_n748), .B1(new_n280), .B2(new_n849), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n741), .B(new_n1203), .C1(new_n857), .C2(new_n750), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1185), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1081), .B(new_n1082), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1078), .A2(new_n1207), .A3(new_n1085), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n965), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(G381));
  NOR2_X1   g1010(.A1(G375), .A2(G378), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1030), .A2(new_n1031), .A3(new_n1054), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1209), .B1(new_n963), .B2(new_n735), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n986), .B(new_n985), .C1(new_n1214), .C2(new_n946), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1215), .A3(new_n945), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1212), .A3(new_n1217), .ZN(G407));
  INV_X1    g1018(.A(G343), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G407), .A2(G213), .A3(new_n1220), .ZN(G409));
  OAI211_X1 g1021(.A(new_n1156), .B(new_n965), .C1(new_n1157), .C2(new_n1126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1183), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1098), .A2(new_n1118), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT126), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1159), .A2(G378), .A3(new_n1183), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT126), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1223), .A2(new_n1229), .A3(new_n1225), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1219), .A2(G213), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1208), .A2(KEYINPUT60), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1083), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT60), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n682), .A3(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(G384), .A3(new_n1206), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n682), .B1(new_n1234), .B2(KEYINPUT60), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(KEYINPUT60), .B2(new_n1208), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n826), .B(new_n851), .C1(new_n1239), .C2(new_n1205), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1231), .A2(new_n1232), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT62), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1219), .A2(G213), .A3(G2897), .ZN(new_n1245));
  AOI211_X1 g1045(.A(KEYINPUT127), .B(new_n1245), .C1(new_n1237), .C2(new_n1240), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT127), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1245), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1241), .B2(new_n1247), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1246), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1231), .A2(new_n1255), .A3(new_n1232), .A4(new_n1242), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1244), .A2(new_n1253), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(G390), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(G393), .B(G396), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1258), .A2(new_n1216), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1258), .B2(new_n1216), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1232), .A4(new_n1242), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1265), .A2(new_n1262), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1243), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1266), .B(new_n1254), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(G375), .A2(new_n1225), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1228), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1262), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1262), .A2(new_n1273), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1241), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1276), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1242), .A3(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(G402));
endmodule


