//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(new_n212), .B2(new_n211), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT67), .B(G77), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G58), .A2(G232), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n220), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G223), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(new_n221), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n247), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n214), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(G274), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(new_n263), .C1(G41), .C2(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n253), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n254), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G200), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT10), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G150), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT71), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT8), .ZN(new_n280));
  OR2_X1    g0080(.A1(KEYINPUT8), .A2(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n278), .B1(new_n282), .B2(new_n284), .C1(new_n283), .C2(new_n204), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n213), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n202), .ZN(new_n291));
  INV_X1    g0091(.A(new_n287), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G1), .B2(new_n283), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n293), .B2(new_n202), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT9), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n272), .B1(new_n297), .B2(new_n271), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n276), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n295), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n298), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(new_n275), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT16), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n201), .B1(new_n279), .B2(G68), .ZN(new_n306));
  INV_X1    g0106(.A(G159), .ZN(new_n307));
  INV_X1    g0107(.A(new_n277), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n306), .A2(new_n283), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G68), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n283), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT7), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n311), .A2(KEYINPUT7), .A3(new_n283), .A4(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n310), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n305), .B1(new_n309), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n321), .B2(new_n283), .ZN(new_n322));
  INV_X1    g0122(.A(new_n316), .ZN(new_n323));
  OAI21_X1  g0123(.A(G68), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n308), .A2(new_n307), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT71), .A2(G58), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT71), .A2(G58), .ZN(new_n327));
  OAI21_X1  g0127(.A(G68), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n216), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(G20), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n318), .A2(new_n287), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n287), .B1(new_n263), .B2(G20), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n282), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n289), .B2(new_n282), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G223), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n248), .ZN(new_n339));
  INV_X1    g0139(.A(G226), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n341), .C1(new_n319), .C2(new_n320), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G87), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT69), .B(G45), .ZN(new_n345));
  AOI21_X1  g0145(.A(G1), .B1(new_n345), .B2(new_n259), .ZN(new_n346));
  INV_X1    g0146(.A(G274), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n253), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n344), .A2(new_n253), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n266), .A2(new_n268), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(G232), .A3(new_n262), .ZN(new_n351));
  AOI21_X1  g0151(.A(G169), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n344), .A2(new_n253), .ZN(new_n354));
  AND4_X1   g0154(.A1(new_n353), .A2(new_n354), .A3(new_n264), .A4(new_n351), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT77), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NOR2_X1   g0157(.A1(G223), .A2(G1698), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n340), .B2(G1698), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n247), .B1(G33), .B2(G87), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n264), .B1(new_n360), .B2(new_n262), .ZN(new_n361));
  INV_X1    g0161(.A(new_n351), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n349), .A2(new_n353), .A3(new_n351), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n337), .A2(new_n356), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT18), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT17), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n361), .B2(new_n362), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n349), .A2(new_n297), .A3(new_n351), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(new_n332), .A3(new_n336), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n369), .B1(new_n374), .B2(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n324), .A2(new_n330), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n292), .B1(new_n376), .B2(new_n305), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n335), .B1(new_n377), .B2(new_n331), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT17), .A4(new_n373), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n337), .A2(new_n356), .A3(new_n381), .A4(new_n366), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n368), .A2(new_n375), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n271), .A2(G179), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n385), .B(new_n295), .C1(new_n357), .C2(new_n271), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n293), .A2(new_n205), .B1(new_n221), .B2(new_n289), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT8), .B(G58), .Z(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n277), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n283), .B2(new_n251), .C1(new_n284), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n287), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G232), .A2(G1698), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n248), .A2(G238), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n247), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n253), .C1(G107), .C2(new_n247), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n269), .A2(G244), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n264), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n393), .B(new_n400), .C1(new_n357), .C2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(G200), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(KEYINPUT72), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n399), .A2(new_n297), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n403), .B2(KEYINPUT72), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n304), .A2(new_n384), .A3(new_n387), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n269), .A2(G238), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n340), .A2(new_n248), .ZN(new_n410));
  INV_X1    g0210(.A(G232), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n412), .C1(new_n319), .C2(new_n320), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT74), .B1(new_n415), .B2(new_n253), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT74), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n417), .B(new_n262), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n409), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n346), .A2(new_n348), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT13), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(G226), .A2(G1698), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n411), .B2(G1698), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n247), .B1(G33), .B2(G97), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n417), .B1(new_n427), .B2(new_n262), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n415), .A2(KEYINPUT74), .A3(new_n253), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n420), .A2(new_n422), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n409), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(KEYINPUT13), .C1(new_n419), .C2(new_n423), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(G169), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n434), .A2(new_n439), .A3(G169), .A4(new_n436), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n424), .A2(G179), .A3(new_n433), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT12), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n290), .B2(new_n310), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n293), .A2(new_n310), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT11), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n308), .A2(new_n202), .B1(new_n283), .B2(G68), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n284), .A2(new_n205), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n287), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n447), .B2(new_n450), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n433), .A2(G190), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n454), .B2(new_n424), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n434), .A2(G200), .A3(new_n436), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n408), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n283), .C1(G33), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT87), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n287), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n287), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT20), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n263), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n289), .A2(new_n472), .A3(new_n213), .A4(new_n286), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n289), .A2(new_n464), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n470), .A2(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n247), .A2(G264), .A3(G1698), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n247), .A2(G257), .A3(new_n248), .ZN(new_n478));
  INV_X1    g0278(.A(G303), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(new_n247), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n253), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n255), .A2(G1), .ZN(new_n482));
  AND2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G270), .A3(new_n262), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n262), .A2(new_n487), .A3(G274), .A4(new_n482), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT86), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT86), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n481), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT21), .A3(G169), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n481), .B(G179), .C1(new_n490), .C2(new_n489), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n476), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT90), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n283), .B2(G107), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT23), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n496), .B(new_n499), .C1(new_n283), .C2(G107), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n283), .A2(KEYINPUT89), .A3(G87), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n311), .B2(new_n312), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(KEYINPUT22), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n283), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n283), .A2(KEYINPUT89), .A3(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n247), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n504), .A2(new_n511), .A3(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n509), .A2(new_n510), .B1(new_n498), .B2(new_n500), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n503), .A2(KEYINPUT22), .B1(new_n283), .B2(new_n506), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n287), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n292), .A2(KEYINPUT80), .A3(new_n289), .A4(new_n472), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n473), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n520), .A3(G107), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n289), .A2(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT25), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n526));
  OAI211_X1 g0326(.A(G250), .B(new_n248), .C1(new_n319), .C2(new_n320), .ZN(new_n527));
  AND2_X1   g0327(.A1(KEYINPUT91), .A2(G294), .ZN(new_n528));
  NOR2_X1   g0328(.A1(KEYINPUT91), .A2(G294), .ZN(new_n529));
  OAI21_X1  g0329(.A(G33), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n253), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n487), .A2(new_n482), .B1(new_n214), .B2(new_n261), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT92), .B1(new_n533), .B2(G264), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n485), .A2(KEYINPUT92), .A3(G264), .A4(new_n262), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n488), .B(new_n532), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n517), .A2(new_n525), .B1(new_n357), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n537), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n353), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT88), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n491), .A2(G169), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(new_n476), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n474), .A2(new_n475), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n287), .A2(new_n465), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n287), .A2(new_n463), .A3(new_n465), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT20), .B1(new_n551), .B2(new_n462), .ZN(new_n552));
  INV_X1    g0352(.A(new_n471), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(G169), .A3(new_n491), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n542), .B1(new_n555), .B2(new_n543), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n495), .B(new_n541), .C1(new_n546), .C2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n491), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n554), .B1(new_n559), .B2(G190), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n370), .B2(new_n559), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n283), .B1(new_n414), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT84), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n565), .B(new_n283), .C1(new_n414), .C2(new_n562), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G87), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT85), .ZN(new_n568));
  INV_X1    g0368(.A(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n564), .B(new_n566), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n283), .A2(G33), .A3(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n562), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n310), .A2(G20), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n321), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n292), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n518), .A2(new_n520), .A3(G87), .ZN(new_n581));
  INV_X1    g0381(.A(new_n391), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(new_n289), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G238), .B(new_n248), .C1(new_n319), .C2(new_n320), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n247), .A2(KEYINPUT83), .A3(G238), .A4(new_n248), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n505), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n262), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n348), .A2(new_n482), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n263), .A2(G45), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n595), .A2(G250), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n262), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(G200), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n348), .A2(new_n482), .B1(new_n262), .B2(new_n596), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n591), .B1(new_n587), .B2(new_n588), .ZN(new_n601));
  OAI211_X1 g0401(.A(G190), .B(new_n600), .C1(new_n601), .C2(new_n262), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n584), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n518), .A2(new_n520), .A3(new_n582), .ZN(new_n604));
  INV_X1    g0404(.A(new_n583), .ZN(new_n605));
  INV_X1    g0405(.A(G87), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n461), .A3(new_n569), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n570), .B1(KEYINPUT84), .B2(new_n563), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n578), .B1(new_n609), .B2(new_n566), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n604), .B(new_n605), .C1(new_n610), .C2(new_n292), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n353), .B(new_n600), .C1(new_n601), .C2(new_n262), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n589), .A2(new_n592), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n598), .B1(new_n613), .B2(new_n253), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n611), .B(new_n612), .C1(new_n614), .C2(G169), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n603), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n537), .A2(new_n370), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n485), .A2(G264), .A3(new_n262), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT92), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n535), .B1(new_n253), .B2(new_n531), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n297), .A3(new_n488), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT24), .B1(new_n504), .B2(new_n511), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n514), .A2(new_n515), .A3(new_n513), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n524), .B1(new_n626), .B2(new_n287), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n623), .A2(new_n627), .A3(KEYINPUT93), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT93), .B1(new_n623), .B2(new_n627), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n616), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n485), .A2(G257), .A3(new_n262), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n488), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT81), .ZN(new_n634));
  OAI211_X1 g0434(.A(G244), .B(new_n248), .C1(new_n319), .C2(new_n320), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT4), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n460), .ZN(new_n638));
  NAND2_X1  g0438(.A1(G250), .A2(G1698), .ZN(new_n639));
  NAND2_X1  g0439(.A1(KEYINPUT4), .A2(G244), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(G1698), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n247), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n634), .B1(new_n643), .B2(new_n253), .ZN(new_n644));
  AOI211_X1 g0444(.A(KEYINPUT81), .B(new_n262), .C1(new_n637), .C2(new_n642), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n633), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT82), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT82), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n648), .B(new_n633), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(G200), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n262), .B1(new_n637), .B2(new_n642), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(new_n632), .A3(new_n297), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n290), .A2(G97), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n518), .A2(new_n520), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(G97), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n569), .A2(KEYINPUT6), .A3(G97), .ZN(new_n656));
  XNOR2_X1  g0456(.A(G97), .B(G107), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT6), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n659), .A2(new_n283), .B1(new_n205), .B2(new_n308), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n569), .B1(new_n315), .B2(new_n316), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n287), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT79), .ZN(new_n663));
  OAI21_X1  g0463(.A(G107), .B1(new_n322), .B2(new_n323), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n308), .A2(new_n205), .ZN(new_n665));
  AND2_X1   g0465(.A1(G97), .A2(G107), .ZN(new_n666));
  NOR2_X1   g0466(.A1(G97), .A2(G107), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n658), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n569), .A2(KEYINPUT6), .A3(G97), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n670), .B2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT79), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n287), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n652), .B(new_n655), .C1(new_n663), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n650), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n655), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n673), .B1(new_n672), .B2(new_n287), .ZN(new_n678));
  AOI211_X1 g0478(.A(KEYINPUT79), .B(new_n292), .C1(new_n664), .C2(new_n671), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n353), .B(new_n633), .C1(new_n644), .C2(new_n645), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n651), .A2(new_n632), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G169), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n676), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n630), .A2(new_n686), .ZN(new_n687));
  AND4_X1   g0487(.A1(new_n459), .A2(new_n558), .A3(new_n561), .A4(new_n687), .ZN(G372));
  NAND2_X1  g0488(.A1(new_n375), .A2(new_n380), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n457), .A2(new_n401), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n453), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n368), .A2(new_n382), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n304), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT96), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(new_n694), .A3(new_n387), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n693), .B2(new_n387), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT94), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n630), .B2(new_n686), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n603), .A2(new_n615), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n623), .A2(new_n627), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n623), .A2(new_n627), .A3(KEYINPUT93), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n663), .A2(new_n674), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n683), .B1(new_n706), .B2(new_n677), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n650), .A2(new_n675), .B1(new_n707), .B2(new_n681), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(KEYINPUT94), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n557), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n543), .B1(new_n544), .B2(new_n476), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT88), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n545), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(KEYINPUT95), .A3(new_n495), .A4(new_n541), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n699), .A2(new_n709), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n615), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n616), .A2(KEYINPUT26), .A3(new_n681), .A4(new_n707), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT26), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n685), .B2(new_n700), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n717), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n459), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n697), .A2(new_n723), .ZN(G369));
  NAND3_X1  g0524(.A1(new_n263), .A2(new_n283), .A3(G13), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G213), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G343), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n541), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT97), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n541), .B1(new_n627), .B2(new_n731), .C1(new_n628), .C2(new_n629), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n494), .B1(new_n713), .B2(new_n545), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n730), .ZN(new_n738));
  INV_X1    g0538(.A(new_n541), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n736), .A2(new_n738), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n737), .A2(new_n561), .B1(new_n554), .B2(new_n730), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n476), .A2(new_n731), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n736), .A3(G330), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT98), .ZN(G399));
  INV_X1    g0546(.A(new_n210), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G41), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n571), .A2(new_n572), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n464), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(G1), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n217), .B2(new_n749), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n557), .A2(new_n705), .A3(new_n708), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n721), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(KEYINPUT29), .A3(new_n731), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n730), .B1(new_n716), .B2(new_n721), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(KEYINPUT29), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n687), .A2(new_n558), .A3(new_n561), .A4(new_n731), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n539), .A2(new_n614), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(new_n353), .A3(new_n491), .A4(new_n646), .ZN(new_n763));
  INV_X1    g0563(.A(new_n493), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n651), .A2(new_n632), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n764), .A2(new_n767), .A3(KEYINPUT30), .A4(new_n614), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT30), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n614), .A2(new_n621), .A3(new_n682), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n493), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n763), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n730), .ZN(new_n773));
  AOI21_X1  g0573(.A(KEYINPUT31), .B1(new_n772), .B2(new_n730), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n761), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n760), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n755), .B1(new_n778), .B2(G1), .ZN(G364));
  NAND2_X1  g0579(.A1(new_n743), .A2(G330), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n283), .A2(G13), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n263), .B1(new_n781), .B2(G45), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n749), .A2(KEYINPUT99), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT99), .ZN(new_n784));
  INV_X1    g0584(.A(new_n782), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n748), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n743), .A2(G330), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n213), .B1(G20), .B2(new_n357), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n283), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n606), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n794), .B1(G97), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n283), .A2(new_n353), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G190), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n321), .B1(new_n802), .B2(new_n221), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n792), .A2(new_n800), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT32), .B1(new_n804), .B2(new_n307), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n798), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n799), .A2(G190), .A3(new_n370), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT101), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n279), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n799), .A2(G200), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G190), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n792), .A2(new_n297), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n812), .A2(G68), .B1(new_n814), .B2(G107), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n804), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n811), .A2(new_n297), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G50), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n806), .A2(new_n810), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  INV_X1    g0620(.A(G329), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n801), .A2(new_n820), .B1(new_n804), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n807), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n247), .B(new_n822), .C1(G322), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n817), .A2(G326), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n812), .A2(new_n826), .B1(new_n814), .B2(G283), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n528), .A2(new_n529), .ZN(new_n828));
  INV_X1    g0628(.A(new_n793), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n797), .A2(new_n828), .B1(new_n829), .B2(G303), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n824), .A2(new_n825), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n791), .B1(new_n819), .B2(new_n831), .ZN(new_n832));
  OR3_X1    g0632(.A1(KEYINPUT100), .A2(G13), .A3(G33), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT100), .B1(G13), .B2(G33), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n790), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n210), .A2(G355), .A3(new_n247), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n747), .A2(new_n247), .ZN(new_n840));
  INV_X1    g0640(.A(new_n345), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n217), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n245), .A2(new_n255), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n839), .B1(G116), .B2(new_n210), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n787), .B(new_n832), .C1(new_n838), .C2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT102), .ZN(new_n846));
  INV_X1    g0646(.A(new_n837), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n743), .A2(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n788), .A2(new_n789), .B1(new_n846), .B2(new_n848), .ZN(G396));
  INV_X1    g0649(.A(new_n787), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n404), .A2(new_n406), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n393), .A2(new_n731), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n401), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n401), .A2(new_n731), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n759), .B(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n850), .B1(new_n858), .B2(new_n777), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n777), .B2(new_n858), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n836), .A2(new_n791), .ZN(new_n861));
  INV_X1    g0661(.A(new_n804), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n247), .B1(new_n862), .B2(G311), .ZN(new_n863));
  INV_X1    g0663(.A(G294), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n464), .B2(new_n801), .C1(new_n864), .C2(new_n807), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n817), .A2(G303), .B1(new_n829), .B2(G107), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n606), .B2(new_n813), .ZN(new_n867));
  INV_X1    g0667(.A(new_n812), .ZN(new_n868));
  INV_X1    g0668(.A(G283), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n868), .A2(new_n869), .B1(new_n461), .B2(new_n796), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n865), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n813), .A2(new_n310), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  INV_X1    g0673(.A(new_n279), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n247), .B1(new_n804), .B2(new_n873), .C1(new_n796), .C2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n872), .B(new_n875), .C1(G50), .C2(new_n829), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT103), .Z(new_n877));
  INV_X1    g0677(.A(KEYINPUT34), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n817), .A2(G137), .B1(new_n802), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G150), .ZN(new_n880));
  INV_X1    g0680(.A(G143), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n880), .B2(new_n868), .C1(new_n808), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n882), .A2(new_n878), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n871), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n850), .B1(G77), .B2(new_n861), .C1(new_n885), .C2(new_n791), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT104), .Z(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n836), .B2(new_n857), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n860), .A2(new_n888), .ZN(G384));
  NAND4_X1  g0689(.A1(new_n328), .A2(G50), .A3(new_n216), .A4(new_n221), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n202), .A2(G68), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n263), .B(G13), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT105), .Z(new_n893));
  INV_X1    g0693(.A(KEYINPUT36), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n464), .B(new_n215), .C1(new_n670), .C2(KEYINPUT35), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(KEYINPUT35), .B2(new_n670), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n442), .A2(new_n452), .A3(new_n731), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT106), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n324), .B2(new_n330), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n292), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n318), .A2(KEYINPUT106), .A3(new_n287), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n331), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n728), .B1(new_n905), .B2(new_n336), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n383), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n336), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n909), .A2(new_n912), .B1(new_n378), .B2(new_n373), .ZN(new_n913));
  INV_X1    g0713(.A(new_n906), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT107), .B1(new_n912), .B2(new_n337), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n337), .A2(new_n356), .A3(KEYINPUT107), .A4(new_n366), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n374), .B(new_n908), .C1(new_n378), .C2(new_n728), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n907), .B(KEYINPUT38), .C1(new_n915), .C2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT108), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n367), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n374), .B1(new_n378), .B2(new_n728), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT107), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n367), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n917), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n929), .B2(new_n919), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n378), .A2(new_n728), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n383), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT39), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n383), .B2(new_n906), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(KEYINPUT108), .C1(new_n915), .C2(new_n920), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n923), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n907), .B1(new_n915), .B2(new_n920), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n934), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n941), .B2(new_n921), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT109), .ZN(new_n944));
  INV_X1    g0744(.A(new_n942), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n923), .A2(new_n935), .A3(new_n937), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n900), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n855), .B1(new_n759), .B2(new_n857), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n452), .A2(new_n730), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n453), .A2(new_n457), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n457), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n452), .B(new_n730), .C1(new_n442), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n941), .A2(new_n921), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n956), .A2(new_n957), .B1(new_n692), .B2(new_n728), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n948), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n459), .B(new_n758), .C1(new_n759), .C2(KEYINPUT29), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n697), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n856), .B1(new_n761), .B2(new_n775), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n963), .A2(new_n954), .A3(KEYINPUT40), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n933), .A2(new_n934), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n923), .A2(new_n937), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n954), .A3(new_n963), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT110), .B(KEYINPUT40), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n459), .A3(new_n776), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(G330), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n971), .B1(new_n459), .B2(new_n776), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n962), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n263), .B2(new_n781), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n962), .A2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n898), .B1(new_n977), .B2(new_n978), .ZN(G367));
  NAND2_X1  g0779(.A1(new_n680), .A2(new_n730), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n708), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n707), .A2(new_n681), .A3(new_n730), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n736), .A2(new_n738), .A3(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n739), .A2(new_n676), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n730), .B1(new_n986), .B2(new_n685), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(KEYINPUT42), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n584), .A2(new_n731), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n616), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n615), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n985), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n983), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n744), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n748), .B(KEYINPUT41), .Z(new_n1001));
  NAND3_X1  g0801(.A1(new_n740), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n740), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n998), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(KEYINPUT44), .A3(new_n998), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n740), .B2(new_n983), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1002), .A2(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT111), .B1(new_n1009), .B2(new_n744), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1005), .A2(new_n1002), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT111), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n744), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n736), .B(new_n738), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT112), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n780), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1017), .B(new_n1019), .Z(new_n1020));
  INV_X1    g0820(.A(new_n778), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1009), .A2(new_n744), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1010), .A2(new_n1016), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1001), .B1(new_n1024), .B2(new_n778), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1000), .B1(new_n1025), .B2(new_n785), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n840), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(new_n237), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n838), .B1(new_n210), .B2(new_n391), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n850), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G137), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n801), .A2(new_n202), .B1(new_n804), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n321), .B(new_n1032), .C1(G150), .C2(new_n823), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n797), .A2(G68), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n221), .A2(new_n814), .B1(new_n829), .B2(new_n279), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n812), .A2(G159), .B1(new_n817), .B2(G143), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(KEYINPUT114), .B(G317), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n321), .B1(new_n804), .B2(new_n1038), .C1(new_n869), .C2(new_n801), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n809), .B2(G303), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n814), .A2(G97), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n812), .A2(new_n828), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G107), .A2(new_n797), .B1(new_n817), .B2(G311), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT113), .B1(new_n793), .B2(new_n464), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT46), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1037), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT47), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1030), .B1(new_n1048), .B2(new_n790), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n847), .B2(new_n992), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1026), .A2(new_n1050), .ZN(G387));
  NAND3_X1  g0851(.A1(new_n751), .A2(new_n210), .A3(new_n247), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(G107), .B2(new_n210), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n389), .A2(new_n202), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT50), .Z(new_n1056));
  AOI21_X1  g0856(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n752), .A3(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n840), .C1(new_n234), .C2(new_n345), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n787), .B1(new_n1060), .B2(new_n838), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n797), .A2(new_n582), .B1(new_n829), .B2(new_n221), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n817), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1041), .C1(new_n307), .C2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n823), .A2(G50), .B1(new_n862), .B2(G150), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n321), .B1(new_n802), .B2(G68), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n282), .C2(new_n868), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n813), .A2(new_n464), .ZN(new_n1069));
  INV_X1    g0869(.A(G326), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n321), .B1(new_n804), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n817), .A2(G322), .B1(new_n802), .B2(G303), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n820), .B2(new_n868), .C1(new_n808), .C2(new_n1038), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n797), .A2(G283), .B1(new_n829), .B2(new_n828), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1069), .B(new_n1071), .C1(new_n1079), .C2(KEYINPUT49), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1079), .A2(KEYINPUT49), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1068), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1061), .B1(new_n1082), .B2(new_n791), .C1(new_n736), .C2(new_n847), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n748), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1083), .B1(new_n782), .B2(new_n1020), .C1(new_n1084), .C2(new_n1085), .ZN(G393));
  NOR2_X1   g0886(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1009), .A2(new_n744), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n782), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n998), .A2(new_n837), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT116), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n838), .B1(new_n461), .B2(new_n210), .C1(new_n1027), .C2(new_n241), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n796), .A2(new_n205), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n389), .B2(new_n802), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n202), .B2(new_n868), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT118), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1063), .A2(new_n880), .B1(new_n307), .B2(new_n807), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n321), .B1(new_n862), .B2(G143), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n310), .B2(new_n793), .C1(new_n606), .C2(new_n813), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G317), .A2(new_n817), .B1(new_n823), .B2(G311), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  OAI22_X1  g0905(.A1(new_n868), .A2(new_n479), .B1(new_n569), .B2(new_n813), .ZN(new_n1106));
  INV_X1    g0906(.A(G322), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n321), .B1(new_n804), .B2(new_n1107), .C1(new_n864), .C2(new_n801), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n796), .A2(new_n464), .B1(new_n793), .B2(new_n869), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1096), .A2(new_n1103), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n850), .B(new_n1092), .C1(new_n1111), .C2(new_n791), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1091), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1089), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n748), .B1(new_n1115), .B2(new_n1022), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1024), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n954), .B1(new_n963), .B2(G330), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n730), .B(new_n853), .C1(new_n756), .C2(new_n721), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n855), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n963), .A2(new_n954), .A3(G330), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT120), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G330), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1127), .B(new_n856), .C1(new_n761), .C2(new_n775), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(KEYINPUT120), .A3(new_n954), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1119), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1130), .B2(new_n949), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n459), .A2(G330), .A3(new_n776), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n960), .B(new_n1132), .C1(new_n695), .C2(new_n696), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n899), .B1(new_n949), .B2(new_n955), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT109), .B1(new_n938), .B2(new_n942), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n945), .A2(new_n944), .A3(new_n946), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n954), .B1(new_n1121), .B2(new_n855), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n966), .A3(new_n899), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT119), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n966), .A3(KEYINPUT119), .A4(new_n899), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1139), .A2(new_n1145), .A3(new_n1123), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT120), .B1(new_n1128), .B2(new_n954), .ZN(new_n1147));
  AND4_X1   g0947(.A1(KEYINPUT120), .A2(new_n963), .A3(G330), .A4(new_n954), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1135), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1149), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1120), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n949), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1133), .B1(new_n1157), .B2(new_n1124), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1139), .A2(new_n1145), .A3(new_n1123), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1152), .A2(new_n1160), .A3(new_n748), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT124), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n282), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n850), .B1(new_n1163), .B2(new_n861), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n817), .A2(G283), .B1(new_n802), .B2(G97), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n569), .B2(new_n868), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT122), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n321), .B1(new_n804), .B2(new_n864), .C1(new_n807), .C2(new_n464), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1168), .A2(new_n794), .A3(new_n1093), .A4(new_n872), .ZN(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n807), .A2(new_n873), .B1(new_n804), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n321), .B(new_n1171), .C1(new_n802), .C2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n793), .A2(new_n880), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT53), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n812), .A2(G137), .B1(new_n814), .B2(G50), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G159), .A2(new_n797), .B1(new_n817), .B2(G128), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1167), .A2(new_n1169), .B1(new_n1179), .B2(KEYINPUT121), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(KEYINPUT121), .B2(new_n1179), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1164), .B1(new_n1181), .B2(new_n790), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT123), .Z(new_n1183));
  NOR2_X1   g0983(.A1(new_n943), .A2(new_n947), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n835), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n785), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1161), .A2(new_n1162), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1162), .B1(new_n1161), .B2(new_n1187), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(G378));
  NAND3_X1  g0990(.A1(new_n967), .A2(new_n970), .A3(G330), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n304), .A2(new_n387), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n295), .A2(new_n728), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n304), .B(new_n387), .C1(new_n295), .C2(new_n728), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(G330), .A3(new_n970), .A4(new_n967), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n959), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n948), .A3(new_n958), .A4(new_n1204), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1202), .A2(new_n835), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n850), .B1(G50), .B2(new_n861), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n321), .B2(new_n259), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n868), .A2(new_n461), .B1(new_n1063), .B2(new_n464), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n279), .B2(new_n814), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G41), .B(new_n247), .C1(new_n802), .C2(new_n582), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n823), .A2(G107), .B1(new_n862), .B2(G283), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n797), .A2(G68), .B1(new_n829), .B2(new_n221), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1212), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n807), .A2(new_n1221), .B1(new_n801), .B2(new_n1031), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n812), .A2(G132), .B1(new_n829), .B2(new_n1173), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1170), .B2(new_n1063), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G150), .C2(new_n797), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n814), .A2(G159), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n862), .C2(G124), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1220), .B1(new_n1219), .B2(new_n1218), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1210), .B1(new_n1232), .B2(new_n790), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1208), .A2(new_n785), .B1(new_n1209), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1133), .B1(new_n1186), .B2(new_n1131), .ZN(new_n1235));
  AND4_X1   g1035(.A1(new_n948), .A2(new_n1203), .A3(new_n958), .A4(new_n1204), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1203), .A2(new_n1204), .B1(new_n948), .B2(new_n958), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n748), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1160), .A2(new_n1134), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1208), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1234), .B1(new_n1239), .B2(new_n1241), .ZN(G375));
  NAND2_X1  g1042(.A1(new_n955), .A2(new_n835), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n809), .A2(G137), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n796), .A2(new_n202), .B1(new_n793), .B2(new_n307), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G132), .B2(new_n817), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n247), .B1(new_n801), .B2(new_n880), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G128), .B2(new_n862), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n812), .A2(new_n1173), .B1(new_n814), .B2(new_n279), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n813), .A2(new_n205), .B1(new_n793), .B2(new_n461), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G116), .B2(new_n812), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n247), .B1(new_n862), .B2(G303), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n823), .A2(G283), .B1(new_n802), .B2(G107), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n582), .A2(new_n797), .B1(new_n817), .B2(G294), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n791), .B1(new_n1250), .B2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n861), .A2(G68), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1257), .A2(new_n787), .A3(new_n1258), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1131), .A2(new_n785), .B1(new_n1243), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1001), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1135), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1262), .B2(new_n1263), .ZN(G381));
  INV_X1    g1064(.A(G390), .ZN(new_n1265));
  INV_X1    g1065(.A(G384), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G387), .A2(new_n1267), .A3(G381), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1161), .A2(new_n1187), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G375), .B(KEYINPUT125), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(G407));
  INV_X1    g1072(.A(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n729), .A2(G213), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT126), .Z(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(new_n1271), .C2(new_n1276), .ZN(G409));
  NAND3_X1  g1077(.A1(new_n1240), .A2(new_n1261), .A3(new_n1208), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1234), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1273), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1270), .A2(KEYINPUT124), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1161), .A2(new_n1187), .A3(new_n1162), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1280), .B1(new_n1283), .B2(G375), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1275), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1157), .A2(KEYINPUT60), .A3(new_n1133), .A4(new_n1124), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1287), .A2(new_n748), .A3(new_n1288), .A4(new_n1135), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1260), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1266), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(G384), .A3(new_n1260), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1284), .A2(new_n1285), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1275), .A2(G2897), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1291), .A2(new_n1300), .A3(new_n1292), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1300), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1298), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1270), .B1(new_n1234), .B2(new_n1278), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1234), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1240), .A2(new_n1208), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT57), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n749), .B1(new_n1240), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1305), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1304), .B1(new_n1311), .B2(G378), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1299), .B(new_n1303), .C1(new_n1312), .C2(new_n1275), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1284), .A2(new_n1314), .A3(new_n1285), .A4(new_n1294), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1296), .A2(new_n1297), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G393), .A2(G396), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1268), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1026), .A2(new_n1050), .A3(G390), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G390), .B1(new_n1026), .B2(new_n1050), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1318), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G387), .A2(new_n1265), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1323), .A2(new_n1268), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1312), .A2(new_n1275), .A3(new_n1293), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(new_n1327), .B2(KEYINPUT63), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1302), .A2(new_n1298), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1284), .A2(new_n1285), .B1(new_n1329), .B2(new_n1301), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1330), .B2(new_n1299), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1295), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1328), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1326), .A2(new_n1334), .ZN(G405));
  NOR2_X1   g1135(.A1(new_n1283), .A2(G375), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(new_n1273), .B2(G375), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1293), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1337), .A2(new_n1293), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1325), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  OR2_X1    g1141(.A1(new_n1337), .A2(new_n1293), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1325), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(new_n1343), .A3(new_n1338), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1344), .ZN(G402));
endmodule


