//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1263, new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n452), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n452), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n460), .A2(KEYINPUT68), .B1(G567), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT69), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n470), .A2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n472), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n465), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n465), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n484), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT71), .Z(G162));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(KEYINPUT72), .B2(G114), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT72), .A2(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n495), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(KEYINPUT73), .C1(new_n493), .C2(new_n492), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n502), .B(new_n503), .C1(new_n472), .C2(new_n471), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n466), .B2(new_n502), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n499), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n510), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(new_n520), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n511), .A2(new_n512), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n522), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n513), .A2(new_n522), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT74), .B(G90), .Z(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(new_n540), .B1(G52), .B2(new_n520), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n515), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n520), .A2(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n523), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n532), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(new_n539), .B2(G91), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n520), .A2(new_n559), .A3(G53), .ZN(new_n560));
  INV_X1    g135(.A(new_n519), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT6), .A2(G651), .ZN(new_n562));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n565), .B1(new_n560), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n558), .B1(new_n566), .B2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  OR2_X1    g144(.A1(new_n516), .A2(new_n525), .ZN(G303));
  NAND2_X1  g145(.A1(new_n539), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n520), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n532), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n539), .B2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n520), .A2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n520), .A2(new_n581), .A3(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(G305));
  XNOR2_X1  g159(.A(KEYINPUT77), .B(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n529), .A2(new_n585), .B1(new_n523), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n515), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n520), .A2(G54), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n515), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n523), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(G868), .B2(new_n600), .ZN(G284));
  OAI21_X1  g176(.A(new_n592), .B1(G868), .B2(new_n600), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n466), .A2(new_n475), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT13), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n483), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n485), .A2(G123), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n620));
  INV_X1    g195(.A(G111), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n620), .B2(new_n619), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n616), .A2(new_n625), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT79), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(KEYINPUT79), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(G401));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n659), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT81), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n671), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(G6), .ZN(new_n688));
  INV_X1    g263(.A(G305), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n682), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n682), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n682), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n694), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n687), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n483), .A2(G131), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n485), .A2(G119), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n708));
  NOR2_X1   g283(.A1(G95), .A2(G2105), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT83), .ZN(new_n710));
  INV_X1    g285(.A(G107), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n474), .B1(new_n711), .B2(G2105), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n708), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n710), .A2(new_n708), .A3(new_n712), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n706), .B(new_n707), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G25), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n682), .A2(G24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n590), .B2(new_n682), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1986), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n704), .A2(new_n705), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT36), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G32), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n483), .A2(G141), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n485), .A2(G129), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT26), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(G105), .B2(new_n475), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(KEYINPUT91), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(KEYINPUT91), .B2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G160), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n728), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT94), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n549), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G16), .B2(G19), .ZN(new_n754));
  INV_X1    g329(.A(G1341), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n682), .A2(G5), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G301), .B2(G16), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n682), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n682), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G1966), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n741), .A2(new_n752), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n728), .A2(G33), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n483), .A2(G139), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  INV_X1    g342(.A(G127), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n479), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(KEYINPUT88), .A3(G2105), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n766), .A2(new_n772), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n765), .B1(new_n777), .B2(new_n728), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT89), .Z(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G2072), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n754), .A2(new_n755), .B1(new_n624), .B2(new_n728), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n749), .A2(new_n750), .B1(new_n758), .B2(new_n756), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n682), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n600), .B2(new_n682), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G1348), .ZN(new_n786));
  INV_X1    g361(.A(G2078), .ZN(new_n787));
  NAND2_X1  g362(.A1(G164), .A2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G27), .B2(G29), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n787), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT31), .B(G11), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n728), .B1(new_n793), .B2(G28), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(G28), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n792), .B(new_n798), .C1(new_n761), .C2(G1966), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G1348), .B2(new_n785), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n783), .A2(new_n790), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n764), .A2(new_n780), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n682), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n604), .B2(new_n682), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT95), .B(G1956), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n728), .A2(G26), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT28), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n485), .A2(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n479), .A2(new_n480), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n812));
  OAI211_X1 g387(.A(G140), .B(new_n465), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(G116), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n810), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n809), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2067), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n805), .A2(new_n806), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n802), .A2(new_n807), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n728), .A2(G35), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G162), .B2(new_n728), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT29), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2090), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n779), .A2(G2072), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT92), .Z(new_n828));
  NOR3_X1   g403(.A1(new_n822), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n727), .A2(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n520), .A2(G55), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n513), .A2(new_n522), .A3(G93), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n513), .A2(G67), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n515), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n832), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n835), .A2(new_n839), .A3(KEYINPUT97), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n599), .A2(new_n598), .ZN(new_n847));
  INV_X1    g422(.A(new_n595), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n607), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI221_X1 g427(.A(new_n546), .B1(new_n523), .B2(new_n547), .C1(new_n544), .C2(new_n515), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n841), .B2(new_n842), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n549), .A2(new_n840), .A3(new_n836), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n852), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n844), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n816), .B1(new_n485), .B2(G128), .ZN(new_n863));
  NAND3_X1  g438(.A1(G164), .A2(new_n813), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(G126), .A2(G2105), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n479), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n502), .B1(new_n471), .B2(new_n472), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT4), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n868), .B2(new_n504), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n496), .A2(new_n498), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n818), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n864), .A2(new_n872), .A3(new_n776), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n776), .B1(new_n864), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n737), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G164), .B1(new_n813), .B2(new_n863), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n818), .A2(new_n871), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n777), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n864), .A2(new_n872), .A3(new_n776), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n738), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n485), .A2(G130), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n485), .A2(KEYINPUT98), .A3(G130), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  INV_X1    g462(.A(G118), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n483), .A2(G142), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n715), .A2(new_n614), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n715), .A2(new_n614), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n881), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT99), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT100), .B1(new_n881), .B2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(new_n900), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n880), .A4(new_n875), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n881), .A2(new_n907), .A3(new_n900), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n902), .A2(new_n903), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n624), .B(new_n748), .ZN(new_n910));
  XNOR2_X1  g485(.A(G162), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n901), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n881), .A2(KEYINPUT101), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n875), .A2(new_n880), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n917), .A3(new_n904), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT102), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n915), .A2(new_n920), .A3(new_n917), .A4(new_n904), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n914), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n913), .B1(new_n922), .B2(KEYINPUT103), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n924));
  AOI211_X1 g499(.A(new_n924), .B(new_n914), .C1(new_n919), .C2(new_n921), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n862), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n919), .A2(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n927), .B2(new_n914), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(KEYINPUT103), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(KEYINPUT40), .A3(new_n929), .A4(new_n913), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n926), .A2(new_n930), .ZN(G395));
  NAND2_X1  g506(.A1(G303), .A2(new_n697), .ZN(new_n932));
  NAND2_X1  g507(.A1(G166), .A2(G288), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G305), .A2(new_n590), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(G305), .A2(new_n590), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n689), .A2(G290), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n939), .A2(new_n933), .A3(new_n932), .A4(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n942));
  NOR2_X1   g517(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n609), .B(KEYINPUT104), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(new_n856), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n600), .B(new_n558), .C1(new_n567), .C2(new_n566), .ZN(new_n947));
  NAND2_X1  g522(.A1(G299), .A2(new_n849), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT41), .B1(new_n947), .B2(new_n948), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n950), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n944), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G868), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g532(.A(new_n956), .B1(G868), .B2(new_n843), .ZN(G331));
  OAI211_X1 g533(.A(new_n538), .B(new_n541), .C1(new_n535), .C2(new_n531), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n539), .A2(new_n540), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n520), .A2(G52), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n537), .A2(new_n515), .ZN(new_n963));
  OAI21_X1  g538(.A(G168), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n854), .A2(new_n855), .A3(new_n959), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n959), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n836), .A2(new_n840), .A3(new_n832), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT97), .B1(new_n835), .B2(new_n839), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n549), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n853), .A2(new_n839), .A3(new_n835), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n949), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n966), .A2(new_n969), .A3(new_n970), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n854), .A2(new_n855), .B1(new_n959), .B2(new_n964), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n953), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n941), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n949), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n965), .A4(new_n971), .ZN(new_n981));
  INV_X1    g556(.A(new_n949), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n973), .B2(new_n974), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n941), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n941), .A3(new_n983), .ZN(new_n988));
  INV_X1    g563(.A(G37), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n976), .B2(new_n941), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(KEYINPUT106), .A3(new_n985), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  MUX2_X1   g570(.A(new_n987), .B(new_n994), .S(new_n995), .Z(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT107), .B1(new_n994), .B2(new_n995), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n984), .B2(new_n985), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n991), .B(new_n941), .C1(new_n981), .C2(new_n983), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n977), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n977), .A2(new_n995), .A3(new_n986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT44), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT108), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n1010), .B(new_n1007), .C1(new_n999), .C2(new_n1004), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n998), .B1(new_n1009), .B2(new_n1011), .ZN(G397));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n499), .B2(new_n507), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT69), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n468), .B(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G125), .ZN(new_n1020));
  INV_X1    g595(.A(new_n472), .ZN(new_n1021));
  NAND2_X1  g596(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(G2105), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(G40), .A3(new_n476), .A4(new_n473), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1013), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G40), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n470), .A2(new_n1027), .A3(new_n477), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1015), .A2(KEYINPUT109), .A3(new_n1016), .A4(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1996), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(KEYINPUT110), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(G1996), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n737), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G2067), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n818), .B(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n737), .A2(G1996), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n715), .B(new_n719), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1034), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n590), .B(G1986), .Z(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1030), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1016), .A2(G1384), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n499), .B2(new_n507), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n869), .B2(new_n870), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1049), .B(new_n1028), .C1(KEYINPUT45), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n686), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(G2090), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n1014), .C1(new_n499), .C2(new_n507), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1028), .A4(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1057), .A3(KEYINPUT111), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G303), .A2(G8), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1028), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1064));
  AOI211_X1 g639(.A(KEYINPUT50), .B(G1384), .C1(new_n869), .C2(new_n870), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(G2090), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1025), .B1(new_n871), .B2(new_n1048), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1971), .B1(new_n1017), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1059), .A2(KEYINPUT112), .A3(new_n1062), .A4(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(G8), .A3(new_n1058), .A4(new_n1062), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1050), .B2(new_n1028), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n697), .A2(G1976), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(G288), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G305), .A2(G1981), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n1085));
  INV_X1    g660(.A(G1981), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n578), .A2(new_n583), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G305), .A2(KEYINPUT113), .A3(G1981), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1075), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1082), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1070), .A2(new_n1073), .A3(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1078), .B(new_n697), .C1(new_n1093), .C2(new_n1090), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1087), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1075), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1966), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1051), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1053), .A2(new_n750), .A3(new_n1028), .A4(new_n1056), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(G168), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  AND2_X1   g680(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(G8), .A3(G286), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1105), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT62), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1051), .B2(G2078), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT53), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1113), .B(new_n1116), .C1(new_n1051), .C2(G2078), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n756), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT51), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1109), .A4(new_n1107), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1112), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1091), .A2(new_n1075), .A3(new_n1092), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1064), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1050), .A2(new_n1130), .A3(new_n1055), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1054), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1074), .B1(new_n1134), .B2(new_n1052), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1128), .B(new_n1129), .C1(new_n1062), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1073), .B2(new_n1070), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1100), .B1(new_n1126), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1050), .A2(new_n1038), .A3(new_n1028), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n600), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n560), .A2(new_n564), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n558), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n560), .B2(new_n564), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT57), .B(new_n558), .C1(new_n566), .C2(new_n567), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1956), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT56), .B(G2072), .Z(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1017), .A2(new_n1067), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1153), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1144), .A2(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1154), .B2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1166), .A2(new_n1053), .A3(new_n1028), .A4(new_n1133), .ZN(new_n1167));
  INV_X1    g742(.A(G1956), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1165), .A2(new_n1169), .A3(KEYINPUT117), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1160), .A2(new_n1161), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT61), .B1(new_n1172), .B2(new_n1159), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1159), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT58), .B(G1341), .Z(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1015), .B2(new_n1025), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1051), .B2(G1996), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT119), .B1(new_n1179), .B2(new_n549), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(KEYINPUT119), .A3(new_n549), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(KEYINPUT59), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT59), .ZN(new_n1183));
  AOI211_X1 g758(.A(KEYINPUT119), .B(new_n1183), .C1(new_n1179), .C2(new_n549), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1176), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1173), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1142), .ZN(new_n1187));
  OAI211_X1 g762(.A(KEYINPUT120), .B(new_n600), .C1(new_n1187), .C2(KEYINPUT60), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n849), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1187), .A2(KEYINPUT60), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1188), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1171), .B1(new_n1186), .B2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1197), .A2(new_n1198), .A3(G301), .A4(new_n1117), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT124), .B1(new_n1119), .B2(G171), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1199), .A2(KEYINPUT54), .A3(new_n1200), .A4(new_n1120), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1123), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1202));
  XNOR2_X1  g777(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1119), .A2(G171), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1203), .B1(new_n1121), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1137), .A2(new_n1201), .A3(new_n1202), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1138), .B1(new_n1196), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1134), .A2(new_n1052), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1062), .B1(new_n1209), .B2(G8), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1211), .B(new_n1080), .C1(new_n1093), .C2(new_n1090), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g788(.A(new_n1074), .B(G286), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1208), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT63), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1108), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1212), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1062), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1069), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1058), .A2(G8), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g800(.A(KEYINPUT115), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT115), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1208), .A2(new_n1227), .A3(new_n1224), .A4(new_n1220), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1217), .A2(new_n1226), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1047), .B1(new_n1207), .B2(new_n1229), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1034), .A2(G1986), .A3(G290), .ZN(new_n1231));
  XNOR2_X1  g806(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1231), .B(new_n1232), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1233), .A2(new_n1037), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT47), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT46), .ZN(new_n1236));
  AOI21_X1  g811(.A(KEYINPUT110), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1237));
  NOR3_X1   g812(.A1(new_n1034), .A2(new_n1033), .A3(G1996), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1032), .A2(KEYINPUT46), .A3(new_n1035), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1034), .B1(new_n738), .B2(new_n1039), .ZN(new_n1242));
  INV_X1    g817(.A(new_n1242), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1235), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  AOI211_X1 g819(.A(KEYINPUT47), .B(new_n1242), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1234), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n716), .A2(new_n719), .ZN(new_n1247));
  XNOR2_X1  g822(.A(new_n1247), .B(KEYINPUT125), .ZN(new_n1248));
  NOR3_X1   g823(.A1(new_n1036), .A2(new_n1041), .A3(new_n1248), .ZN(new_n1249));
  NOR2_X1   g824(.A1(new_n818), .A2(G2067), .ZN(new_n1250));
  OAI21_X1  g825(.A(new_n1030), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g826(.A(new_n1251), .ZN(new_n1252));
  OAI21_X1  g827(.A(KEYINPUT127), .B1(new_n1246), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1254), .A2(KEYINPUT47), .ZN(new_n1255));
  NAND3_X1  g830(.A1(new_n1241), .A2(new_n1235), .A3(new_n1243), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1258));
  NAND4_X1  g833(.A1(new_n1257), .A2(new_n1258), .A3(new_n1251), .A4(new_n1234), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1253), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g835(.A1(new_n1230), .A2(new_n1260), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g836(.A1(new_n928), .A2(new_n929), .A3(new_n913), .ZN(new_n1263));
  OR2_X1    g837(.A1(new_n463), .A2(G227), .ZN(new_n1264));
  NOR3_X1   g838(.A1(G229), .A2(G401), .A3(new_n1264), .ZN(new_n1265));
  AND3_X1   g839(.A1(new_n1263), .A2(new_n996), .A3(new_n1265), .ZN(G308));
  NAND3_X1  g840(.A1(new_n1263), .A2(new_n996), .A3(new_n1265), .ZN(G225));
endmodule


