//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  AOI21_X1  g004(.A(G131), .B1(new_n189), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT65), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT64), .B1(new_n203), .B2(G146), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n200), .B(new_n202), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G143), .B2(new_n199), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n210), .B2(new_n201), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n192), .A2(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n189), .A2(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  AND4_X1   g030(.A1(new_n187), .A2(new_n198), .A3(new_n212), .A4(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n196), .A2(new_n197), .B1(G131), .B2(new_n215), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n187), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g034(.A(G116), .B(G119), .Z(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT2), .B(G113), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n221), .A2(new_n226), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n190), .A2(new_n193), .A3(new_n214), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n198), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n199), .B2(G143), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(G143), .B2(new_n199), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n236), .A2(new_n238), .B1(new_n240), .B2(new_n208), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n229), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n220), .A2(KEYINPUT28), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n232), .A2(new_n241), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n198), .A2(new_n212), .A3(new_n216), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n229), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n246), .B2(new_n229), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n218), .A2(new_n187), .A3(new_n212), .ZN(new_n260));
  INV_X1    g074(.A(new_n229), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n259), .A2(new_n244), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n255), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n246), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n259), .A2(new_n244), .A3(KEYINPUT30), .A4(new_n260), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n229), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT31), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT68), .B1(new_n262), .B2(new_n255), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT31), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n258), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  NOR2_X1   g092(.A1(G472), .A2(G902), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n257), .B1(new_n283), .B2(new_n275), .ZN(new_n284));
  INV_X1    g098(.A(new_n279), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT32), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n256), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n259), .A2(new_n260), .A3(new_n244), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n220), .A2(new_n242), .B1(new_n290), .B2(new_n229), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n249), .B(new_n289), .C1(new_n291), .C2(new_n248), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n243), .A2(new_n255), .A3(new_n249), .A4(new_n247), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n288), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n255), .B1(new_n271), .B2(new_n262), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n292), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n300), .A3(G472), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n287), .A2(new_n302), .A3(KEYINPUT70), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT70), .B1(new_n287), .B2(new_n302), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT16), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G125), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(G146), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n307), .A2(KEYINPUT72), .A3(G146), .A4(new_n310), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G128), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(G128), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n316), .B(new_n318), .C1(new_n319), .C2(KEYINPUT23), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n201), .A2(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT24), .B(G110), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n321), .A2(new_n325), .B1(new_n199), .B2(new_n306), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G953), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(G221), .A3(G234), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT73), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT22), .B(G137), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n332), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n323), .A2(new_n324), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n307), .A2(new_n310), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n199), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n338), .B2(new_n311), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n320), .A2(G110), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT71), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n327), .B(new_n335), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT74), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n342), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n349), .A2(new_n339), .B1(new_n315), .B2(new_n326), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n343), .B(new_n293), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n347), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n293), .A4(new_n343), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(new_n293), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n343), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  OAI21_X1  g180(.A(G221), .B1(new_n366), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n375), .B2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n374), .A3(KEYINPUT3), .A4(G104), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n372), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n371), .B1(new_n375), .B2(new_n370), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n210), .A2(new_n201), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n206), .B1(new_n236), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n372), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n369), .A2(G107), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n388), .B2(new_n377), .ZN(new_n389));
  INV_X1    g203(.A(new_n378), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n370), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n376), .B2(new_n378), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n391), .B(KEYINPUT4), .C1(new_n393), .C2(new_n371), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n370), .B1(new_n389), .B2(new_n390), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n241), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n196), .A2(new_n197), .B1(G131), .B2(new_n230), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n381), .A2(KEYINPUT10), .A3(new_n212), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n386), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n328), .A2(G227), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n402), .B(new_n403), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n206), .B(new_n211), .C1(new_n379), .C2(new_n380), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n384), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n232), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n405), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n386), .A2(new_n398), .A3(new_n400), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT77), .A3(new_n232), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT77), .B1(new_n413), .B2(new_n232), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n401), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n404), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n419), .A2(G469), .A3(G902), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n232), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT77), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n405), .B1(new_n424), .B2(new_n414), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n404), .B(KEYINPUT75), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n411), .A2(new_n408), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n401), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n421), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n405), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n415), .B2(new_n416), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT12), .B1(new_n407), .B2(new_n232), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n410), .B(new_n399), .C1(new_n384), .C2(new_n406), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n401), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n426), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(KEYINPUT78), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n430), .A2(new_n437), .A3(new_n293), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G469), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n420), .B1(new_n439), .B2(KEYINPUT79), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n441), .A3(G469), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n368), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n446));
  OAI21_X1  g260(.A(G131), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n446), .ZN(new_n448));
  INV_X1    g262(.A(G131), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n444), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT17), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(KEYINPUT17), .B(G131), .C1(new_n445), .C2(new_n446), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n338), .A3(new_n311), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n369), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n306), .B(new_n199), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT18), .B(G131), .C1(new_n445), .C2(new_n446), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n444), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n456), .B1(new_n454), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n293), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G475), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n447), .A2(new_n450), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n306), .A2(KEYINPUT19), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n306), .A2(KEYINPUT19), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n199), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n467), .A2(new_n313), .A3(new_n314), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n461), .ZN(new_n472));
  INV_X1    g286(.A(new_n456), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n476));
  NOR2_X1   g290(.A1(G475), .A2(G902), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n466), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G122), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT92), .B1(new_n483), .B2(G116), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n485));
  INV_X1    g299(.A(G116), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(G122), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n488), .A2(KEYINPUT14), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n488), .A2(KEYINPUT14), .B1(G116), .B2(new_n483), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n374), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n483), .A2(G116), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n374), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT93), .B1(new_n201), .B2(G143), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT93), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n203), .A3(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n201), .A2(G143), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n189), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n189), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n493), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n374), .B1(new_n488), .B2(new_n492), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n497), .A2(new_n506), .B1(new_n201), .B2(G143), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT13), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n189), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n491), .A2(new_n502), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n366), .A2(new_n358), .A3(G953), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI221_X1 g327(.A(new_n511), .B1(new_n505), .B2(new_n509), .C1(new_n491), .C2(new_n502), .ZN(new_n514));
  AOI21_X1  g328(.A(G902), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G478), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n515), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n482), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n328), .A2(G952), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT21), .B(G898), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G214), .B1(G237), .B2(G902), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT80), .Z(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT81), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G125), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n206), .A2(new_n211), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT86), .B1(new_n241), .B2(new_n534), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT86), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n236), .A2(new_n238), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n240), .A2(new_n208), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n539), .B(G125), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n328), .A2(G224), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n543), .B(new_n544), .Z(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(G116), .A3(new_n317), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT84), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n546), .A2(new_n549), .A3(G116), .A4(new_n317), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(G113), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n546), .B1(new_n222), .B2(new_n225), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n381), .A2(new_n228), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G122), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n227), .A2(new_n228), .B1(new_n395), .B2(new_n396), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n557), .A2(KEYINPUT82), .A3(new_n394), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT82), .B1(new_n557), .B2(new_n394), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n555), .B(new_n556), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n556), .B(KEYINPUT85), .Z(new_n562));
  AOI22_X1  g376(.A1(new_n560), .A2(KEYINPUT6), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n561), .A2(KEYINPUT6), .A3(new_n562), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n545), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n394), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n557), .A2(KEYINPUT82), .A3(new_n394), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n568), .A2(new_n569), .B1(new_n554), .B2(new_n553), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n542), .A2(new_n538), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n571), .A2(new_n537), .B1(KEYINPUT90), .B2(new_n544), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n570), .A2(new_n556), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n544), .A2(KEYINPUT90), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n543), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n223), .A2(KEYINPUT5), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n551), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G113), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n547), .B2(KEYINPUT84), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT89), .B1(new_n584), .B2(new_n550), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n554), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n228), .B1(new_n551), .B2(new_n552), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n379), .B2(new_n380), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n556), .B(KEYINPUT8), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n576), .A2(new_n577), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n574), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n565), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n565), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n533), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT91), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n565), .A2(new_n592), .ZN(new_n598));
  INV_X1    g412(.A(new_n593), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n565), .A2(new_n592), .A3(new_n593), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n533), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n529), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n305), .A2(new_n365), .A3(new_n443), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  OAI21_X1  g421(.A(G472), .B1(new_n284), .B2(G902), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n285), .B2(new_n284), .ZN(new_n609));
  INV_X1    g423(.A(new_n365), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n443), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n531), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n527), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n512), .B2(KEYINPUT94), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n513), .A2(new_n514), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n513), .B2(new_n514), .ZN(new_n619));
  OAI21_X1  g433(.A(G478), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n516), .A2(new_n293), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n515), .B2(new_n516), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n481), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT95), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n612), .A2(new_n615), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n518), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n466), .A2(KEYINPUT96), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n475), .A2(new_n477), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT20), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n478), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n466), .A2(KEYINPUT96), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n630), .A2(new_n631), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n612), .A2(new_n615), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n354), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n357), .A2(new_n359), .B1(new_n363), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n609), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n605), .A2(new_n443), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  AOI21_X1  g461(.A(new_n278), .B1(new_n277), .B2(new_n279), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n300), .B1(new_n297), .B2(G472), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n297), .A2(new_n300), .A3(G472), .ZN(new_n651));
  OAI22_X1  g465(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT70), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT97), .B(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n523), .B1(new_n655), .B2(new_n525), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n636), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n643), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n602), .A2(new_n657), .A3(new_n613), .A4(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n287), .A2(new_n302), .A3(KEYINPUT70), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n654), .A2(new_n659), .A3(new_n443), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XOR2_X1   g476(.A(new_n656), .B(KEYINPUT39), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n443), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n602), .B(KEYINPUT38), .ZN(new_n667));
  INV_X1    g481(.A(G472), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n281), .B1(new_n255), .B2(new_n291), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n293), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n287), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n482), .A2(new_n531), .A3(new_n518), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n643), .A2(new_n667), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n665), .A2(new_n666), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  INV_X1    g491(.A(new_n656), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n481), .A2(new_n620), .A3(new_n622), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n643), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n602), .A2(new_n680), .A3(new_n613), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n305), .A2(new_n677), .A3(new_n443), .A4(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n654), .A2(new_n443), .A3(new_n660), .A4(new_n682), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT98), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT99), .B(G146), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G48));
  OR3_X1    g502(.A1(new_n419), .A2(G469), .A3(G902), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n419), .B2(G902), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n367), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n654), .A2(new_n660), .A3(new_n365), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n615), .A2(new_n626), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT41), .B(G113), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND2_X1  g511(.A1(new_n615), .A2(new_n637), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n486), .ZN(G18));
  NOR2_X1   g514(.A1(new_n529), .A2(new_n643), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n614), .A2(new_n691), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n654), .A2(new_n701), .A3(new_n660), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  NAND2_X1  g518(.A1(new_n602), .A2(new_n673), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n691), .A3(new_n527), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n249), .B1(new_n291), .B2(new_n248), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n283), .A2(new_n275), .B1(new_n707), .B2(new_n256), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT100), .B1(new_n708), .B2(new_n285), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n256), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n272), .B2(new_n276), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT100), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n279), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n709), .A2(new_n713), .A3(new_n608), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n706), .A2(new_n365), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NOR3_X1   g530(.A1(new_n614), .A2(new_n691), .A3(new_n679), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n709), .A2(new_n713), .A3(new_n608), .A4(new_n658), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  NAND2_X1  g537(.A1(new_n652), .A2(new_n365), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(G469), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n435), .A2(KEYINPUT102), .A3(new_n426), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT102), .B1(new_n435), .B2(new_n426), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n432), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n729), .B2(new_n293), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n367), .B1(new_n420), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n600), .A2(new_n601), .A3(new_n613), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n679), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n654), .A2(new_n733), .A3(new_n660), .A4(new_n365), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT103), .B1(new_n735), .B2(new_n736), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT104), .B(G131), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G33));
  NOR2_X1   g556(.A1(new_n731), .A2(new_n732), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n305), .A2(new_n365), .A3(new_n657), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT43), .B1(new_n482), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n482), .A2(new_n624), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n643), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n751), .B(new_n609), .C1(new_n750), .C2(new_n749), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT108), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n732), .B1(new_n752), .B2(new_n753), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  OAI21_X1  g572(.A(G469), .B1(new_n729), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n430), .A2(new_n437), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n726), .A2(new_n293), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n689), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n367), .A3(new_n663), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT105), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n757), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  NAND2_X1  g584(.A1(new_n766), .A2(new_n367), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n305), .A2(new_n365), .A3(new_n679), .A4(new_n732), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n309), .ZN(G42));
  AND2_X1   g590(.A1(new_n722), .A2(new_n661), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n705), .A2(new_n731), .A3(new_n656), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n643), .A3(new_n672), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n686), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n722), .A2(new_n661), .A3(new_n779), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n683), .B2(new_n685), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n781), .B1(new_n783), .B2(KEYINPUT52), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n703), .B(new_n715), .C1(new_n693), .C2(new_n694), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n699), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n605), .A2(new_n443), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n654), .A2(new_n660), .A3(new_n365), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n597), .A2(new_n604), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n519), .B1(new_n482), .B2(new_n624), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n527), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n443), .A2(new_n790), .A3(new_n611), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n645), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT111), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n606), .A2(new_n796), .A3(new_n645), .A4(new_n793), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n786), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n732), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n631), .A2(new_n634), .A3(new_n635), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n643), .A2(new_n800), .A3(new_n630), .A4(new_n656), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n305), .A2(new_n443), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n718), .B(new_n719), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n733), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n744), .A2(new_n802), .A3(KEYINPUT53), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n735), .A2(new_n736), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT103), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n737), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n805), .B1(new_n809), .B2(new_n734), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n784), .A2(new_n798), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n784), .A2(new_n798), .A3(KEYINPUT114), .A4(new_n810), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n744), .A2(new_n802), .A3(new_n804), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n740), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n786), .A2(new_n795), .A3(new_n797), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n722), .A2(new_n661), .A3(new_n779), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n819), .A2(new_n686), .A3(KEYINPUT52), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(new_n819), .B2(new_n686), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n686), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n819), .A2(new_n686), .A3(KEYINPUT52), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n818), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n813), .A2(new_n814), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n829), .A2(new_n830), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n818), .A2(new_n784), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n830), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n835), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n833), .B1(new_n840), .B2(new_n832), .ZN(new_n841));
  INV_X1    g655(.A(new_n672), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n691), .A2(new_n732), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n365), .A3(new_n523), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n626), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n520), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n749), .A2(new_n523), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT115), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n691), .A3(new_n732), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n725), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT48), .Z(new_n851));
  NAND2_X1  g665(.A1(new_n714), .A2(new_n365), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n846), .B(new_n851), .C1(new_n702), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n799), .ZN(new_n855));
  INV_X1    g669(.A(new_n773), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n689), .A2(new_n368), .A3(new_n690), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n667), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(new_n531), .A3(new_n859), .A4(new_n692), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT50), .Z(new_n861));
  NOR3_X1   g675(.A1(new_n844), .A2(new_n481), .A3(new_n624), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n849), .B2(new_n803), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(KEYINPUT51), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n863), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n857), .B(KEYINPUT116), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n855), .B1(new_n856), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI221_X1 g682(.A(new_n854), .B1(new_n858), .B2(new_n864), .C1(KEYINPUT51), .C2(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n841), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n610), .A2(new_n748), .A3(new_n368), .A4(new_n532), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT110), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n689), .A2(new_n690), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(KEYINPUT49), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n874), .B(new_n859), .C1(KEYINPUT49), .C2(new_n873), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n870), .B1(new_n672), .B2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n328), .A2(G952), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n831), .A2(new_n293), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n563), .A2(new_n564), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n545), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT117), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n878), .B(KEYINPUT118), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n599), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT56), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n877), .B(new_n885), .C1(new_n887), .C2(new_n890), .ZN(G51));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n761), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT121), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n831), .B(new_n832), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n762), .B(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n419), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(KEYINPUT120), .B2(new_n896), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n877), .B1(new_n893), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  INV_X1    g714(.A(new_n475), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n877), .ZN(G60));
  OR2_X1    g718(.A1(new_n618), .A2(new_n619), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n621), .B(KEYINPUT59), .Z(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n841), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n894), .A2(new_n906), .A3(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n877), .A3(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n813), .A2(new_n814), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n829), .A2(new_n830), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n642), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n361), .B1(new_n831), .B2(new_n912), .ZN(new_n917));
  INV_X1    g731(.A(new_n877), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT61), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(new_n918), .C1(new_n915), .C2(new_n362), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n916), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n917), .B2(new_n918), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT123), .B(new_n920), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n915), .B2(new_n362), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n922), .A3(new_n916), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT123), .B1(new_n929), .B2(new_n920), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n919), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT124), .B(new_n919), .C1(new_n926), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  NAND2_X1  g749(.A1(G224), .A2(G953), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n817), .A2(G953), .B1(new_n526), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n880), .B1(G898), .B2(new_n328), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT125), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n937), .B(new_n939), .ZN(G69));
  INV_X1    g754(.A(new_n775), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n769), .A2(new_n744), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n686), .A2(new_n777), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n768), .A2(new_n602), .A3(new_n673), .A4(new_n725), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n942), .A2(new_n740), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n328), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n328), .A2(G900), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT127), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n269), .A2(new_n270), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n468), .A2(new_n469), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G227), .A2(G900), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n952), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n791), .B(KEYINPUT126), .Z(new_n957));
  NOR4_X1   g771(.A1(new_n788), .A2(new_n664), .A3(new_n957), .A4(new_n732), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n958), .B(new_n775), .C1(new_n757), .C2(new_n768), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n943), .A2(new_n675), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n956), .B1(new_n964), .B2(G953), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n953), .A2(new_n955), .A3(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(G953), .B(new_n954), .C1(new_n949), .C2(new_n956), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n945), .B2(new_n817), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n256), .A3(new_n262), .A4(new_n271), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n963), .B2(new_n817), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n256), .B1(new_n271), .B2(new_n262), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n918), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n840), .ZN(new_n977));
  INV_X1    g791(.A(new_n970), .ZN(new_n978));
  INV_X1    g792(.A(new_n296), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n281), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n977), .B2(new_n980), .ZN(G57));
endmodule


