//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G50), .B(G68), .Z(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  NAND3_X1  g0040(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(new_n210), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n245), .A2(new_n247), .B1(G150), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n203), .A2(G20), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n243), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT67), .B(G1), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n242), .B1(new_n252), .B2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G50), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(G13), .A4(G20), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(G50), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT9), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT70), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n256), .A3(new_n258), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G226), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n255), .A2(G274), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT66), .B(G45), .Z(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n268), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G222), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G223), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n266), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n276), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G190), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n261), .A2(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(G200), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n263), .A2(new_n294), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n294), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n300), .A2(new_n263), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n261), .B1(new_n305), .B2(new_n292), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n293), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n247), .A2(G77), .B1(G20), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n248), .A2(G50), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n243), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n315), .B(KEYINPUT11), .Z(new_n316));
  INV_X1    g0116(.A(new_n259), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n312), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n253), .A2(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n275), .A2(G238), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n226), .A2(G1698), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G226), .B2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n326), .B2(new_n288), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n279), .B1(new_n327), .B2(new_n267), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n323), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n323), .B2(new_n328), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n322), .B(G169), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n323), .A2(new_n328), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G179), .A3(new_n330), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n330), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n322), .B1(new_n338), .B2(G169), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n321), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(G200), .ZN(new_n341));
  INV_X1    g0141(.A(new_n321), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n338), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n253), .A2(G77), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G77), .B2(new_n259), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n245), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT69), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT15), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G87), .ZN(new_n351));
  INV_X1    g0151(.A(G87), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(KEYINPUT15), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(KEYINPUT15), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(G87), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT69), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n247), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n348), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n347), .B1(new_n360), .B2(new_n242), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n275), .A2(G244), .ZN(new_n362));
  NOR2_X1   g0162(.A1(G232), .A2(G1698), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n282), .A2(G238), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n280), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G107), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n266), .B1(new_n288), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n279), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n361), .B1(new_n305), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(new_n368), .A3(new_n307), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(G200), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n361), .C1(new_n343), .C2(new_n369), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n311), .A2(new_n345), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n259), .A2(new_n244), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n253), .B2(new_n244), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT72), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n285), .A2(new_n287), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n246), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n211), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n385), .A3(new_n211), .A4(new_n382), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(G68), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G58), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n312), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n201), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n248), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n243), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n385), .B1(new_n280), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n312), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(new_n392), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n379), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(G223), .A2(G1698), .ZN(new_n401));
  INV_X1    g0201(.A(G226), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n381), .B2(new_n382), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n246), .A2(new_n352), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n267), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT68), .B1(new_n252), .B2(new_n270), .ZN(new_n408));
  AND4_X1   g0208(.A1(KEYINPUT68), .A2(new_n270), .A3(new_n256), .A4(new_n258), .ZN(new_n409));
  OAI211_X1 g0209(.A(G232), .B(new_n266), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n279), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n407), .A2(new_n410), .A3(new_n343), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT17), .B1(new_n400), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n246), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n280), .B2(new_n380), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n385), .B1(new_n420), .B2(new_n211), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n386), .A2(G68), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n394), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n399), .A3(new_n242), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n378), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n412), .A2(G169), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n279), .B1(new_n275), .B2(G232), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(G179), .A3(new_n407), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT18), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n425), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n400), .A2(new_n416), .A3(KEYINPUT17), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n418), .A2(new_n431), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n376), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G257), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G250), .B2(G1698), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n382), .B2(new_n381), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G294), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT88), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT88), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(new_n442), .C1(new_n420), .C2(new_n440), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n267), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G274), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n264), .B2(new_n265), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT5), .B(G41), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n252), .A4(G45), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n256), .A2(new_n258), .A3(G45), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G41), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n266), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G264), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n447), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n305), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n447), .A2(new_n307), .A3(new_n451), .A4(new_n459), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT86), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(KEYINPUT25), .C1(new_n259), .C2(G107), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n256), .A2(new_n258), .A3(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(KEYINPUT25), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT25), .ZN(new_n467));
  AOI21_X1  g0267(.A(G107), .B1(new_n467), .B2(KEYINPUT86), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(G13), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n256), .A2(new_n258), .A3(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n259), .A2(new_n243), .A3(new_n470), .A4(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n464), .A2(new_n469), .A3(KEYINPUT87), .A4(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT22), .A2(G87), .ZN(new_n478));
  AOI211_X1 g0278(.A(G20), .B(new_n478), .C1(new_n381), .C2(new_n382), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n352), .A2(G20), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n288), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n211), .B2(G107), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n366), .A2(KEYINPUT23), .A3(G20), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n485), .A2(new_n486), .B1(new_n247), .B2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n477), .B1(new_n479), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n486), .ZN(new_n490));
  INV_X1    g0290(.A(G116), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n359), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT22), .B1(new_n280), .B2(new_n481), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n381), .A2(new_n382), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT24), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n497), .A3(new_n242), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n476), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n461), .A2(new_n462), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n461), .A2(new_n499), .A3(KEYINPUT89), .A4(new_n462), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n438), .A2(new_n282), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n458), .A2(G1698), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n495), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G303), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n280), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n267), .ZN(new_n512));
  OAI211_X1 g0312(.A(G270), .B(new_n266), .C1(new_n452), .C2(new_n456), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n451), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n513), .B2(new_n451), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  INV_X1    g0319(.A(G97), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n211), .C1(G33), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n491), .A2(G20), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n242), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT20), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(KEYINPUT85), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n259), .A2(new_n491), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n259), .A2(new_n243), .A3(new_n470), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(new_n491), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT85), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n523), .A2(new_n532), .A3(new_n524), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n518), .A2(new_n534), .A3(KEYINPUT21), .A4(G169), .ZN(new_n535));
  INV_X1    g0335(.A(new_n517), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n515), .B1(new_n267), .B2(new_n511), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(G179), .A3(new_n534), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n518), .A2(new_n534), .A3(G169), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n534), .B1(new_n518), .B2(G200), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n343), .B2(new_n518), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n499), .ZN(new_n546));
  INV_X1    g0346(.A(new_n459), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n442), .B1(new_n420), .B2(new_n440), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n266), .B1(new_n548), .B2(KEYINPUT88), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n549), .B2(new_n446), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT90), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n343), .A4(new_n451), .ZN(new_n552));
  AOI21_X1  g0352(.A(G200), .B1(new_n550), .B2(new_n451), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n447), .A2(new_n343), .A3(new_n451), .A4(new_n459), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT90), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n546), .B(new_n552), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n504), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g0357(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n282), .A2(G244), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n495), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G250), .A2(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n280), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n519), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n267), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(new_n266), .C1(new_n452), .C2(new_n456), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n451), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n568), .A2(KEYINPUT75), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT75), .B1(new_n568), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n305), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n259), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n530), .B2(G97), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n280), .A2(new_n385), .A3(G20), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT7), .B1(new_n288), .B2(new_n211), .ZN(new_n578));
  OAI21_X1  g0378(.A(G107), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  AND2_X1   g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G97), .A2(G107), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(KEYINPUT6), .A2(G97), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(G107), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT73), .B1(new_n589), .B2(new_n242), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT73), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n591), .B(new_n243), .C1(new_n579), .C2(new_n588), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n576), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n558), .B1(new_n420), .B2(new_n560), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n565), .A2(new_n280), .B1(G33), .B2(G283), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n266), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n596), .A2(G179), .A3(new_n570), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n574), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT76), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n366), .B1(new_n396), .B2(new_n397), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n248), .A2(G77), .ZN(new_n602));
  XNOR2_X1  g0402(.A(G97), .B(G107), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n585), .B1(new_n603), .B2(new_n580), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n604), .B2(new_n211), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n242), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n591), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n589), .A2(KEYINPUT73), .A3(new_n242), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n597), .B1(new_n609), .B2(new_n576), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT76), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n574), .ZN(new_n612));
  INV_X1    g0412(.A(new_n576), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n607), .B2(new_n608), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n568), .A2(new_n571), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT75), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n596), .B2(new_n570), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n568), .A2(KEYINPUT75), .A3(new_n571), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n614), .B(new_n616), .C1(new_n620), .C2(new_n343), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n600), .A2(new_n612), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n452), .A2(G250), .A3(new_n266), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n449), .A2(G45), .A3(new_n252), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT77), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n623), .B2(new_n624), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT83), .ZN(new_n630));
  INV_X1    g0430(.A(G244), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G1698), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G238), .B2(G1698), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n381), .B2(new_n382), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n246), .A2(new_n491), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n267), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n629), .A2(new_n630), .A3(G190), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(new_n624), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT77), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n636), .A3(G190), .A4(new_n626), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT83), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n636), .A3(new_n626), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G200), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n495), .A2(new_n211), .A3(G68), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT19), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n359), .B2(new_n520), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n324), .B2(new_n211), .ZN(new_n648));
  NOR2_X1   g0448(.A1(G87), .A2(G97), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n649), .A2(KEYINPUT78), .A3(new_n366), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT78), .B1(new_n649), .B2(new_n366), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n645), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(new_n242), .B1(new_n317), .B2(new_n358), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n529), .A2(new_n352), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n644), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n642), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT80), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT79), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT69), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT69), .B1(new_n355), .B2(new_n356), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n354), .A2(KEYINPUT79), .A3(new_n357), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n666), .B2(new_n530), .ZN(new_n667));
  AOI211_X1 g0467(.A(KEYINPUT80), .B(new_n529), .C1(new_n664), .C2(new_n665), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n654), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT81), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT81), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n654), .B(new_n671), .C1(new_n667), .C2(new_n668), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n643), .A2(G179), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n305), .B2(new_n643), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n659), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n622), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n437), .A2(new_n557), .A3(new_n677), .ZN(G372));
  AND3_X1   g0478(.A1(new_n425), .A2(new_n429), .A3(new_n432), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n432), .B1(new_n425), .B2(new_n429), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n344), .A2(new_n371), .A3(new_n370), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n340), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n400), .A2(new_n416), .A3(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n417), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n681), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n304), .ZN(new_n688));
  INV_X1    g0488(.A(new_n672), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n662), .A2(new_n663), .A3(new_n661), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT79), .B1(new_n354), .B2(new_n357), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n530), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT80), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n666), .A2(new_n660), .A3(new_n530), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n671), .B1(new_n695), .B2(new_n654), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n675), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n644), .A2(new_n657), .A3(new_n654), .A4(new_n640), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n697), .A2(new_n556), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(G169), .B1(new_n618), .B2(new_n619), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n700), .A2(new_n614), .A3(KEYINPUT76), .A4(new_n597), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n611), .B1(new_n610), .B2(new_n574), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n539), .A2(new_n500), .A3(new_n542), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n699), .A2(new_n703), .A3(new_n621), .A4(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n700), .A2(new_n614), .A3(new_n597), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n697), .A2(new_n706), .A3(new_n707), .A4(new_n698), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n673), .A2(new_n710), .A3(new_n675), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n697), .B1(new_n658), .B2(new_n642), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT26), .B1(new_n703), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n705), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n310), .B(new_n688), .C1(new_n437), .C2(new_n716), .ZN(G369));
  NAND2_X1  g0517(.A1(new_n539), .A2(new_n542), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n211), .A2(G13), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n252), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G213), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G343), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n534), .A2(new_n725), .ZN(new_n726));
  MUX2_X1   g0526(.A(new_n718), .B(new_n545), .S(new_n726), .Z(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n556), .A2(new_n502), .A3(new_n503), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n725), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n546), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n500), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n725), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n718), .A2(new_n732), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n730), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n734), .B2(new_n732), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(G399));
  INV_X1    g0541(.A(new_n207), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G41), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G1), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n650), .A2(new_n651), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n491), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n747), .B1(new_n214), .B2(new_n744), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n502), .A2(new_n503), .A3(new_n542), .A4(new_n539), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n622), .A2(new_n699), .A3(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n676), .B(new_n707), .C1(new_n702), .C2(new_n701), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n709), .A2(new_n711), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n697), .A2(new_n698), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT26), .B1(new_n754), .B2(new_n599), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n732), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT29), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n715), .A2(new_n759), .A3(new_n732), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G330), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n460), .A2(new_n615), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT92), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n460), .A2(KEYINPUT92), .A3(new_n615), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n639), .A2(new_n636), .A3(new_n626), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n537), .A2(new_n767), .A3(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT30), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n550), .A2(new_n537), .A3(G179), .A4(new_n767), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n620), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n572), .A2(new_n573), .ZN(new_n773));
  AND3_X1   g0573(.A1(new_n767), .A2(new_n459), .A3(new_n447), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n512), .B(G179), .C1(new_n516), .C2(new_n517), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT30), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n778), .A2(KEYINPUT31), .A3(new_n725), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT31), .B1(new_n778), .B2(new_n725), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n730), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n783), .A2(new_n622), .A3(new_n676), .A4(new_n732), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n762), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n761), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n749), .B1(new_n788), .B2(G1), .ZN(G364));
  AOI21_X1  g0589(.A(new_n255), .B1(new_n719), .B2(G45), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n743), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n729), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G330), .B2(new_n727), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n210), .B1(G20), .B2(new_n305), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n211), .A2(new_n343), .A3(new_n413), .A4(G179), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n352), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n211), .A2(G190), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n307), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n801), .A2(G20), .A3(G190), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n280), .B1(new_n802), .B2(new_n289), .C1(new_n388), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n211), .A2(new_n307), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n343), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n799), .B(new_n804), .C1(G68), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G179), .A2(G200), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n211), .B1(new_n809), .B2(G190), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT95), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G97), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n800), .A2(new_n809), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n211), .A2(new_n413), .A3(G179), .A4(G190), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n366), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n805), .A2(G190), .A3(G200), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(G50), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n808), .A2(new_n812), .A3(new_n817), .A4(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G322), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n803), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n288), .B1(new_n802), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n813), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n828), .C1(G329), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n822), .A2(G326), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n807), .A2(new_n832), .B1(new_n797), .B2(G303), .ZN(new_n833));
  INV_X1    g0633(.A(new_n810), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(G294), .B1(new_n818), .B2(G283), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n796), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(G13), .A2(G33), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(G20), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n795), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n420), .A2(new_n207), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT93), .ZN(new_n844));
  INV_X1    g0644(.A(new_n278), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n269), .B2(new_n236), .C1(new_n215), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n742), .A2(new_n288), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G355), .B1(new_n491), .B2(new_n742), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n842), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n792), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n837), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n840), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n727), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n794), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NOR2_X1   g0655(.A1(new_n372), .A2(new_n725), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n374), .B1(new_n361), .B2(new_n732), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n372), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n716), .B2(new_n725), .ZN(new_n861));
  INV_X1    g0661(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n715), .A2(new_n732), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n792), .B1(new_n864), .B2(new_n786), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n786), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n795), .A2(new_n838), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n850), .B1(new_n289), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G294), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n812), .B1(new_n869), .B2(new_n803), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT96), .ZN(new_n871));
  INV_X1    g0671(.A(G283), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n798), .A2(new_n366), .B1(new_n872), .B2(new_n806), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n288), .B1(new_n813), .B2(new_n827), .C1(new_n491), .C2(new_n802), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n819), .A2(new_n352), .B1(new_n508), .B2(new_n821), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n803), .ZN(new_n877));
  INV_X1    g0677(.A(new_n802), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(G143), .B1(new_n878), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n880), .B2(new_n821), .C1(new_n881), .C2(new_n806), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT34), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n798), .A2(new_n202), .B1(new_n819), .B2(new_n312), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT97), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  INV_X1    g0687(.A(G132), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n495), .B1(new_n388), .B2(new_n810), .C1(new_n888), .C2(new_n813), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n871), .A2(new_n876), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n868), .B1(new_n796), .B2(new_n891), .C1(new_n862), .C2(new_n839), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n866), .A2(new_n892), .ZN(G384));
  OAI211_X1 g0693(.A(G116), .B(new_n212), .C1(new_n587), .C2(KEYINPUT35), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT98), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n587), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(KEYINPUT98), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  OAI21_X1  g0699(.A(G77), .B1(new_n388), .B2(new_n312), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n900), .A2(new_n214), .B1(G50), .B2(new_n312), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n252), .A2(G13), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n321), .A2(new_n725), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n340), .A2(new_n344), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n340), .B2(new_n344), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n863), .B2(new_n857), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(new_n723), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n423), .A2(new_n242), .ZN(new_n912));
  INV_X1    g0712(.A(new_n392), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT16), .B1(new_n387), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n378), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n911), .A2(new_n915), .B1(new_n400), .B2(new_n416), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n429), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n425), .A2(new_n911), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n400), .A2(new_n416), .ZN(new_n920));
  AND4_X1   g0720(.A1(new_n910), .A2(new_n430), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n387), .A2(new_n913), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n393), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n379), .B1(new_n924), .B2(new_n395), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n723), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n681), .B2(new_n685), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n909), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n723), .B2(new_n925), .ZN(new_n930));
  INV_X1    g0730(.A(new_n917), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n430), .A2(new_n919), .A3(new_n920), .A4(new_n910), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n435), .A2(new_n926), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT38), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(KEYINPUT99), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT99), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(new_n909), .C1(new_n922), .C2(new_n928), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n681), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n908), .A2(new_n941), .B1(new_n942), .B2(new_n723), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n430), .A2(new_n919), .A3(new_n920), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n910), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n919), .B1(new_n681), .B2(new_n685), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT39), .B1(new_n948), .B2(new_n936), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n940), .B2(KEYINPUT39), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n340), .A2(new_n725), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n943), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT101), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n943), .A2(KEYINPUT101), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n437), .B1(new_n758), .B2(new_n760), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n688), .A2(new_n310), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n958), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n778), .A2(new_n725), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT31), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n778), .A2(KEYINPUT31), .A3(new_n725), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n703), .A2(new_n621), .A3(new_n676), .A4(new_n732), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n966), .C1(new_n967), .C2(new_n557), .ZN(new_n968));
  INV_X1    g0768(.A(new_n906), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n340), .A2(new_n344), .A3(new_n904), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n860), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n937), .A2(new_n968), .A3(new_n939), .A4(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT40), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n862), .B1(new_n905), .B2(new_n906), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n781), .B2(new_n784), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n973), .B1(new_n948), .B2(new_n936), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT102), .Z(new_n980));
  NAND3_X1  g0780(.A1(new_n376), .A2(new_n436), .A3(new_n968), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT103), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n762), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n980), .B2(new_n982), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n962), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n252), .B2(new_n719), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n962), .A2(new_n984), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n903), .B1(new_n986), .B2(new_n987), .ZN(G367));
  OAI21_X1  g0788(.A(new_n622), .B1(new_n614), .B2(new_n732), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n706), .A2(new_n725), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n739), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT42), .Z(new_n993));
  INV_X1    g0793(.A(new_n991), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n703), .B1(new_n994), .B2(new_n504), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n732), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n732), .B1(new_n654), .B2(new_n657), .ZN(new_n998));
  MUX2_X1   g0798(.A(new_n754), .B(new_n753), .S(new_n998), .Z(new_n999));
  INV_X1    g0799(.A(KEYINPUT43), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT105), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n999), .A2(KEYINPUT104), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n999), .A2(KEYINPUT104), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n997), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n737), .B2(new_n994), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n737), .A2(new_n994), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n743), .B(KEYINPUT41), .Z(new_n1014));
  INV_X1    g0814(.A(KEYINPUT107), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT106), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n728), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n739), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n733), .A2(new_n735), .A3(new_n738), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1018), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1021), .A2(new_n1016), .A3(new_n728), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n788), .A2(new_n1015), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT45), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n740), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n994), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n991), .A2(new_n740), .A3(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n994), .A2(new_n1026), .A3(KEYINPUT44), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT44), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n991), .B2(new_n740), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1029), .A2(new_n737), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n737), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1023), .A2(new_n786), .A3(new_n761), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT107), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1024), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1014), .B1(new_n1039), .B2(new_n788), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1011), .B(new_n1013), .C1(new_n1040), .C2(new_n791), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n999), .A2(new_n840), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n844), .A2(new_n232), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n841), .C1(new_n207), .C2(new_n358), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n792), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT108), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n819), .A2(new_n289), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n798), .A2(new_n388), .B1(new_n814), .B2(new_n806), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G143), .C2(new_n822), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n811), .A2(G68), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n288), .B1(new_n877), .B2(G150), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT109), .B(G137), .Z(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n829), .A2(new_n1053), .B1(new_n878), .B2(G50), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n797), .A2(G116), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT46), .Z(new_n1057));
  OAI22_X1  g0857(.A1(new_n819), .A2(new_n520), .B1(new_n827), .B2(new_n821), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G294), .B2(new_n807), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n803), .A2(new_n508), .B1(new_n802), .B2(new_n872), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G317), .B2(new_n829), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n495), .B1(G107), .B2(new_n834), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1055), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n795), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1042), .B(new_n1046), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1041), .A2(new_n1069), .ZN(G387));
  AND2_X1   g0870(.A1(new_n1037), .A2(new_n743), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n788), .B2(new_n1023), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n733), .A2(new_n735), .A3(new_n840), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n747), .A2(new_n847), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(G107), .B2(new_n207), .ZN(new_n1075));
  AOI211_X1 g0875(.A(G45), .B(new_n747), .C1(G68), .C2(G77), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT111), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(KEYINPUT111), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n244), .A2(G50), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n844), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n229), .B2(new_n845), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1075), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n792), .B1(new_n1084), .B2(new_n842), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n797), .A2(G77), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n814), .B2(new_n821), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n245), .B2(new_n807), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n666), .A2(new_n811), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n802), .A2(new_n312), .B1(new_n813), .B2(new_n881), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G50), .B2(new_n877), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n420), .B1(G97), .B2(new_n818), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n797), .A2(G294), .B1(new_n834), .B2(G283), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n877), .A2(G317), .B1(new_n878), .B2(G303), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n827), .B2(new_n806), .C1(new_n825), .C2(new_n821), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT48), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT112), .Z(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(KEYINPUT49), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n495), .B1(G326), .B2(new_n829), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n491), .C2(new_n819), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT49), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1093), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1085), .B1(new_n1105), .B2(new_n795), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1023), .A2(new_n791), .B1(new_n1073), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1072), .A2(new_n1107), .ZN(G393));
  OAI21_X1  g0908(.A(new_n841), .B1(new_n520), .B2(new_n207), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n844), .B2(new_n239), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT113), .Z(new_n1111));
  OAI22_X1  g0911(.A1(new_n798), .A2(new_n312), .B1(new_n819), .B2(new_n352), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n420), .B(new_n1112), .C1(G143), .C2(new_n829), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n806), .A2(new_n202), .B1(new_n802), .B2(new_n244), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT114), .Z(new_n1115));
  OAI22_X1  g0915(.A1(new_n821), .A2(new_n881), .B1(new_n803), .B2(new_n814), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT51), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n811), .A2(G77), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G317), .A2(new_n822), .B1(new_n877), .B2(G311), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT52), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n798), .A2(new_n872), .B1(new_n491), .B2(new_n810), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n820), .B(new_n1122), .C1(G303), .C2(new_n807), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n288), .B1(new_n813), .B2(new_n825), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G294), .B2(new_n878), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n796), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1111), .A2(new_n1127), .A3(new_n850), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n991), .B2(new_n852), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1036), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n790), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n744), .B1(new_n1130), .B2(new_n1037), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1039), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(G390));
  NAND3_X1  g0934(.A1(new_n968), .A2(G330), .A3(new_n862), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n907), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n908), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n950), .B1(new_n1137), .B2(new_n951), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n948), .A2(new_n936), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n951), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n859), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n857), .B1(new_n757), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n907), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1136), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n950), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n952), .B2(new_n908), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n785), .A2(new_n862), .A3(new_n1143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1144), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(new_n790), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n867), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n819), .A2(new_n312), .B1(new_n869), .B2(new_n813), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT116), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT116), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1155), .A2(new_n1118), .A3(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n288), .B1(new_n802), .B2(new_n520), .C1(new_n491), .C2(new_n803), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n798), .A2(new_n352), .B1(new_n366), .B2(new_n806), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G283), .C2(new_n822), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n807), .A2(new_n1053), .B1(G50), .B2(new_n818), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n821), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n280), .B1(new_n803), .B2(new_n888), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n802), .A2(new_n1165), .B1(new_n813), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT53), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n798), .B2(new_n881), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n797), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G159), .A2(new_n811), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1157), .A2(new_n1160), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n792), .B1(new_n245), .B2(new_n1153), .C1(new_n1173), .C2(new_n796), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1146), .B2(new_n838), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1152), .A2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n622), .A2(new_n699), .A3(new_n750), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n725), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n856), .B1(new_n1179), .B2(new_n859), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1135), .A2(new_n907), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1148), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(KEYINPUT115), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT115), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1143), .B1(new_n785), .B2(new_n862), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1136), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n1186), .B2(new_n1180), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1181), .A2(new_n1148), .B1(new_n857), .B2(new_n863), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n437), .A2(new_n786), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n959), .A2(new_n1191), .A3(new_n960), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n1145), .A3(new_n1150), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1186), .A2(new_n1184), .A3(new_n1180), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1182), .A2(KEYINPUT115), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1192), .B(new_n1194), .C1(new_n1195), .C2(new_n1188), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1151), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1197), .A3(new_n743), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1176), .A2(new_n1198), .ZN(G378));
  NOR2_X1   g0999(.A1(new_n261), .A2(new_n723), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n311), .B(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1201), .B(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n762), .B1(new_n976), .B2(new_n977), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n974), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT119), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n974), .A2(KEYINPUT119), .A3(new_n1205), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1204), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT119), .B1(new_n974), .B2(new_n1205), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1201), .B(new_n1202), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n956), .B(new_n957), .C1(new_n1210), .C2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n974), .A2(KEYINPUT119), .A3(new_n1205), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1212), .B1(new_n1215), .B2(new_n1211), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1208), .A2(new_n1204), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n908), .A2(new_n941), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n942), .A2(new_n723), .ZN(new_n1219));
  AND4_X1   g1019(.A1(KEYINPUT101), .A2(new_n953), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT101), .B1(new_n943), .B2(new_n953), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1216), .B(new_n1217), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1214), .A2(KEYINPUT120), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1194), .B1(new_n1195), .B2(new_n1188), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1192), .B1(new_n1151), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT120), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n958), .A2(new_n1226), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1193), .B2(new_n1192), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1214), .A2(new_n1222), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n744), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1223), .A2(new_n791), .A3(new_n1227), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1212), .A2(new_n838), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n792), .B1(G50), .B2(new_n1153), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n420), .B2(new_n268), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n807), .A2(G97), .B1(G58), .B2(new_n818), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n491), .B2(new_n821), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1086), .B1(new_n366), .B2(new_n803), .C1(new_n872), .C2(new_n813), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1241), .A2(new_n1242), .A3(G41), .A4(new_n495), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n666), .A2(new_n878), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1050), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT58), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1239), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n798), .A2(new_n1165), .B1(new_n1162), .B2(new_n803), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT118), .Z(new_n1249));
  OAI22_X1  g1049(.A1(new_n806), .A2(new_n888), .B1(new_n802), .B2(new_n880), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT117), .Z(new_n1251));
  AOI22_X1  g1051(.A1(new_n811), .A2(G150), .B1(G125), .B2(new_n822), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n818), .A2(G159), .ZN(new_n1255));
  AOI211_X1 g1055(.A(G33), .B(G41), .C1(new_n829), .C2(G124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1247), .B1(new_n1246), .B2(new_n1245), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1237), .B1(new_n1259), .B2(new_n795), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1236), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1235), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1234), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT121), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1262), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT121), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1266), .A2(new_n1270), .ZN(G375));
  XNOR2_X1  g1071(.A(new_n790), .B(KEYINPUT122), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n907), .A2(new_n838), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n819), .A2(new_n289), .B1(new_n806), .B2(new_n491), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n288), .B1(new_n802), .B2(new_n366), .C1(new_n872), .C2(new_n803), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(G294), .C2(new_n822), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(G303), .A2(new_n829), .B1(new_n797), .B2(G97), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(KEYINPUT123), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1089), .A3(new_n1279), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n888), .A2(new_n821), .B1(new_n806), .B2(new_n1165), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G159), .B2(new_n797), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n811), .A2(G50), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1052), .A2(new_n803), .B1(new_n813), .B2(new_n1162), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G150), .B2(new_n878), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n420), .B1(G58), .B2(new_n818), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1282), .A2(new_n1283), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n796), .B1(new_n1280), .B2(new_n1287), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n850), .B(new_n1288), .C1(new_n312), .C2(new_n867), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1190), .A2(new_n1273), .B1(new_n1274), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1196), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1291), .A2(new_n1014), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1192), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1224), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1290), .B1(new_n1292), .B2(new_n1295), .ZN(G381));
  AND3_X1   g1096(.A1(new_n1176), .A2(new_n1198), .A3(KEYINPUT124), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT124), .B1(new_n1176), .B2(new_n1198), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1041), .A2(new_n1069), .A3(new_n1133), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1072), .A2(new_n854), .A3(new_n1107), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(new_n1300), .A2(G384), .A3(G381), .A4(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1299), .B(new_n1302), .C1(new_n1266), .C2(new_n1270), .ZN(G407));
  OAI21_X1  g1103(.A(new_n1299), .B1(new_n1266), .B2(new_n1270), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G407), .B(G213), .C1(new_n1304), .C2(G343), .ZN(G409));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1232), .A2(new_n1273), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1261), .B(new_n1307), .C1(new_n1228), .C2(new_n1014), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1267), .A2(G378), .B1(new_n1299), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n724), .A2(G213), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1306), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1234), .A2(G378), .A3(new_n1263), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1298), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1176), .A2(new_n1198), .A3(KEYINPUT124), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1308), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1311), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT125), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1294), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n743), .B(new_n1196), .C1(new_n1294), .C2(new_n1319), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1290), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n866), .A3(new_n892), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G384), .B(new_n1290), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1311), .A2(G2897), .ZN(new_n1327));
  XOR2_X1   g1127(.A(new_n1327), .B(KEYINPUT126), .Z(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1324), .A2(new_n1325), .A3(new_n1328), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1312), .A2(new_n1318), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1301), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n854), .B1(new_n1072), .B2(new_n1107), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1041), .A2(new_n1069), .A3(new_n1133), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1133), .B1(new_n1041), .B2(new_n1069), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1337), .B(new_n1338), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G387), .A2(G390), .ZN(new_n1342));
  OAI21_X1  g1142(.A(KEYINPUT127), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1342), .A2(new_n1300), .A3(new_n1343), .A4(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT61), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1341), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1326), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1310), .A3(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1347), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1349), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1334), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT62), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1317), .A2(new_n1355), .A3(new_n1349), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1346), .B1(new_n1317), .B2(new_n1332), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1355), .B1(new_n1317), .B2(new_n1349), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1356), .A2(new_n1357), .A3(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1354), .B1(new_n1359), .B2(new_n1361), .ZN(G405));
  NAND3_X1  g1162(.A1(new_n1265), .A2(new_n1269), .A3(new_n1299), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1363), .A2(new_n1313), .A3(new_n1326), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1326), .B1(new_n1363), .B2(new_n1313), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1360), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1366), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1368), .A2(new_n1361), .A3(new_n1364), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1367), .A2(new_n1369), .ZN(G402));
endmodule


