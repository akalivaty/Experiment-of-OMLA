//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n214), .A2(G50), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n211), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n220), .B1(new_n223), .B2(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n218), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT67), .Z(G361));
  XOR2_X1   g0032(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT69), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(KEYINPUT70), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT70), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n253), .B(new_n205), .C1(new_n256), .C2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(G226), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n251), .A2(new_n252), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n257), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n265), .B1(new_n266), .B2(new_n263), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n259), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(G190), .ZN(new_n274));
  XOR2_X1   g0074(.A(KEYINPUT8), .B(G58), .Z(new_n275));
  NAND2_X1  g0075(.A1(new_n206), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n275), .A2(new_n277), .B1(G150), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n212), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n205), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  XOR2_X1   g0090(.A(new_n290), .B(KEYINPUT71), .Z(new_n291));
  OAI221_X1 g0091(.A(new_n284), .B1(G50), .B2(new_n285), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n273), .B(new_n274), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT73), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n273), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n295), .B(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT72), .B1(new_n271), .B2(G169), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n271), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT72), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n303), .B(new_n292), .C1(new_n304), .C2(new_n302), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G68), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n286), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n266), .B2(new_n276), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n287), .A2(G68), .A3(new_n289), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT11), .B1(new_n311), .B2(new_n283), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n256), .ZN(new_n318));
  INV_X1    g0118(.A(G45), .ZN(new_n319));
  AOI21_X1  g0119(.A(G1), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n261), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n253), .A2(new_n320), .B1(new_n321), .B2(G238), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n263), .A2(G226), .A3(new_n264), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n270), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n322), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n322), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(G169), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n322), .A2(new_n327), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n322), .A2(new_n327), .A3(new_n328), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n331), .A2(KEYINPUT14), .B1(new_n335), .B2(new_n301), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n335), .B2(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n317), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(G200), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n333), .A2(G190), .A3(new_n334), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n316), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n275), .A2(new_n289), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n288), .A2(new_n344), .B1(new_n285), .B2(new_n275), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT16), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n263), .B2(G20), .ZN(new_n348));
  INV_X1    g0148(.A(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n307), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G58), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n307), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n357), .B2(new_n201), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n278), .A2(G159), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n346), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n283), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n348), .A2(new_n354), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(G68), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT74), .B1(new_n364), .B2(KEYINPUT16), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n345), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G232), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n257), .B1(new_n369), .B2(new_n261), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n350), .A2(new_n352), .A3(G226), .A4(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n268), .A2(G1698), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n263), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n350), .A3(new_n352), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n374), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n371), .B(new_n301), .C1(new_n380), .C2(new_n259), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n377), .ZN(new_n382));
  INV_X1    g0182(.A(new_n374), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n259), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n370), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n385), .B2(G169), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT18), .B1(new_n368), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n363), .A2(G68), .ZN(new_n388));
  INV_X1    g0188(.A(new_n360), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n392), .A2(new_n283), .A3(new_n367), .A4(new_n361), .ZN(new_n393));
  INV_X1    g0193(.A(new_n345), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n386), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n371), .B(new_n399), .C1(new_n380), .C2(new_n259), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n272), .B1(new_n384), .B2(new_n370), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n393), .A2(new_n394), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT76), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n393), .A2(new_n394), .A3(new_n402), .A4(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n387), .A2(new_n398), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n287), .A2(G77), .A3(new_n289), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G77), .B2(new_n285), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n282), .A2(new_n212), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n275), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n277), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n321), .A2(G244), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n257), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n263), .A2(G232), .A3(new_n264), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  INV_X1    g0222(.A(G238), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n421), .B1(new_n422), .B2(new_n263), .C1(new_n267), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n420), .B1(new_n424), .B2(new_n270), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n418), .B1(new_n425), .B2(G190), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n272), .B2(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n424), .A2(new_n270), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n420), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n425), .A2(new_n301), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n418), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n306), .A2(new_n343), .A3(new_n409), .A4(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n350), .A2(new_n352), .A3(G257), .A4(G1698), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n350), .A2(new_n352), .A3(G250), .A4(new_n264), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G294), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n270), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT5), .B1(new_n254), .B2(new_n255), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT5), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n205), .B(G45), .C1(new_n441), .C2(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(G264), .B(new_n259), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n255), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT70), .A2(G41), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n442), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n253), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT82), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n439), .A2(new_n453), .A3(new_n443), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n452), .A2(new_n454), .A3(G179), .A4(new_n449), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n350), .A2(new_n352), .A3(new_n206), .A4(G87), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT22), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT80), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G116), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G20), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n206), .A2(KEYINPUT80), .A3(G33), .A4(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n263), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n422), .A3(G20), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n458), .A2(new_n464), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n471), .A2(new_n473), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n283), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n205), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n412), .A2(KEYINPUT78), .A3(new_n285), .A4(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n285), .A2(new_n477), .A3(new_n212), .A4(new_n282), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT25), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n285), .B2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n422), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n482), .A2(G107), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n451), .A2(new_n455), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n476), .A2(new_n486), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n439), .A2(new_n399), .A3(new_n449), .A4(new_n443), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n439), .A2(new_n453), .A3(new_n443), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n453), .B1(new_n439), .B2(new_n443), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n490), .A2(new_n491), .A3(new_n450), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(G200), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n487), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n350), .A2(new_n352), .A3(G244), .A4(new_n264), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n264), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n270), .ZN(new_n502));
  OAI211_X1 g0302(.A(G257), .B(new_n259), .C1(new_n440), .C2(new_n442), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n503), .A2(new_n449), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n504), .A3(new_n399), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n449), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n270), .B2(new_n501), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n507), .B2(G200), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n278), .A2(G77), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n510), .A2(new_n511), .A3(G107), .ZN(new_n512));
  XNOR2_X1  g0312(.A(G97), .B(G107), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n510), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n514), .B2(new_n206), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n422), .B1(new_n348), .B2(new_n354), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n283), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n478), .A2(new_n481), .A3(G97), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n285), .A2(G97), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n508), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n206), .B1(new_n325), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G87), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n511), .A3(new_n422), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n350), .A2(new_n352), .A3(new_n206), .A4(G68), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n526), .B1(new_n276), .B2(new_n511), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n283), .B1(new_n286), .B2(new_n414), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n478), .A2(new_n481), .A3(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n205), .A2(new_n250), .A3(G45), .ZN(new_n537));
  INV_X1    g0337(.A(G250), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n319), .B2(G1), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n259), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n350), .A2(new_n352), .A3(G244), .A4(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n350), .A2(new_n352), .A3(G238), .A4(new_n264), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n460), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n399), .B(new_n540), .C1(new_n543), .C2(new_n270), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n270), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n259), .A2(new_n537), .A3(new_n539), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n478), .A2(new_n481), .A3(new_n415), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n540), .B1(new_n543), .B2(new_n270), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n534), .A2(new_n550), .B1(new_n551), .B2(new_n301), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n428), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n545), .A2(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n502), .A2(new_n504), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n428), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n507), .A2(new_n301), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n523), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n525), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G270), .B(new_n259), .C1(new_n440), .C2(new_n442), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n560), .A2(new_n449), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n353), .A2(G303), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n350), .A2(new_n352), .A3(G257), .A4(new_n264), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n350), .A2(new_n352), .A3(G264), .A4(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n263), .A2(KEYINPUT79), .A3(G264), .A4(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n561), .B(G190), .C1(new_n569), .C2(new_n259), .ZN(new_n570));
  INV_X1    g0370(.A(G116), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n286), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n479), .B2(new_n571), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n282), .A2(new_n212), .B1(G20), .B2(new_n571), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n499), .B(new_n206), .C1(G33), .C2(new_n511), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n564), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n567), .A2(new_n568), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n259), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n560), .A2(new_n449), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n570), .B(new_n580), .C1(new_n585), .C2(new_n272), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n583), .A2(new_n301), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(new_n576), .ZN(new_n588));
  INV_X1    g0388(.A(new_n573), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(G169), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n585), .A2(new_n592), .A3(KEYINPUT21), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n561), .B1(new_n569), .B2(new_n259), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n580), .A2(new_n428), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n586), .B(new_n591), .C1(new_n593), .C2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n559), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n434), .A2(new_n494), .A3(new_n599), .ZN(G372));
  AND3_X1   g0400(.A1(new_n340), .A2(new_n316), .A3(new_n341), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n339), .B1(new_n601), .B2(new_n432), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n406), .A2(new_n408), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n386), .B1(new_n393), .B2(new_n394), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n397), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n368), .A2(KEYINPUT18), .A3(new_n386), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n299), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(new_n305), .ZN(new_n611));
  INV_X1    g0411(.A(new_n546), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n547), .A2(KEYINPUT83), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n259), .A2(new_n614), .A3(new_n537), .A4(new_n539), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n428), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n552), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n507), .A2(new_n301), .B1(new_n517), .B2(new_n522), .ZN(new_n619));
  OAI21_X1  g0419(.A(G200), .B1(new_n612), .B2(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n533), .A2(new_n283), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n414), .A2(new_n286), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n535), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n551), .A2(G190), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n619), .A2(new_n618), .A3(new_n625), .A4(new_n556), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n618), .B1(new_n626), .B2(KEYINPUT26), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n556), .A2(new_n557), .A3(new_n523), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n554), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT84), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n545), .A2(new_n549), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n552), .A2(new_n553), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT26), .B1(new_n634), .B2(new_n558), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n545), .A2(new_n620), .B1(new_n552), .B2(new_n617), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n628), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n637), .A3(new_n638), .A4(new_n618), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n455), .A2(new_n451), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n476), .A2(new_n486), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT21), .B1(new_n585), .B2(new_n592), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n595), .A2(new_n596), .A3(new_n594), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n645), .A3(new_n591), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n525), .A2(new_n636), .A3(new_n558), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n493), .A2(new_n488), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n631), .A2(new_n639), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n434), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n611), .A2(new_n651), .ZN(G369));
  OAI21_X1  g0452(.A(new_n591), .B1(new_n593), .B2(new_n597), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(G213), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n494), .B1(new_n488), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n487), .A2(new_n659), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT85), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n661), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n642), .A2(new_n659), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n667), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n660), .A2(new_n580), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n653), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n598), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(G399));
  NAND2_X1  g0478(.A1(new_n209), .A2(new_n318), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n529), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n216), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n556), .A2(new_n619), .B1(new_n508), .B2(new_n524), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n648), .A2(new_n684), .A3(new_n636), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n653), .A2(new_n487), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT89), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n646), .A2(new_n647), .A3(new_n688), .A4(new_n648), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n628), .B1(new_n634), .B2(new_n558), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n690), .B(KEYINPUT88), .C1(new_n628), .C2(new_n626), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n626), .A2(KEYINPUT88), .A3(new_n628), .ZN(new_n692));
  INV_X1    g0492(.A(new_n618), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n687), .A2(new_n689), .A3(new_n691), .A4(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n660), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT90), .B1(new_n695), .B2(new_n660), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT29), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT87), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n650), .A2(new_n660), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI211_X1 g0502(.A(KEYINPUT87), .B(KEYINPUT29), .C1(new_n650), .C2(new_n660), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n599), .A2(new_n494), .A3(new_n660), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n551), .A2(G179), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n585), .A2(new_n710), .A3(new_n507), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n452), .A2(new_n454), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n452), .A2(new_n454), .A3(new_n449), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n612), .A2(new_n616), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n716), .A3(new_n595), .A4(new_n555), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n595), .A2(new_n709), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n490), .A2(new_n491), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n507), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n713), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n659), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n707), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n659), .A2(KEYINPUT31), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT86), .B1(new_n713), .B2(new_n717), .ZN(new_n727));
  INV_X1    g0527(.A(new_n720), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n713), .A2(KEYINPUT86), .A3(new_n717), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(G330), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n706), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n683), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n679), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n206), .A2(G13), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n205), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n676), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G330), .B2(new_n674), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n209), .A2(new_n263), .ZN(new_n742));
  INV_X1    g0542(.A(G355), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n743), .B1(G116), .B2(new_n209), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n245), .A2(new_n319), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n209), .A2(new_n353), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n217), .B2(new_n319), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n744), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n212), .B1(G20), .B2(new_n428), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n739), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n206), .A2(new_n301), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n399), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G50), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n206), .A2(new_n399), .A3(new_n272), .A4(G179), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n759), .A2(new_n760), .B1(new_n528), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n756), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n764), .A2(new_n399), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n263), .B1(new_n766), .B2(new_n356), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G20), .A3(new_n399), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n763), .B(new_n767), .C1(KEYINPUT32), .C2(new_n772), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n206), .A2(new_n272), .A3(G179), .A4(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n422), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n206), .B1(new_n768), .B2(G190), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n772), .A2(KEYINPUT32), .B1(new_n511), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n757), .A2(G190), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n776), .B(new_n778), .C1(G68), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT91), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT91), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n773), .B(new_n780), .C1(new_n266), .C2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n769), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G329), .ZN(new_n787));
  INV_X1    g0587(.A(new_n781), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n263), .B(new_n790), .C1(G322), .C2(new_n765), .ZN(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n779), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n777), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n761), .A2(G303), .B1(new_n796), .B2(G294), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n758), .A2(G326), .B1(G283), .B2(new_n774), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n791), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n785), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n755), .B1(new_n800), .B2(new_n752), .ZN(new_n801));
  INV_X1    g0601(.A(new_n751), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n674), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n741), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n432), .A2(KEYINPUT93), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n418), .A2(new_n659), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT93), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n430), .A2(new_n431), .A3(new_n808), .A4(new_n418), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n806), .A2(new_n427), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n432), .A2(new_n660), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT94), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n810), .A2(KEYINPUT94), .A3(new_n811), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n700), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n806), .A2(new_n809), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(new_n427), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n650), .A2(new_n660), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n739), .B1(new_n820), .B2(new_n732), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n732), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n752), .A2(new_n749), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n739), .B1(G77), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT92), .Z(new_n826));
  INV_X1    g0626(.A(new_n779), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n766), .A2(new_n830), .B1(new_n759), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n784), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n829), .B(new_n832), .C1(new_n833), .C2(G159), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n263), .B1(new_n769), .B2(new_n837), .C1(new_n356), .C2(new_n777), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n762), .A2(new_n760), .B1(new_n775), .B2(new_n307), .ZN(new_n839));
  OR4_X1    g0639(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n833), .A2(G116), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n827), .A2(new_n842), .B1(new_n422), .B2(new_n762), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G303), .B2(new_n758), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n353), .B1(new_n769), .B2(new_n789), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n765), .B2(G294), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n796), .A2(G97), .B1(new_n774), .B2(G87), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n841), .A2(new_n844), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n752), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n826), .B1(new_n750), .B2(new_n812), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n822), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  INV_X1    g0653(.A(new_n514), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT35), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(KEYINPUT35), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(G116), .A3(new_n213), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT36), .Z(new_n858));
  OR3_X1    g0658(.A1(new_n216), .A2(new_n266), .A3(new_n357), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n760), .A2(G68), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n205), .B(G13), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n698), .A2(new_n704), .A3(new_n434), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n611), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT97), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n605), .B1(new_n368), .B2(new_n402), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n657), .B(KEYINPUT96), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n395), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n605), .ZN(new_n871));
  INV_X1    g0671(.A(new_n657), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n395), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n871), .A2(new_n873), .A3(new_n403), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n874), .B2(new_n867), .ZN(new_n875));
  INV_X1    g0675(.A(new_n873), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n409), .A2(KEYINPUT95), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT95), .B1(new_n409), .B2(new_n876), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT38), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n867), .B1(new_n866), .B2(new_n869), .ZN(new_n881));
  AND4_X1   g0681(.A1(new_n867), .A2(new_n871), .A3(new_n869), .A4(new_n403), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n869), .B1(new_n608), .B2(new_n603), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n880), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n331), .A2(KEYINPUT14), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n335), .A2(new_n337), .A3(G169), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n892), .B(new_n893), .C1(new_n301), .C2(new_n335), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n317), .A3(new_n660), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n608), .A2(new_n868), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n890), .A2(new_n879), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n817), .A2(new_n659), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n819), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n317), .B(new_n659), .C1(new_n894), .C2(new_n601), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n317), .A2(new_n659), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n339), .A2(new_n342), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n898), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n865), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n409), .A2(new_n876), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT95), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n409), .A2(KEYINPUT95), .A3(new_n876), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n915), .B2(new_n875), .ZN(new_n916));
  INV_X1    g0716(.A(new_n879), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n902), .A2(new_n904), .B1(new_n811), .B2(new_n810), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n721), .A2(KEYINPUT98), .A3(new_n659), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT98), .B1(new_n721), .B2(new_n659), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT31), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n707), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n919), .B(new_n920), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n812), .B(new_n905), .C1(new_n923), .C2(new_n925), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n879), .B2(new_n885), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n918), .A2(new_n926), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT31), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n707), .A2(new_n924), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n434), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n927), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n920), .B1(new_n886), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n926), .B1(new_n890), .B2(new_n879), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n434), .A2(new_n932), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(G330), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n910), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n205), .B2(new_n736), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n910), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n862), .B1(new_n942), .B2(new_n943), .ZN(G367));
  NAND2_X1  g0744(.A1(new_n536), .A2(new_n659), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n636), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT99), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n618), .A2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(KEYINPUT99), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n751), .ZN(new_n952));
  INV_X1    g0752(.A(new_n241), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n753), .B1(new_n209), .B2(new_n414), .C1(new_n953), .C2(new_n746), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n739), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n796), .A2(G68), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n762), .B2(new_n356), .C1(new_n759), .C2(new_n830), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n263), .B1(new_n766), .B2(new_n828), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G137), .B2(new_n786), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n779), .A2(G159), .B1(G77), .B2(new_n774), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n760), .C2(new_n784), .ZN(new_n962));
  INV_X1    g0762(.A(G303), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n353), .B1(new_n766), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G317), .B2(new_n786), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n761), .A2(G116), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(new_n842), .C2(new_n784), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n758), .A2(G311), .B1(G107), .B2(new_n796), .ZN(new_n969));
  INV_X1    g0769(.A(G294), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n969), .B1(new_n511), .B2(new_n775), .C1(new_n970), .C2(new_n827), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n958), .A2(new_n962), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT47), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n850), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n956), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n952), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n661), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n671), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n669), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n684), .B1(new_n524), .B2(new_n660), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n629), .A2(new_n659), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT102), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT102), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n670), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n983), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT103), .B1(new_n670), .B2(new_n983), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT44), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  INV_X1    g0797(.A(new_n995), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n983), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n993), .A2(new_n677), .A3(new_n996), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT104), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n676), .B1(new_n668), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n668), .A2(new_n1002), .A3(new_n676), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n671), .A2(new_n978), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1005), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1006), .B1(new_n1009), .B2(new_n1003), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n733), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1000), .A2(new_n991), .A3(new_n996), .A4(new_n992), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n677), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1001), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n733), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n679), .B(KEYINPUT41), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n738), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n983), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n677), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n668), .A2(new_n983), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT42), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n983), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n558), .B1(new_n981), .B2(new_n642), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n660), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT43), .B1(new_n1031), .B2(KEYINPUT100), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(KEYINPUT100), .A3(KEYINPUT43), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n951), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1031), .A2(new_n950), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1033), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1023), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1033), .A2(new_n1037), .A3(new_n1034), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1023), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1040), .A2(new_n1035), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n977), .B1(new_n1021), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT106), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(G387));
  NAND3_X1  g0846(.A1(new_n665), .A2(new_n667), .A3(new_n751), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n742), .A2(new_n680), .B1(G107), .B2(new_n209), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n238), .A2(G45), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n275), .A2(new_n760), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT50), .Z(new_n1051));
  INV_X1    g0851(.A(new_n680), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n1052), .C1(G68), .C2(G77), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n746), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1048), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n739), .B1(new_n1055), .B2(new_n754), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n765), .B1(new_n779), .B2(G311), .ZN(new_n1057));
  INV_X1    g0857(.A(G322), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n759), .C1(new_n784), .C2(new_n963), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n761), .A2(G294), .B1(new_n796), .B2(G283), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n775), .A2(new_n571), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n263), .B(new_n1068), .C1(G326), .C2(new_n786), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n788), .A2(new_n307), .B1(new_n828), .B2(new_n769), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n353), .B(new_n1071), .C1(G50), .C2(new_n765), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n761), .A2(G77), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n779), .A2(new_n275), .B1(new_n415), .B2(new_n796), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n758), .A2(G159), .B1(G97), .B2(new_n774), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1070), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1056), .B1(new_n1077), .B2(new_n752), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1011), .A2(new_n738), .B1(new_n1047), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n706), .A2(new_n732), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n735), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT107), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1082), .A2(new_n1083), .B1(new_n733), .B2(new_n1011), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT107), .B1(new_n1012), .B2(new_n735), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(G393));
  NAND3_X1  g0886(.A1(new_n1001), .A2(new_n1016), .A3(new_n738), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n753), .B1(new_n511), .B2(new_n209), .C1(new_n248), .C2(new_n746), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n739), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n263), .B1(new_n830), .B2(new_n769), .C1(new_n775), .C2(new_n528), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n833), .B2(new_n275), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n777), .A2(new_n266), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n779), .B2(G50), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n307), .C2(new_n762), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n765), .A2(G159), .B1(new_n758), .B2(G150), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(KEYINPUT109), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(KEYINPUT109), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n765), .A2(G311), .B1(new_n758), .B2(G317), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT52), .Z(new_n1102));
  OAI21_X1  g0902(.A(new_n353), .B1(new_n769), .B2(new_n1058), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n781), .B2(G294), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n762), .A2(new_n842), .B1(new_n571), .B2(new_n777), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n776), .B(new_n1105), .C1(G303), .C2(new_n779), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1099), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1089), .B1(new_n1108), .B2(new_n752), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n983), .B2(new_n802), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1017), .A2(new_n735), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1013), .B1(new_n1001), .B2(new_n1016), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1087), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(G390));
  NAND3_X1  g0913(.A1(new_n932), .A2(G330), .A3(new_n919), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n886), .A2(new_n895), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n812), .B1(new_n696), .B2(new_n697), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n900), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n905), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n819), .A2(new_n900), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n896), .B1(new_n1120), .B2(new_n905), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n888), .B2(new_n891), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1115), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1116), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n900), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n695), .A2(new_n660), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT90), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n660), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1125), .B1(new_n1130), .B2(new_n812), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1124), .B1(new_n1131), .B2(new_n906), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n888), .A2(new_n891), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1121), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n812), .C1(new_n725), .C2(new_n731), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1136), .A2(new_n906), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1123), .A2(new_n1138), .A3(new_n738), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n749), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n739), .B1(new_n275), .B2(new_n824), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n766), .A2(new_n837), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n353), .B(new_n1142), .C1(G125), .C2(new_n786), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n827), .A2(new_n831), .B1(new_n777), .B2(new_n770), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n759), .A2(new_n1145), .B1(new_n760), .B2(new_n775), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n833), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n761), .A2(G150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT53), .Z(new_n1152));
  NAND4_X1  g0952(.A1(new_n1143), .A2(new_n1147), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n422), .A2(new_n827), .B1(new_n759), .B2(new_n842), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n833), .B2(G97), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT113), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n353), .B1(new_n769), .B2(new_n970), .C1(new_n766), .C2(new_n571), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n762), .A2(new_n528), .B1(new_n775), .B2(new_n307), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1157), .A2(new_n1092), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1153), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT114), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n850), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1141), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1140), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1139), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1123), .A2(new_n1138), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n814), .A2(new_n815), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(G330), .C1(new_n923), .C2(new_n925), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT111), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n906), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT111), .B1(new_n1173), .B2(new_n905), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1131), .A2(new_n1137), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT110), .ZN(new_n1176));
  INV_X1    g0976(.A(G330), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n930), .B2(new_n931), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1178), .A2(new_n919), .B1(new_n1136), .B2(new_n906), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1176), .B1(new_n1179), .B2(new_n901), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1136), .A2(new_n906), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1114), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(KEYINPUT110), .A3(new_n1120), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1175), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n434), .A2(new_n1178), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n863), .A2(new_n611), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n679), .B1(new_n1168), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT112), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1187), .B1(new_n1175), .B2(new_n1184), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1138), .A3(new_n1123), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1191), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1167), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT115), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1168), .A2(new_n1189), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n735), .A3(new_n1193), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT112), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1166), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT115), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1197), .A2(new_n1204), .ZN(G378));
  NAND2_X1  g1005(.A1(new_n1193), .A2(new_n1188), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n897), .A2(new_n908), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n292), .A2(new_n872), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT55), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n299), .A2(new_n305), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1211), .B1(new_n299), .B2(new_n305), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1209), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n1208), .A3(new_n1212), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n929), .B2(G330), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G330), .B(new_n1218), .C1(new_n935), .C2(new_n936), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1207), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT119), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1218), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n937), .B2(new_n1177), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n909), .A3(new_n1220), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n909), .A3(KEYINPUT119), .A4(new_n1220), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1206), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n679), .B1(new_n1232), .B2(new_n1206), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1227), .A2(new_n738), .A3(new_n1228), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n738), .B(new_n735), .C1(new_n760), .C2(new_n823), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n759), .A2(new_n571), .B1(new_n356), .B2(new_n775), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G97), .B2(new_n779), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n422), .A2(new_n766), .B1(new_n788), .B2(new_n414), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n318), .B(new_n353), .C1(new_n842), .C2(new_n769), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1241), .A3(new_n957), .A4(new_n1073), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT58), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n760), .B1(G33), .B2(G41), .C1(new_n256), .C2(new_n263), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1145), .A2(new_n766), .B1(new_n788), .B2(new_n831), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G125), .A2(new_n758), .B1(new_n779), .B2(G132), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n828), .B2(new_n777), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(new_n761), .C2(new_n1149), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT116), .Z(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT117), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(G124), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(G124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n786), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G33), .A2(G41), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n770), .C2(new_n775), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1252), .B2(KEYINPUT59), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1244), .B(new_n1247), .C1(new_n1253), .C2(new_n1260), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1236), .B1(new_n850), .B2(new_n1261), .C1(new_n1218), .C2(new_n750), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1235), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1234), .A2(new_n1264), .ZN(G375));
  NOR2_X1   g1065(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT120), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT120), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1020), .A3(new_n1189), .A4(new_n1269), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(KEYINPUT121), .Z(new_n1271));
  NOR2_X1   g1071(.A1(new_n905), .A2(new_n750), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT122), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n833), .A2(G107), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n759), .A2(new_n970), .B1(new_n511), .B2(new_n762), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G116), .B2(new_n779), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n353), .B1(new_n769), .B2(new_n963), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n765), .B2(G283), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n796), .A2(new_n415), .B1(new_n774), .B2(G77), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1276), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n781), .A2(G150), .B1(G128), .B2(new_n786), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n353), .B1(new_n765), .B2(G137), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n779), .A2(new_n1149), .B1(G58), .B2(new_n774), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n761), .A2(G159), .B1(new_n796), .B2(G50), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n758), .A2(G132), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT123), .Z(new_n1287));
  OAI21_X1  g1087(.A(new_n1280), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n850), .B1(new_n1288), .B2(KEYINPUT124), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(KEYINPUT124), .B2(new_n1288), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n823), .A2(new_n307), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1273), .A2(new_n739), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1175), .A2(new_n1184), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n737), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1271), .A2(new_n1295), .ZN(G381));
  OAI211_X1 g1096(.A(new_n804), .B(new_n1079), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G381), .A2(G384), .A3(G390), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1045), .A2(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1299), .A2(KEYINPUT125), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(KEYINPUT125), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1199), .A2(new_n1167), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(G375), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1301), .A3(new_n1303), .ZN(G407));
  INV_X1    g1104(.A(G213), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1303), .B2(new_n658), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G407), .A2(new_n1306), .ZN(G409));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1305), .A2(G343), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G375), .B1(new_n1204), .B2(new_n1197), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1229), .A2(new_n1019), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1262), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1314), .B2(new_n738), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1302), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(KEYINPUT126), .B(new_n1310), .C1(new_n1311), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1268), .A2(new_n1269), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n679), .B1(new_n1266), .B2(KEYINPUT60), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1295), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n852), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(G384), .A3(new_n1295), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1309), .A2(G2897), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1325), .B(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1317), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1263), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1330));
  AOI211_X1 g1130(.A(KEYINPUT115), .B(new_n1166), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1329), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1316), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT126), .B1(new_n1334), .B2(new_n1310), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1308), .B1(new_n1328), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1316), .B1(G378), .B2(new_n1329), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1337), .B1(new_n1338), .B2(new_n1309), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1339), .A2(KEYINPUT127), .A3(new_n1327), .A4(new_n1317), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1325), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1341), .B(new_n1310), .C1(new_n1311), .C2(new_n1316), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  OR2_X1    g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n737), .ZN(new_n1346));
  OR2_X1    g1146(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1347));
  AOI22_X1  g1147(.A1(new_n1346), .A2(new_n1347), .B1(new_n952), .B2(new_n976), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G393), .A2(G396), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1297), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT106), .ZN(new_n1351));
  AOI21_X1  g1151(.A(G390), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1112), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(new_n735), .A3(new_n1017), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1087), .A2(new_n1110), .ZN(new_n1355));
  AOI22_X1  g1155(.A1(new_n1354), .A2(new_n1355), .B1(new_n1349), .B2(new_n1297), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1348), .B1(new_n1352), .B2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1350), .A2(G390), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT106), .B1(new_n1349), .B2(new_n1297), .ZN(new_n1359));
  OAI211_X1 g1159(.A(new_n1358), .B(new_n1044), .C1(G390), .C2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT61), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1357), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1362), .B1(new_n1343), .B2(new_n1342), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1336), .A2(new_n1340), .A3(new_n1344), .A4(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1357), .A2(new_n1360), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1342), .A2(KEYINPUT62), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1327), .B1(new_n1338), .B2(new_n1309), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1366), .A2(new_n1367), .A3(new_n1361), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1342), .A2(KEYINPUT62), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1365), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1364), .A2(new_n1370), .ZN(G405));
  NAND3_X1  g1171(.A1(G375), .A2(new_n1167), .A3(new_n1199), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1332), .A2(new_n1372), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1373), .B(new_n1341), .ZN(new_n1374));
  XNOR2_X1  g1174(.A(new_n1374), .B(new_n1365), .ZN(G402));
endmodule


