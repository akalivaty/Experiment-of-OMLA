//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G101), .A3(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n472), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(G160));
  NAND4_X1  g057(.A1(new_n466), .A2(new_n468), .A3(G2105), .A4(new_n469), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n479), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n470), .B2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  OAI221_X1 g067(.A(new_n485), .B1(new_n486), .B2(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n479), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n483), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n479), .A2(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n475), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n466), .A2(new_n468), .A3(new_n502), .A4(new_n469), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n507));
  AOI211_X1 g082(.A(KEYINPUT71), .B(new_n498), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  INV_X1    g085(.A(new_n500), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n498), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n508), .A2(new_n514), .ZN(G164));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT6), .B1(KEYINPUT72), .B2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n524), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  INV_X1    g104(.A(new_n520), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n533), .B(new_n534), .C1(new_n522), .C2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT5), .B(G543), .Z(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n526), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n543), .B1(new_n542), .B2(new_n541), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n519), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n517), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n530), .A2(G90), .B1(G52), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n547), .A2(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI221_X1 g128(.A(new_n551), .B1(new_n552), .B2(new_n526), .C1(new_n553), .C2(new_n520), .ZN(new_n554));
  INV_X1    g129(.A(G860), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n554), .A2(new_n555), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(KEYINPUT74), .A2(G53), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n522), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n522), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n539), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n530), .A2(G91), .B1(new_n567), .B2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  XNOR2_X1  g145(.A(G168), .B(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G286));
  NAND2_X1  g147(.A1(new_n530), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n547), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n547), .A2(G48), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  OAI221_X1 g154(.A(new_n577), .B1(new_n520), .B2(new_n578), .C1(new_n526), .C2(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT76), .ZN(G305));
  AOI22_X1  g156(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n582), .A2(new_n583), .A3(new_n526), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT78), .B(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n530), .A2(new_n585), .B1(G47), .B2(new_n547), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n583), .B1(new_n582), .B2(new_n526), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n520), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n547), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n600), .A2(G54), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n539), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n598), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n598), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n597), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n593), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n593), .B1(new_n610), .B2(G868), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n571), .B2(G868), .ZN(G297));
  XNOR2_X1  g189(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g190(.A(new_n597), .ZN(new_n616));
  INV_X1    g191(.A(new_n609), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n607), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(G559), .B2(new_n555), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT83), .ZN(G148));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n554), .B(new_n622), .S(G868), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n484), .A2(G123), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT86), .Z(new_n626));
  INV_X1    g201(.A(new_n491), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G135), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n479), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(G2100), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n636), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n638), .B2(new_n637), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n640), .B1(new_n642), .B2(new_n639), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n632), .A2(new_n633), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT88), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT18), .ZN(new_n669));
  OAI21_X1  g244(.A(KEYINPUT17), .B1(new_n660), .B2(new_n661), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(new_n663), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n663), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n662), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT20), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT89), .Z(new_n686));
  NOR3_X1   g261(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G32), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n627), .A2(G141), .ZN(new_n699));
  INV_X1    g274(.A(G105), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n700), .A2(new_n465), .A3(G2105), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT26), .ZN(new_n703));
  AOI211_X1 g278(.A(new_n701), .B(new_n703), .C1(new_n484), .C2(G129), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(new_n697), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G29), .A2(G35), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G162), .B2(G29), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT29), .B(G2090), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n708), .B(new_n713), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(G20), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT98), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G299), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1956), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  NAND2_X1  g299(.A1(G160), .A2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n726), .B2(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(KEYINPUT24), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n718), .B(new_n723), .C1(new_n724), .C2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n717), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n724), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT97), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n610), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G4), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1348), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n733), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n697), .A2(G27), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G164), .B2(new_n697), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2078), .ZN(new_n742));
  NAND2_X1  g317(.A1(G115), .A2(G2104), .ZN(new_n743));
  INV_X1    g318(.A(G127), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n475), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT25), .ZN(new_n746));
  NAND2_X1  g321(.A1(G103), .A2(G2104), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G2105), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n479), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n745), .A2(G2105), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G139), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n491), .B2(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G33), .B(new_n752), .S(G29), .Z(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G2072), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n709), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n709), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G1966), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(G1966), .ZN(new_n758));
  MUX2_X1   g333(.A(G19), .B(new_n554), .S(G16), .Z(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT94), .B(G1341), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n697), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n627), .A2(G140), .ZN(new_n765));
  NOR2_X1   g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT95), .ZN(new_n767));
  INV_X1    g342(.A(G116), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n465), .B1(new_n768), .B2(G2105), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n484), .A2(G128), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n631), .A2(new_n697), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n759), .A2(new_n761), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT96), .B(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(KEYINPUT30), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n754), .A2(new_n762), .A3(new_n773), .A4(new_n781), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n731), .A2(new_n739), .A3(new_n742), .A4(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT99), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n709), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n709), .ZN(new_n786));
  INV_X1    g361(.A(G1971), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n709), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(G288), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n709), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT33), .B(G1976), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n709), .A2(G6), .ZN(new_n797));
  INV_X1    g372(.A(G305), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n709), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n788), .B(new_n793), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n796), .B2(new_n799), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n484), .A2(G119), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n479), .A2(G107), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(G131), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n803), .B1(new_n804), .B2(new_n805), .C1(new_n491), .C2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G25), .B(new_n807), .S(G29), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT35), .B(G1991), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G24), .B(G290), .S(G16), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT92), .ZN(new_n813));
  INV_X1    g388(.A(G1986), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n802), .B(new_n815), .C1(new_n814), .C2(new_n813), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n784), .A2(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  XOR2_X1   g394(.A(KEYINPUT100), .B(G93), .Z(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n520), .A2(new_n820), .B1(new_n522), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT101), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n526), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NOR2_X1   g402(.A1(new_n618), .A2(new_n621), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT102), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n825), .B(new_n554), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n555), .B1(new_n833), .B2(KEYINPUT39), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n827), .B1(new_n834), .B2(new_n835), .ZN(G145));
  XNOR2_X1  g411(.A(new_n705), .B(new_n752), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n484), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n479), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(G142), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n838), .B1(new_n839), .B2(new_n840), .C1(new_n491), .C2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(new_n635), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n837), .B(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n771), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n807), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n844), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(G162), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n631), .ZN(new_n851));
  AOI21_X1  g426(.A(G37), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n849), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g429(.A(G868), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n825), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G290), .B(new_n798), .ZN(new_n857));
  XNOR2_X1  g432(.A(G303), .B(G288), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(KEYINPUT42), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n862), .B(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n831), .B(new_n622), .Z(new_n867));
  INV_X1    g442(.A(G299), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT103), .B1(new_n618), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n610), .A2(new_n870), .A3(G299), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n618), .A2(new_n868), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n869), .B2(new_n871), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n873), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n610), .A2(KEYINPUT104), .A3(G299), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n618), .B2(new_n868), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(new_n882), .B2(new_n872), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n875), .B1(new_n888), .B2(new_n867), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n866), .B1(KEYINPUT107), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(KEYINPUT107), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(new_n866), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n856), .B1(new_n892), .B2(new_n855), .ZN(G295));
  OAI21_X1  g468(.A(new_n856), .B1(new_n892), .B2(new_n855), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  INV_X1    g472(.A(G168), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(G171), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(G301), .A2(KEYINPUT108), .A3(G168), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n899), .B(new_n900), .C1(new_n571), .C2(G301), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(new_n831), .Z(new_n902));
  INV_X1    g477(.A(new_n887), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n885), .ZN(new_n904));
  INV_X1    g479(.A(new_n863), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n902), .A2(new_n874), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n863), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n896), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n901), .B(new_n831), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n872), .B2(new_n873), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n914), .A2(new_n915), .B1(new_n882), .B2(new_n877), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n874), .B2(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n902), .A2(new_n874), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n863), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n907), .A2(new_n920), .A3(new_n908), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n895), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n895), .B1(new_n921), .B2(KEYINPUT43), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n911), .A2(new_n896), .A3(new_n908), .A4(new_n907), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(G397));
  AOI21_X1  g504(.A(G1384), .B1(new_n512), .B2(new_n513), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(KEYINPUT45), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n472), .A2(new_n478), .A3(G40), .A4(new_n480), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n705), .B(G1996), .ZN(new_n935));
  INV_X1    g510(.A(G2067), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n771), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n938), .A2(new_n810), .A3(new_n807), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n765), .A2(new_n936), .A3(new_n770), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n938), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n807), .B(new_n809), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n934), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n934), .A2(G290), .A3(G1986), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n944), .A2(new_n945), .B1(KEYINPUT48), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(KEYINPUT48), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n934), .B2(G1996), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT126), .Z(new_n953));
  NOR3_X1   g528(.A1(new_n934), .A2(new_n951), .A3(G1996), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT127), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n937), .A2(new_n705), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n953), .B(new_n955), .C1(new_n934), .C2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n950), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n950), .B2(new_n957), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(G1384), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n933), .B1(new_n845), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT70), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(new_n966), .A3(new_n500), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT71), .B1(new_n967), .B2(new_n498), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n512), .A2(new_n509), .A3(new_n513), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n508), .B2(new_n514), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n960), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(KEYINPUT111), .A3(new_n964), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n787), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G2090), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n932), .B1(new_n930), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n979), .B(new_n981), .C1(new_n970), .C2(new_n980), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n985), .A2(KEYINPUT112), .A3(new_n979), .A4(new_n981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(G166), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n994));
  NAND3_X1  g569(.A1(G303), .A2(G8), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n978), .A2(new_n987), .A3(KEYINPUT113), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n990), .A2(G8), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n930), .A2(new_n933), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(G1976), .B2(new_n790), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n580), .B(G1981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1009));
  MUX2_X1   g584(.A(new_n1008), .B(new_n1006), .S(new_n1009), .Z(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n1002), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(G288), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1005), .B(new_n1011), .C1(new_n1003), .C2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1012), .B(new_n790), .C1(new_n1010), .C2(new_n1002), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n580), .A2(G1981), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(new_n1002), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(KEYINPUT116), .A3(new_n1016), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1000), .A2(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n933), .B1(new_n930), .B2(KEYINPUT45), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n961), .B1(new_n508), .B2(new_n514), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT118), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1966), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n724), .B(new_n981), .C1(new_n970), .C2(new_n980), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1021), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1966), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n974), .B1(new_n967), .B2(new_n498), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n932), .B1(new_n1033), .B2(new_n960), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1023), .A2(KEYINPUT118), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT124), .A3(new_n1029), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(G168), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(new_n992), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G168), .A2(new_n992), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n1040), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1037), .A2(new_n1029), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT111), .B1(new_n976), .B2(new_n964), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n972), .B(new_n963), .C1(new_n975), .C2(new_n960), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1056), .B2(G2078), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1053), .A2(G2078), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n981), .B1(new_n970), .B2(new_n980), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(new_n1059), .B1(new_n712), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(G301), .B(KEYINPUT54), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n712), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1034), .B(new_n1059), .C1(new_n845), .C2(new_n962), .ZN(new_n1065));
  XOR2_X1   g640(.A(new_n1065), .B(KEYINPUT125), .Z(new_n1066));
  AND3_X1   g641(.A1(new_n1057), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(new_n1062), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n980), .B(new_n974), .C1(new_n508), .C2(new_n514), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n932), .B1(new_n1033), .B2(KEYINPUT50), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT57), .B1(new_n868), .B2(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(G299), .B2(KEYINPUT120), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(KEYINPUT57), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n964), .B(new_n1082), .C1(new_n970), .C2(KEYINPUT45), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1074), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1001), .A2(G2067), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n1060), .B2(new_n736), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n618), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1081), .B1(new_n1074), .B2(new_n1083), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1069), .B(new_n1084), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT122), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1074), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n1088), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1086), .A2(KEYINPUT60), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1348), .B1(new_n985), .B2(new_n981), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1085), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1098), .A3(new_n610), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1082), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1100), .B(new_n963), .C1(new_n975), .C2(new_n960), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1956), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1079), .B(new_n1080), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(KEYINPUT61), .A3(new_n1084), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1094), .A2(new_n1099), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1001), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT58), .B(G1341), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n971), .A2(G1996), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n554), .A2(KEYINPUT123), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1111), .A2(new_n1112), .B1(new_n610), .B2(new_n1095), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1089), .B(new_n1091), .C1(new_n1105), .C2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1052), .A2(new_n1068), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1072), .A2(G2090), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1056), .B2(new_n787), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT117), .B(new_n996), .C1(new_n1117), .C2(new_n992), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1116), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n992), .B1(new_n978), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1121), .B2(new_n997), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(new_n999), .A3(new_n1014), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1020), .B1(new_n1115), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1049), .A2(new_n1126), .A3(new_n1051), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1047), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT62), .B1(new_n1128), .B2(new_n1050), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G301), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1123), .A2(new_n999), .A3(new_n1014), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1134), .A2(new_n992), .A3(G286), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n999), .A3(new_n1014), .A4(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n999), .A2(new_n1014), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(KEYINPUT63), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n990), .A2(G8), .A3(new_n998), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(new_n996), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1125), .A2(new_n1133), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n944), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G290), .B(new_n814), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n934), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n959), .B1(new_n1143), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g722(.A1(new_n912), .A2(new_n922), .ZN(new_n1149));
  NOR4_X1   g723(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n1150), .A2(new_n853), .ZN(new_n1151));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1151), .ZN(G308));
  OR2_X1    g726(.A1(new_n1149), .A2(new_n1151), .ZN(G225));
endmodule


