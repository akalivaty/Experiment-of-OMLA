//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g027(.A1(G221), .A2(G219), .A3(G220), .A4(G218), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(KEYINPUT70), .A3(G125), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n465), .B2(G125), .ZN(new_n473));
  INV_X1    g048(.A(G113), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n467), .ZN(new_n475));
  INV_X1    g050(.A(new_n464), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(G160));
  XOR2_X1   g052(.A(KEYINPUT3), .B(G2104), .Z(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n467), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n483), .B1(new_n482), .B2(new_n481), .C1(new_n464), .C2(G112), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n478), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n461), .A2(new_n463), .A3(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n495), .A3(G138), .A4(new_n465), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT73), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n507), .A2(new_n509), .A3(new_n514), .A4(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n505), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n501), .B1(new_n513), .B2(new_n515), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G88), .B1(new_n517), .B2(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n505), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  XOR2_X1   g101(.A(KEYINPUT76), .B(G89), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT75), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n532), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n531), .A2(new_n529), .A3(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n505), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n528), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT77), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n537), .B1(G51), .B2(new_n517), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(new_n543), .A3(new_n528), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n516), .A2(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n517), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n505), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(new_n523), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n505), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n516), .A2(G81), .B1(new_n556), .B2(new_n523), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n517), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G53), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n513), .B2(new_n515), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI211_X1 g144(.A(KEYINPUT78), .B(new_n566), .C1(new_n513), .C2(new_n515), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT79), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(new_n566), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n511), .B1(new_n522), .B2(KEYINPUT6), .ZN(new_n574));
  AND4_X1   g149(.A1(new_n514), .A2(new_n507), .A3(new_n509), .A4(KEYINPUT6), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n567), .B2(new_n572), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n574), .A2(new_n575), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT78), .B1(new_n581), .B2(new_n566), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n567), .A2(new_n568), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(KEYINPUT9), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n571), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G65), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n505), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n516), .A2(G91), .B1(new_n589), .B2(G651), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT81), .B1(new_n586), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(G299));
  INV_X1    g168(.A(G168), .ZN(G286));
  NAND2_X1  g169(.A1(new_n516), .A2(G87), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n517), .A2(G49), .ZN(new_n596));
  INV_X1    g171(.A(new_n505), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n597), .B2(G74), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(G288));
  OAI211_X1 g174(.A(G48), .B(G543), .C1(new_n574), .C2(new_n575), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g176(.A1(G73), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n505), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n516), .A2(G86), .B1(new_n604), .B2(new_n523), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n516), .A2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n517), .A2(G47), .ZN(new_n608));
  NAND2_X1  g183(.A1(G72), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G60), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n505), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n523), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n516), .A2(G92), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT10), .Z(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n505), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(G651), .A2(new_n619), .B1(new_n517), .B2(G54), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n614), .B1(new_n621), .B2(G868), .ZN(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NOR2_X1   g199(.A1(G168), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(new_n626));
  INV_X1    g201(.A(G299), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n621), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n559), .A2(new_n624), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n616), .A2(new_n620), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(new_n624), .ZN(G323));
  XOR2_X1   g210(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n636));
  XNOR2_X1  g211(.A(G323), .B(new_n636), .ZN(G282));
  AOI22_X1  g212(.A1(G123), .A2(new_n479), .B1(new_n485), .B2(G135), .ZN(new_n638));
  OAI221_X1 g213(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n465), .A2(new_n468), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT85), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n665), .B(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n674), .B2(new_n671), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n671), .A3(new_n668), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n670), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  INV_X1    g262(.A(new_n682), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n687), .B(new_n691), .C1(new_n688), .C2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT33), .Z(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(G1976), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(G1976), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n699), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n699), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n704), .A2(new_n707), .A3(new_n708), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n479), .A2(G119), .ZN(new_n719));
  OAI221_X1 g294(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n485), .A2(G131), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n699), .A2(G24), .ZN(new_n727));
  INV_X1    g302(.A(G290), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n699), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT88), .B(G1986), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n715), .A2(new_n716), .A3(new_n726), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT36), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n699), .A2(G20), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT23), .Z(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G299), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1956), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n717), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n479), .A2(G129), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n485), .A2(G141), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n468), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NAND4_X1  g321(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n717), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n717), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n741), .B1(new_n717), .B2(new_n640), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  OR2_X1    g328(.A1(G29), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT91), .Z(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT25), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT25), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  INV_X1    g334(.A(G127), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n478), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n761), .A2(new_n476), .B1(new_n485), .B2(G139), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n757), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n754), .B1(new_n763), .B2(new_n717), .ZN(new_n764));
  INV_X1    g339(.A(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT24), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G160), .B2(new_n717), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G2084), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n717), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n717), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT29), .Z(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n753), .A2(new_n766), .A3(new_n772), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G171), .A2(new_n699), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G5), .B2(new_n699), .ZN(new_n780));
  INV_X1    g355(.A(G1961), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n717), .A2(G27), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n717), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G2078), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n780), .A2(new_n781), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n717), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AOI22_X1  g364(.A1(G128), .A2(new_n479), .B1(new_n485), .B2(G140), .ZN(new_n790));
  OAI221_X1 g365(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n782), .A2(new_n785), .A3(new_n786), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n775), .A2(new_n776), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n764), .A2(new_n765), .B1(G2084), .B2(new_n771), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n778), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT92), .B1(G16), .B2(G21), .ZN(new_n799));
  NAND2_X1  g374(.A1(G168), .A2(G16), .ZN(new_n800));
  MUX2_X1   g375(.A(KEYINPUT92), .B(new_n799), .S(new_n800), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1966), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G19), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n560), .B2(G16), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1341), .Z(new_n805));
  NOR2_X1   g380(.A1(new_n621), .A2(new_n699), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G4), .B2(new_n699), .ZN(new_n807));
  INV_X1    g382(.A(G1348), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  AND4_X1   g385(.A1(new_n737), .A2(new_n798), .A3(new_n802), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n733), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT93), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(G311));
  XNOR2_X1  g389(.A(new_n812), .B(KEYINPUT94), .ZN(G150));
  NAND2_X1  g390(.A1(new_n516), .A2(G93), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n505), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n523), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT95), .B(G55), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n517), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n816), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NOR2_X1   g400(.A1(new_n633), .A2(new_n630), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n559), .A2(new_n823), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n516), .A2(G93), .B1(new_n819), .B2(new_n523), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n557), .A2(new_n829), .A3(new_n558), .A4(new_n822), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n827), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT96), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n833), .B2(new_n834), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n825), .B1(new_n836), .B2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(G160), .B(KEYINPUT97), .ZN(new_n840));
  XNOR2_X1  g415(.A(G162), .B(new_n640), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n722), .B(KEYINPUT99), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n643), .ZN(new_n844));
  AOI22_X1  g419(.A1(G130), .A2(new_n479), .B1(new_n485), .B2(G142), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n844), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n494), .A2(new_n496), .ZN(new_n849));
  INV_X1    g424(.A(new_n492), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n792), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n747), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n848), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n848), .A2(new_n857), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n842), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(G37), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n859), .A2(KEYINPUT100), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(KEYINPUT100), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n858), .A4(new_n842), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(G395));
  XOR2_X1   g443(.A(new_n831), .B(KEYINPUT102), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n634), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n633), .B1(new_n591), .B2(new_n592), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n586), .A2(new_n590), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT81), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n590), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n621), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT41), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n871), .B2(new_n876), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n878), .B1(new_n870), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(G303), .B(G288), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(G305), .A2(new_n728), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n601), .A2(new_n605), .A3(G290), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT103), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n883), .A2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(G868), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n823), .A2(new_n624), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(G295));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(G331));
  INV_X1    g473(.A(new_n891), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n543), .B1(new_n542), .B2(new_n528), .ZN(new_n900));
  AND4_X1   g475(.A1(new_n543), .A2(new_n528), .A3(new_n538), .A4(new_n539), .ZN(new_n901));
  OAI21_X1  g476(.A(G301), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n541), .A2(new_n544), .A3(G171), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n831), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n902), .A2(new_n831), .A3(new_n906), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n832), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n877), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT41), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n904), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n877), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n899), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n879), .B2(new_n880), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n899), .B1(new_n910), .B2(new_n877), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n916), .B1(new_n912), .B2(new_n913), .ZN(new_n926));
  INV_X1    g501(.A(new_n877), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n899), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n930), .B2(new_n922), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n922), .A3(new_n925), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n930), .A2(new_n922), .A3(KEYINPUT106), .A4(new_n925), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n925), .B1(new_n923), .B2(KEYINPUT107), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n919), .A2(new_n922), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n891), .B1(new_n927), .B2(new_n928), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n926), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n928), .B1(new_n879), .B2(new_n880), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n891), .B1(new_n950), .B2(new_n917), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT107), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AND4_X1   g527(.A1(KEYINPUT108), .A2(new_n952), .A3(KEYINPUT43), .A4(new_n945), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n936), .B(new_n942), .C1(new_n946), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n945), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n952), .A2(new_n945), .A3(KEYINPUT108), .A4(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n936), .B1(new_n960), .B2(new_n942), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n935), .B1(new_n955), .B2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  NAND3_X1  g538(.A1(G160), .A2(new_n963), .A3(G40), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n466), .A2(new_n469), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n474), .A2(new_n467), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT70), .ZN(new_n967));
  INV_X1    g542(.A(G125), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n478), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(new_n471), .ZN(new_n970));
  OAI211_X1 g545(.A(G40), .B(new_n965), .C1(new_n970), .C2(new_n464), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(G1384), .ZN(new_n974));
  NOR2_X1   g549(.A1(G164), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT45), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n748), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n792), .A2(G2067), .ZN(new_n983));
  INV_X1    g558(.A(G2067), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n790), .A2(new_n984), .A3(new_n791), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n979), .B2(new_n748), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n982), .A2(new_n725), .A3(new_n723), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n989), .B2(new_n985), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n981), .B(KEYINPUT46), .Z(new_n991));
  INV_X1    g566(.A(new_n986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n977), .B1(new_n747), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n722), .B(new_n725), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n982), .B(new_n988), .C1(new_n978), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n990), .B(new_n996), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT45), .B1(new_n851), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NOR3_X1   g583(.A1(G164), .A2(new_n1008), .A3(new_n974), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n973), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n711), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n851), .A2(new_n1005), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n964), .A2(new_n972), .B1(KEYINPUT50), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n776), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1004), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(KEYINPUT113), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1013), .B1(new_n964), .B2(new_n972), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n1004), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G288), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1025), .B(new_n1030), .C1(new_n1027), .C2(G288), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  INV_X1    g607(.A(G1981), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n601), .A2(new_n1033), .A3(new_n605), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1034), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1025), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1023), .A2(new_n1029), .A3(new_n1031), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1017), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1022), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1017), .A2(new_n1042), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1966), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1013), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT45), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1006), .B1(new_n964), .B2(new_n972), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT116), .B(new_n1006), .C1(new_n964), .C2(new_n972), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n963), .B1(G160), .B2(G40), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1015), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1058), .A2(G2084), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1004), .B(G286), .C1(new_n1054), .C2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1041), .A2(new_n1046), .A3(KEYINPUT63), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1060), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1015), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1014), .A2(KEYINPUT115), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n776), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1004), .B1(new_n1068), .B2(new_n1012), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(new_n1022), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1062), .A2(new_n1070), .A3(new_n1040), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1061), .B1(new_n1071), .B2(KEYINPUT63), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1029), .A2(new_n1031), .A3(new_n1039), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n1023), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1039), .A2(new_n1027), .A3(new_n701), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1034), .B(KEYINPUT114), .Z(new_n1076));
  AOI21_X1  g651(.A(new_n1026), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1956), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1015), .B1(new_n1014), .B2(KEYINPUT115), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1050), .A2(new_n1010), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n872), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n586), .A2(KEYINPUT57), .A3(new_n590), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1956), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1095), .B2(new_n1086), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT61), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT120), .B(new_n1093), .C1(new_n1095), .C2(new_n1086), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1006), .B(new_n1009), .C1(new_n964), .C2(new_n972), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n973), .A2(new_n1048), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  AOI22_X1  g678(.A1(new_n1101), .A2(new_n979), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT59), .B1(new_n1104), .B2(new_n559), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1011), .A2(G1996), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1106), .B(new_n560), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1058), .A2(new_n808), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1024), .A2(new_n984), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1111), .A2(new_n633), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n633), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1084), .A2(new_n1116), .A3(new_n1092), .A4(new_n1087), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n633), .A2(KEYINPUT60), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1118), .A3(new_n1112), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1110), .A2(new_n1115), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1093), .A2(KEYINPUT119), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1092), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1088), .A2(new_n1121), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n1067), .A3(new_n1015), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1086), .B1(new_n1127), .B2(new_n1081), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1114), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1100), .A2(new_n1120), .B1(new_n1130), .B2(new_n1094), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1011), .B2(G2078), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1058), .A2(new_n781), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(G2078), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(G301), .B(KEYINPUT54), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n965), .A2(G40), .A3(new_n1137), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1009), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n464), .B1(new_n475), .B2(KEYINPUT122), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(KEYINPUT122), .B2(new_n475), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1142), .B(new_n1144), .C1(KEYINPUT45), .C2(new_n975), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1145), .B2(KEYINPUT123), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(KEYINPUT123), .B2(new_n1145), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1138), .A2(new_n1140), .B1(new_n1135), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1054), .A2(G168), .A3(new_n1059), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT51), .ZN(new_n1151));
  AOI21_X1  g726(.A(G168), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(KEYINPUT51), .ZN(new_n1154));
  OAI211_X1 g729(.A(G8), .B(new_n1149), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1148), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1138), .A2(G301), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(KEYINPUT62), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1151), .A2(new_n1161), .A3(new_n1155), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1131), .A2(new_n1156), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1041), .B(KEYINPUT124), .C1(new_n1069), .C2(new_n1022), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1070), .B2(new_n1040), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1080), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(G290), .B(G1986), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n998), .B1(new_n977), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT125), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1097), .B1(new_n1128), .B2(new_n1092), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(new_n1116), .A3(new_n1099), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1094), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1120), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1088), .A2(new_n1121), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n1129), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1114), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1094), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1156), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1159), .A2(KEYINPUT62), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1182), .A2(new_n1162), .A3(new_n1157), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1167), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT125), .B(new_n1170), .C1(new_n1184), .C2(new_n1079), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1003), .B1(new_n1171), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  OR3_X1    g763(.A1(G401), .A2(new_n1189), .A3(G227), .ZN(new_n1190));
  NOR4_X1   g764(.A1(new_n866), .A2(G229), .A3(new_n932), .A4(new_n1190), .ZN(G308));
  NOR3_X1   g765(.A1(new_n866), .A2(G229), .A3(new_n1190), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1192), .A2(new_n933), .ZN(G225));
endmodule


