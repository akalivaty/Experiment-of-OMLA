//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(G104), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT90), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT90), .A2(G143), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT90), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(G237), .A2(G953), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(G214), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(G131), .B1(new_n194), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n189), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n198), .A2(G214), .B1(KEYINPUT90), .B2(G143), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n201), .B(new_n202), .C1(new_n203), .C2(new_n189), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT94), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(KEYINPUT74), .A3(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(G125), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT74), .B1(new_n211), .B2(G125), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n205), .A2(new_n206), .B1(new_n217), .B2(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(KEYINPUT74), .A3(G125), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n207), .B2(G140), .ZN(new_n221));
  OAI211_X1 g035(.A(KEYINPUT92), .B(new_n219), .C1(new_n221), .C2(new_n208), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n213), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT92), .B1(new_n224), .B2(new_n219), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT19), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n211), .A2(G125), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n208), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n207), .A2(G140), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n231), .A3(KEYINPUT75), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n200), .A2(KEYINPUT94), .A3(new_n204), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(G146), .B1(new_n223), .B2(new_n225), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT76), .B1(new_n233), .B2(new_n227), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT76), .ZN(new_n241));
  AOI211_X1 g055(.A(new_n241), .B(G146), .C1(new_n230), .C2(new_n232), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT18), .A2(G131), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n201), .B1(new_n203), .B2(new_n189), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(KEYINPUT91), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(KEYINPUT91), .B2(new_n245), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n244), .B(KEYINPUT93), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT96), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n238), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n238), .B2(new_n250), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n188), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT97), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT97), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n188), .C1(new_n252), .C2(new_n253), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n217), .A2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n224), .A2(new_n219), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT16), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n227), .B1(new_n260), .B2(new_n210), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n245), .A2(KEYINPUT17), .A3(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n205), .A2(KEYINPUT17), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(new_n188), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n257), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n270));
  NOR2_X1   g084(.A1(G475), .A2(G902), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n271), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n254), .B2(KEYINPUT97), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n257), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n272), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n281), .A2(G122), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT14), .A3(G107), .ZN(new_n283));
  AND2_X1   g097(.A1(KEYINPUT67), .A2(G116), .ZN(new_n284));
  NOR2_X1   g098(.A1(KEYINPUT67), .A2(G116), .ZN(new_n285));
  OAI21_X1  g099(.A(G122), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G107), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n286), .A2(new_n287), .A3(new_n282), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n286), .B2(new_n282), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n283), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n286), .A2(KEYINPUT14), .A3(G107), .A4(new_n282), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n196), .A2(G128), .ZN(new_n292));
  INV_X1    g106(.A(G128), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G143), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n294), .A3(G134), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n291), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n290), .A2(KEYINPUT98), .A3(new_n291), .A4(new_n299), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n288), .A2(new_n289), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT13), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n294), .A2(new_n305), .A3(G134), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n298), .A3(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n292), .A2(new_n294), .A3(new_n305), .A4(G134), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AND4_X1   g125(.A1(new_n280), .A2(new_n302), .A3(new_n303), .A4(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n300), .B2(new_n301), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n280), .B1(new_n313), .B2(new_n303), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT9), .B(G234), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n312), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n302), .A2(new_n303), .A3(new_n311), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT99), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n280), .A3(new_n303), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT100), .B(new_n279), .C1(new_n320), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G478), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT15), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n319), .B1(new_n312), .B2(new_n314), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n318), .A3(new_n323), .ZN(new_n330));
  AOI21_X1  g144(.A(G902), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n327), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(KEYINPUT100), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G952), .ZN(new_n334));
  AOI211_X1 g148(.A(G953), .B(new_n334), .C1(G234), .C2(G237), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT21), .B(G898), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n279), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n328), .A2(new_n333), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G475), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n266), .B(new_n188), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n279), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n278), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G221), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n315), .B2(new_n279), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT81), .A3(G107), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n287), .B2(G104), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n350), .A2(G107), .ZN(new_n354));
  OAI211_X1 g168(.A(G101), .B(new_n351), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n287), .A2(G104), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n350), .A2(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n352), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n360), .A2(KEYINPUT82), .A3(G101), .A4(new_n351), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n287), .A2(G104), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n350), .B2(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n287), .A2(KEYINPUT3), .A3(G104), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT80), .B(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n357), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT69), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n227), .A2(G143), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n196), .A2(G146), .ZN(new_n373));
  AND4_X1   g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(G128), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n375), .A2(G128), .B1(new_n372), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n371), .B1(G143), .B2(new_n227), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n196), .A2(G146), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n227), .A2(G143), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n378), .A2(new_n293), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G143), .B(G146), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G128), .A3(new_n375), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n369), .A2(new_n385), .A3(KEYINPUT10), .ZN(new_n386));
  INV_X1    g200(.A(G137), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT11), .B1(new_n296), .B2(G137), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT11), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n387), .A3(G134), .ZN(new_n391));
  AOI211_X1 g205(.A(G131), .B(new_n388), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n391), .ZN(new_n393));
  INV_X1    g207(.A(new_n388), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n202), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n287), .A2(KEYINPUT3), .A3(G104), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT3), .B1(new_n287), .B2(G104), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n359), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(G101), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  INV_X1    g217(.A(G101), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n366), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n366), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(KEYINPUT0), .A2(G128), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n372), .A2(new_n373), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT0), .B(G128), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n382), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n381), .A2(new_n383), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(new_n357), .A3(new_n361), .A4(new_n368), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT10), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n386), .A2(new_n396), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n416), .A2(new_n415), .B1(new_n407), .B2(new_n412), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n419), .B(new_n396), .C1(new_n420), .C2(new_n386), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n374), .A2(new_n376), .A3(new_n370), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT69), .B1(new_n381), .B2(new_n383), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT10), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n357), .A2(new_n361), .A3(new_n368), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n417), .B(new_n413), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n396), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT83), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n418), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n191), .A2(G227), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n414), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n415), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT12), .B1(new_n436), .B2(new_n427), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n438));
  AOI211_X1 g252(.A(new_n438), .B(new_n396), .C1(new_n435), .C2(new_n415), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n418), .A2(new_n432), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n429), .A2(new_n433), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(G469), .A3(G902), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n421), .B2(new_n428), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n418), .B1(new_n437), .B2(new_n439), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n433), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(G469), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G469), .A2(G902), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n349), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G119), .B1(new_n284), .B2(new_n285), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n281), .A2(G119), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT65), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT2), .ZN(new_n456));
  INV_X1    g270(.A(G113), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT2), .A2(G113), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n454), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT67), .B(G116), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n452), .B1(new_n467), .B2(G119), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n458), .A2(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n407), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n355), .A2(new_n356), .B1(new_n366), .B2(new_n367), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n451), .A2(KEYINPUT5), .A3(new_n453), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT5), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n452), .A2(KEYINPUT84), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G119), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n477), .A3(G116), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n457), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n473), .A2(new_n481), .A3(new_n470), .A4(new_n361), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G122), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n472), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT86), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n472), .A2(new_n486), .A3(new_n482), .A4(new_n483), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n485), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n480), .A2(new_n476), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n493), .A2(new_n474), .B1(new_n468), .B2(new_n469), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n494), .A2(new_n369), .B1(new_n407), .B2(new_n471), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n492), .B1(new_n495), .B2(new_n483), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n472), .A2(new_n482), .ZN(new_n497));
  INV_X1    g311(.A(new_n483), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n491), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n374), .A2(new_n376), .A3(G125), .ZN(new_n501));
  INV_X1    g315(.A(G224), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n408), .ZN(new_n504));
  OR2_X1    g318(.A1(KEYINPUT0), .A2(G128), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n505), .C1(new_n379), .C2(new_n380), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n207), .B1(new_n506), .B2(new_n409), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n501), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n503), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n411), .A2(G125), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n381), .A2(new_n383), .A3(new_n207), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n488), .A2(new_n500), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G210), .B1(G237), .B2(G902), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n485), .A2(new_n487), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n516));
  OAI22_X1  g330(.A1(new_n501), .A2(new_n507), .B1(new_n516), .B2(new_n503), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT7), .A4(new_n509), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n474), .A2(KEYINPUT87), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT87), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n451), .A2(new_n521), .A3(KEYINPUT5), .A4(new_n453), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n493), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n470), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n369), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n483), .B(KEYINPUT8), .Z(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n494), .B2(new_n425), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n515), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n513), .A2(new_n514), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n514), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n508), .A2(new_n512), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n483), .B(new_n492), .C1(new_n472), .C2(new_n482), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n485), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n486), .B1(new_n495), .B2(new_n483), .ZN(new_n538));
  INV_X1    g352(.A(new_n487), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n528), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n279), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n531), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT88), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT88), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n450), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n477), .A2(G128), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n551), .A2(new_n552), .B1(G119), .B2(new_n293), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT24), .B(G110), .Z(new_n554));
  NOR3_X1   g368(.A1(new_n477), .A2(KEYINPUT23), .A3(G128), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT23), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(G119), .B2(new_n293), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n553), .A2(new_n554), .B1(new_n558), .B2(G110), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n258), .B2(new_n261), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n217), .A2(G146), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n553), .A2(new_n554), .B1(G110), .B2(new_n558), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(new_n562), .C1(new_n240), .C2(new_n242), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT22), .B(G137), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n279), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT77), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n569), .A2(new_n279), .A3(new_n570), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n317), .B1(G234), .B2(new_n279), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n569), .A2(new_n570), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n581), .A2(KEYINPUT78), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(KEYINPUT78), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT64), .B1(new_n387), .B2(G134), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT64), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n296), .A3(G137), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n387), .A2(G134), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G131), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n390), .B1(G134), .B2(new_n387), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n296), .A2(KEYINPUT11), .A3(G137), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n202), .B(new_n394), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n385), .A2(KEYINPUT70), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT70), .B1(new_n385), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n412), .B1(new_n392), .B2(new_n395), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT68), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n412), .B(KEYINPUT68), .C1(new_n392), .C2(new_n395), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n588), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n414), .A2(new_n597), .A3(new_n594), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT30), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n471), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT31), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n598), .B1(new_n422), .B2(new_n423), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT70), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n471), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n385), .A2(KEYINPUT70), .A3(new_n598), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n606), .A2(new_n615), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n198), .A2(G210), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n404), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n620), .B(new_n621), .Z(new_n622));
  NAND4_X1  g436(.A1(new_n611), .A2(new_n612), .A3(new_n618), .A4(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n606), .A2(new_n615), .A3(new_n617), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n610), .B1(new_n624), .B2(KEYINPUT30), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n618), .B(new_n622), .C1(new_n625), .C2(new_n616), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT31), .ZN(new_n627));
  INV_X1    g441(.A(new_n622), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT28), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT71), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n609), .A2(new_n630), .A3(new_n471), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n609), .B2(new_n471), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n629), .B1(new_n634), .B2(new_n618), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n471), .B1(new_n427), .B2(new_n412), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT28), .B1(new_n636), .B2(new_n613), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n628), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n623), .A2(new_n627), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(G472), .A2(G902), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT32), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n618), .B1(new_n625), .B2(new_n616), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n628), .ZN(new_n645));
  INV_X1    g459(.A(new_n618), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n609), .A2(new_n471), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT71), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n631), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT28), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n637), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n622), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT29), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n645), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n624), .A2(new_n471), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT72), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n618), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n624), .A2(KEYINPUT72), .A3(new_n471), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(KEYINPUT28), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(KEYINPUT29), .A3(new_n651), .A4(new_n622), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n654), .A2(new_n279), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n639), .A2(KEYINPUT32), .A3(new_n640), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n643), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n346), .A2(new_n549), .A3(new_n587), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(new_n367), .Z(G3));
  INV_X1    g480(.A(G472), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n639), .A2(new_n279), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n639), .B2(new_n279), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n429), .A2(new_n433), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n440), .A2(new_n441), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G469), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n449), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n676), .A2(new_n586), .A3(new_n348), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  AOI211_X1 g492(.A(KEYINPUT20), .B(new_n275), .C1(new_n276), .C2(new_n257), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n274), .B1(new_n269), .B2(new_n271), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n345), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n331), .A2(G478), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n329), .A2(KEYINPUT33), .A3(new_n330), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT33), .B1(new_n329), .B2(new_n330), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n326), .A2(G902), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n687), .B1(new_n278), .B2(new_n345), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n545), .A2(new_n339), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n678), .A2(new_n691), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT34), .B(G104), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G6));
  NOR2_X1   g511(.A1(new_n325), .A2(new_n327), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n332), .B1(new_n331), .B2(KEYINPUT100), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n345), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n269), .A2(new_n271), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n273), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n273), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n678), .A2(new_n694), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT35), .B(G107), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G9));
  NOR2_X1   g522(.A1(new_n568), .A2(KEYINPUT36), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n564), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n583), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n580), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n669), .A2(new_n713), .A3(new_n670), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n346), .A2(new_n714), .A3(new_n549), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT37), .B(G110), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G12));
  AOI21_X1  g531(.A(new_n344), .B1(new_n328), .B2(new_n333), .ZN(new_n718));
  INV_X1    g532(.A(G900), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n338), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n335), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n718), .B(new_n722), .C1(new_n702), .C2(new_n680), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n450), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n713), .A2(new_n545), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n724), .A2(new_n664), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT103), .B(G128), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G30));
  AOI22_X1  g543(.A1(new_n278), .A2(new_n345), .B1(new_n333), .B2(new_n328), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT40), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n722), .B(KEYINPUT39), .Z(new_n733));
  NOR2_X1   g547(.A1(new_n450), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n644), .A2(new_n622), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n279), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n622), .B1(new_n657), .B2(new_n658), .ZN(new_n738));
  OAI21_X1  g552(.A(G472), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n643), .A2(new_n663), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n543), .B(new_n741), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n544), .A2(new_n740), .A3(new_n713), .A4(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n735), .B(new_n743), .C1(new_n732), .C2(new_n734), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G143), .ZN(G45));
  AND3_X1   g559(.A1(new_n639), .A2(KEYINPUT32), .A3(new_n640), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT32), .B1(new_n639), .B2(new_n640), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n450), .B1(new_n748), .B2(new_n662), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n681), .A2(new_n688), .A3(new_n722), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n726), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  NAND3_X1  g566(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n753));
  OAI21_X1  g567(.A(G469), .B1(new_n442), .B2(G902), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n426), .A2(new_n427), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n419), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n426), .A2(KEYINPUT83), .A3(new_n427), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n432), .B1(new_n758), .B2(new_n418), .ZN(new_n759));
  INV_X1    g573(.A(new_n673), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n675), .B(new_n279), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n664), .A2(new_n587), .A3(new_n349), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT41), .B(G113), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G15));
  NAND3_X1  g580(.A1(new_n754), .A2(new_n761), .A3(new_n349), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n545), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n586), .A2(new_n339), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n705), .A2(new_n664), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G116), .ZN(G18));
  NAND4_X1  g585(.A1(new_n346), .A2(new_n664), .A3(new_n712), .A4(new_n768), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G119), .ZN(G21));
  AND2_X1   g587(.A1(new_n623), .A2(new_n627), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n659), .A2(new_n651), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n628), .ZN(new_n776));
  AOI211_X1 g590(.A(G472), .B(G902), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n667), .B1(new_n639), .B2(new_n279), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n730), .A3(new_n768), .A4(new_n769), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  NOR3_X1   g595(.A1(new_n777), .A2(new_n713), .A3(new_n778), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n750), .A2(new_n782), .A3(new_n768), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G125), .ZN(G27));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n643), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n747), .A2(KEYINPUT107), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n663), .A3(new_n662), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n676), .B2(new_n348), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n447), .A2(new_n448), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n761), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT105), .A3(new_n349), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n791), .A2(KEYINPUT42), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n795), .A3(new_n587), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n530), .A2(new_n542), .A3(new_n544), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n530), .A2(new_n542), .A3(KEYINPUT106), .A4(new_n544), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n750), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n785), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n662), .A2(new_n663), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT107), .B1(new_n641), .B2(new_n642), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n586), .B1(new_n807), .B2(new_n788), .ZN(new_n808));
  INV_X1    g622(.A(new_n722), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n689), .A2(new_n809), .A3(new_n801), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n808), .A2(KEYINPUT108), .A3(new_n810), .A4(new_n795), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n586), .B1(new_n748), .B2(new_n662), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT105), .B1(new_n793), .B2(new_n349), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n790), .B(new_n348), .C1(new_n761), .C2(new_n792), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n814), .A3(new_n801), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n815), .A3(new_n750), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT42), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n804), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT109), .B(G131), .Z(new_n820));
  XNOR2_X1  g634(.A(new_n819), .B(new_n820), .ZN(G33));
  NAND3_X1  g635(.A1(new_n812), .A2(new_n815), .A3(new_n724), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G134), .ZN(G36));
  AOI21_X1  g637(.A(new_n344), .B1(new_n704), .B2(new_n272), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n688), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT43), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n671), .A2(new_n713), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT44), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(KEYINPUT44), .A3(new_n828), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n444), .A2(new_n446), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT45), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT45), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(G469), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n448), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT46), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n443), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n837), .A2(KEYINPUT110), .A3(KEYINPUT46), .A4(new_n448), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n349), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n733), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n831), .A2(new_n802), .A3(new_n832), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G137), .ZN(G39));
  XOR2_X1   g661(.A(new_n844), .B(KEYINPUT47), .Z(new_n848));
  NOR3_X1   g662(.A1(new_n803), .A2(new_n587), .A3(new_n664), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n211), .ZN(G42));
  XOR2_X1   g665(.A(new_n762), .B(KEYINPUT49), .Z(new_n852));
  INV_X1    g666(.A(new_n742), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n587), .A3(new_n544), .A4(new_n349), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n852), .A2(new_n854), .A3(new_n740), .A4(new_n825), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT111), .Z(new_n856));
  NOR2_X1   g670(.A1(new_n801), .A2(new_n767), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n827), .A2(new_n335), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT48), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n858), .B(new_n808), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n586), .A2(new_n721), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n827), .A2(new_n779), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n768), .ZN(new_n865));
  INV_X1    g679(.A(new_n740), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n863), .A3(new_n857), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n691), .A3(new_n693), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(G952), .A3(new_n191), .A4(new_n868), .ZN(new_n869));
  AOI211_X1 g683(.A(KEYINPUT115), .B(KEYINPUT48), .C1(new_n858), .C2(new_n808), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n862), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n762), .A2(new_n348), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n848), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n864), .A2(new_n802), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n742), .A2(new_n544), .A3(new_n767), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n864), .A2(KEYINPUT50), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n881), .A3(KEYINPUT114), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n681), .A2(new_n688), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n858), .A2(new_n782), .B1(new_n867), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT51), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n882), .B2(KEYINPUT51), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n871), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n749), .B(new_n726), .C1(new_n750), .C2(new_n724), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n450), .A2(new_n712), .A3(new_n809), .ZN(new_n891));
  INV_X1    g705(.A(new_n545), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n730), .A3(new_n892), .A4(new_n740), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n783), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n890), .A2(KEYINPUT52), .A3(new_n783), .A4(new_n893), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n815), .A2(new_n750), .A3(new_n782), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n344), .A2(new_n809), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n712), .A2(new_n333), .A3(new_n900), .A4(new_n328), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n704), .B2(new_n703), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n664), .A3(new_n725), .A4(new_n802), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n822), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT112), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n278), .A2(new_n905), .A3(new_n718), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n679), .A2(new_n680), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT112), .B1(new_n907), .B2(new_n700), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n692), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n339), .B1(new_n546), .B2(new_n548), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n671), .A3(new_n677), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n665), .B(new_n715), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n780), .A2(new_n772), .A3(new_n770), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n764), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n819), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n889), .B1(new_n898), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n664), .A2(new_n768), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n824), .A2(new_n341), .A3(new_n712), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n769), .B(new_n718), .C1(new_n702), .C2(new_n680), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(new_n780), .C1(new_n753), .C2(new_n763), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n923), .A2(new_n912), .A3(new_n904), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n896), .A2(new_n897), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT53), .A4(new_n819), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT54), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT113), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n917), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  OAI211_X1 g744(.A(KEYINPUT113), .B(new_n889), .C1(new_n898), .C2(new_n916), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n932), .B2(KEYINPUT54), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n888), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(G952), .A2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n856), .B1(new_n934), .B2(new_n935), .ZN(G75));
  NAND3_X1  g750(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n488), .A2(new_n500), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT116), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n532), .B(KEYINPUT117), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n937), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n937), .B2(new_n938), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n191), .A2(G952), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G51));
  XOR2_X1   g761(.A(new_n448), .B(KEYINPUT57), .Z(new_n948));
  AND2_X1   g762(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n759), .B2(new_n760), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n837), .B(KEYINPUT118), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n932), .A2(G902), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n946), .B1(new_n952), .B2(new_n954), .ZN(G54));
  NAND4_X1  g769(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n956));
  INV_X1    g770(.A(new_n269), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n946), .ZN(G60));
  XNOR2_X1  g774(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n326), .A2(new_n279), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n685), .B(KEYINPUT119), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n963), .B(new_n964), .C1(new_n949), .C2(new_n950), .ZN(new_n965));
  INV_X1    g779(.A(new_n946), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n964), .B1(new_n933), .B2(new_n963), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  NAND3_X1  g785(.A1(new_n930), .A2(new_n931), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n582), .A2(new_n584), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n930), .A2(KEYINPUT121), .A3(new_n931), .A4(new_n971), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n966), .ZN(new_n978));
  INV_X1    g792(.A(new_n710), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n974), .B2(new_n976), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT122), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n978), .B(new_n981), .C1(new_n982), .C2(KEYINPUT61), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n977), .A2(new_n982), .A3(new_n966), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n977), .A2(new_n966), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n984), .B(new_n985), .C1(new_n986), .C2(new_n980), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n987), .ZN(G66));
  OAI21_X1  g802(.A(G953), .B1(new_n337), .B2(new_n502), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n923), .A2(new_n912), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(G953), .ZN(new_n991));
  INV_X1    g805(.A(new_n940), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(G898), .B2(new_n191), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n991), .B(new_n993), .ZN(G69));
  INV_X1    g808(.A(new_n845), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n808), .A2(new_n892), .A3(new_n730), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n890), .A2(new_n783), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n848), .A2(new_n849), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1002), .A2(new_n822), .A3(new_n846), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1001), .A2(new_n1003), .A3(new_n819), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1001), .A2(new_n1003), .A3(KEYINPUT127), .A4(new_n819), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(new_n191), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n226), .A2(new_n235), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT123), .Z(new_n1010));
  XOR2_X1   g824(.A(new_n625), .B(new_n1010), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(G900), .B2(G953), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n909), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n812), .A3(new_n734), .A4(new_n802), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n846), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT124), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n999), .A2(new_n744), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n850), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(G953), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT125), .ZN(new_n1025));
  OR3_X1    g839(.A1(new_n1024), .A2(new_n1025), .A3(new_n1011), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1024), .B2(new_n1011), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1014), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1029), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1014), .A2(new_n1026), .A3(new_n1031), .A4(new_n1027), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(G72));
  NAND3_X1  g847(.A1(new_n1006), .A2(new_n990), .A3(new_n1007), .ZN(new_n1034));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  AOI211_X1 g850(.A(new_n622), .B(new_n644), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1019), .A2(new_n990), .A3(new_n1023), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n736), .B1(new_n1038), .B2(new_n1036), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n645), .A2(new_n626), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n927), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n966), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(G57));
endmodule


