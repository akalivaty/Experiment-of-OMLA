//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT72), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(G197gat), .ZN(new_n210));
  INV_X1    g009(.A(G204gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI211_X1 g015(.A(KEYINPUT70), .B(new_n209), .C1(new_n212), .C2(new_n213), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n208), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n207), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G226gat), .ZN(new_n222));
  INV_X1    g021(.A(G233gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT27), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT28), .ZN(new_n229));
  NOR4_X1   g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .A4(G190gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT66), .B1(new_n225), .B2(KEYINPUT27), .ZN(new_n231));
  AOI21_X1  g030(.A(G190gat), .B1(new_n225), .B2(KEYINPUT27), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(new_n227), .A3(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n231), .A2(new_n232), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n236), .A2(new_n229), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n230), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT26), .ZN(new_n244));
  INV_X1    g043(.A(G169gat), .ZN(new_n245));
  INV_X1    g044(.A(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248));
  INV_X1    g047(.A(G190gat), .ZN(new_n249));
  OAI22_X1  g048(.A1(new_n247), .A2(new_n248), .B1(new_n225), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n241), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n243), .B2(KEYINPUT23), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(KEYINPUT65), .A3(new_n253), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n225), .A2(new_n249), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT64), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT25), .B1(new_n258), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n257), .A2(new_n256), .ZN(new_n270));
  INV_X1    g069(.A(new_n254), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT25), .B1(new_n261), .B2(new_n263), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI22_X1  g073(.A1(new_n240), .A2(new_n252), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n224), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n224), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n239), .A2(new_n229), .A3(new_n236), .ZN(new_n279));
  INV_X1    g078(.A(new_n230), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n251), .ZN(new_n282));
  INV_X1    g081(.A(new_n267), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n259), .B(new_n260), .C1(new_n263), .C2(new_n266), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n270), .B(new_n271), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n273), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n258), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n278), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n277), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n285), .A2(new_n286), .B1(new_n258), .B2(new_n288), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n252), .B1(new_n279), .B2(new_n280), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n276), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT71), .B1(new_n295), .B2(new_n278), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n221), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n278), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n224), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n221), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n206), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n300), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n304), .B2(KEYINPUT71), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n301), .B(new_n205), .C1(new_n305), .C2(new_n221), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT30), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n298), .A2(new_n302), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n205), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT85), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT40), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G141gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(new_n325), .B2(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n318), .A2(G141gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n314), .A2(G148gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n322), .ZN(new_n333));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n328), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT2), .B1(new_n315), .B2(new_n319), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n325), .A2(new_n322), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(KEYINPUT73), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n327), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT75), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT73), .B1(new_n337), .B2(new_n338), .ZN(new_n342));
  XNOR2_X1  g141(.A(G141gat), .B(G148gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n335), .B(new_n328), .C1(new_n343), .C2(KEYINPUT2), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n327), .ZN(new_n347));
  XOR2_X1   g146(.A(G127gat), .B(G134gat), .Z(new_n348));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(KEYINPUT1), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G113gat), .B(G120gat), .Z(new_n351));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n341), .A2(KEYINPUT77), .A3(new_n347), .A4(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n345), .A2(new_n346), .A3(new_n327), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n346), .B1(new_n345), .B2(new_n327), .ZN(new_n358));
  INV_X1    g157(.A(new_n355), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n342), .A2(new_n344), .B1(new_n326), .B2(new_n321), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n359), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT39), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n341), .A2(new_n369), .A3(KEYINPUT3), .A4(new_n347), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n357), .A2(new_n358), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT76), .B1(new_n361), .B2(new_n371), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n355), .B(new_n370), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n350), .A2(new_n354), .A3(KEYINPUT68), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT68), .B1(new_n350), .B2(new_n354), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(KEYINPUT78), .A3(new_n378), .A4(new_n361), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n362), .B2(KEYINPUT4), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT68), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n350), .A2(new_n354), .A3(KEYINPUT68), .ZN(new_n384));
  AND4_X1   g183(.A1(new_n378), .A2(new_n383), .A3(new_n361), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n379), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n366), .B1(new_n374), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n368), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT0), .ZN(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT39), .ZN(new_n395));
  AOI211_X1 g194(.A(KEYINPUT84), .B(new_n394), .C1(new_n387), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n357), .A2(new_n358), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n373), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n370), .A2(new_n355), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n386), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n366), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n403), .B2(new_n393), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n389), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n311), .B1(new_n313), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n362), .A2(new_n378), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n383), .A2(new_n361), .A3(KEYINPUT4), .A4(new_n384), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n366), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n399), .B2(new_n400), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n402), .B(new_n356), .C1(new_n360), .C2(new_n364), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT5), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n374), .A2(new_n386), .A3(new_n414), .ZN(new_n415));
  AOI211_X1 g214(.A(KEYINPUT86), .B(new_n393), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n370), .A2(new_n355), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n369), .B1(new_n340), .B2(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n341), .A2(new_n347), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(new_n371), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n409), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n412), .A2(KEYINPUT5), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n415), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n417), .B1(new_n424), .B2(new_n394), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n313), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n389), .C1(new_n396), .C2(new_n404), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT87), .B1(new_n406), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(KEYINPUT39), .B(new_n366), .C1(new_n374), .C2(new_n386), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT84), .B1(new_n431), .B2(new_n394), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n403), .A2(new_n397), .A3(new_n393), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n388), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n310), .B(new_n307), .C1(new_n434), .C2(new_n427), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(new_n428), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT31), .B(G50gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G228gat), .A2(G233gat), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n218), .B2(new_n220), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n341), .B(new_n347), .C1(new_n445), .C2(KEYINPUT3), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n276), .B1(new_n340), .B2(KEYINPUT3), .ZN(new_n447));
  INV_X1    g246(.A(new_n221), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n361), .B2(new_n371), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n444), .B1(new_n451), .B2(new_n221), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n212), .A2(new_n213), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT70), .B1(new_n453), .B2(new_n209), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n207), .B1(new_n454), .B2(new_n219), .ZN(new_n455));
  INV_X1    g254(.A(new_n220), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n276), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n361), .B1(new_n457), .B2(new_n371), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(G22gat), .B1(new_n450), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n340), .B1(new_n445), .B2(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n449), .A3(new_n444), .ZN(new_n462));
  INV_X1    g261(.A(G22gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n371), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n464), .A2(new_n398), .B1(new_n448), .B2(new_n447), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n462), .B(new_n463), .C1(new_n465), .C2(new_n444), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n443), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n460), .A2(KEYINPUT81), .A3(new_n466), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n469), .B2(new_n468), .ZN(new_n473));
  INV_X1    g272(.A(new_n443), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n440), .B(new_n471), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n466), .A3(KEYINPUT81), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT82), .B1(new_n478), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n424), .A2(new_n394), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT86), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n393), .B1(new_n413), .B2(new_n415), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n417), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n415), .B(new_n393), .C1(new_n422), .C2(new_n423), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n426), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n394), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n301), .B1(new_n305), .B2(new_n221), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n206), .B1(new_n494), .B2(KEYINPUT37), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n305), .A2(new_n221), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n304), .A2(KEYINPUT89), .A3(new_n448), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n221), .B1(new_n299), .B2(new_n300), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT38), .B1(new_n501), .B2(KEYINPUT37), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n494), .A2(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT38), .B1(new_n504), .B2(new_n495), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n505), .A3(new_n306), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n480), .B1(new_n493), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT90), .B1(new_n439), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n406), .A2(new_n429), .A3(KEYINPUT87), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n437), .B1(new_n435), .B2(new_n436), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n503), .A2(new_n505), .A3(new_n306), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(new_n492), .A3(new_n491), .A4(new_n489), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .A4(new_n480), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n485), .A2(new_n486), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n492), .B1(new_n517), .B2(new_n483), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n311), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n311), .A2(new_n518), .A3(KEYINPUT79), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT83), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT83), .B1(new_n475), .B2(new_n479), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G43gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n275), .A2(new_n377), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n282), .B(new_n290), .C1(new_n375), .C2(new_n376), .ZN(new_n531));
  INV_X1    g330(.A(G227gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(new_n223), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n529), .B1(new_n534), .B2(KEYINPUT32), .ZN(new_n535));
  INV_X1    g334(.A(new_n534), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(KEYINPUT33), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n530), .B2(new_n531), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT34), .ZN(new_n539));
  INV_X1    g338(.A(new_n529), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT69), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(KEYINPUT69), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT33), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n534), .A2(KEYINPUT32), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n539), .B1(new_n544), .B2(new_n537), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT36), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n526), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n516), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n480), .A2(new_n521), .A3(new_n522), .A4(new_n548), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT35), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n554), .B2(KEYINPUT35), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n546), .B2(new_n547), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n544), .ZN(new_n560));
  INV_X1    g359(.A(new_n539), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(KEYINPUT91), .A3(new_n545), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT35), .B1(new_n307), .B2(new_n310), .ZN(new_n565));
  AND4_X1   g364(.A1(new_n480), .A2(new_n493), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n556), .A2(new_n557), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(G1gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT16), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(G8gat), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n573), .B(new_n575), .C1(new_n572), .C2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(G8gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n580));
  AOI21_X1  g379(.A(G36gat), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G29gat), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n582), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G43gat), .B(G50gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(KEYINPUT93), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n581), .A2(new_n583), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT94), .B(G50gat), .Z(new_n594));
  OAI211_X1 g393(.A(new_n584), .B(new_n593), .C1(G43gat), .C2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n597), .A3(new_n595), .ZN(new_n598));
  INV_X1    g397(.A(new_n577), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n576), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n592), .B2(new_n595), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n570), .B(new_n596), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT18), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n602), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n600), .A3(new_n598), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n607), .A2(KEYINPUT18), .A3(new_n570), .A4(new_n596), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n595), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n600), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n596), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n570), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n605), .A2(new_n608), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G197gat), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT11), .B(G169gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n603), .A2(new_n604), .B1(new_n611), .B2(new_n614), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n621), .A3(new_n608), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(G57gat), .A2(G64gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G57gat), .A2(G64gat), .ZN(new_n628));
  INV_X1    g427(.A(G71gat), .ZN(new_n629));
  INV_X1    g428(.A(G78gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n627), .B(new_n628), .C1(new_n631), .C2(KEYINPUT9), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n633));
  XNOR2_X1  g432(.A(G71gat), .B(G78gat), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n578), .B1(KEYINPUT21), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT98), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n323), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n640), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT21), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G127gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n643), .A2(new_n655), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n592), .A2(new_n595), .ZN(new_n660));
  XOR2_X1   g459(.A(G99gat), .B(G106gat), .Z(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n662));
  INV_X1    g461(.A(G85gat), .ZN(new_n663));
  INV_X1    g462(.A(G92gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G99gat), .A2(G106gat), .ZN(new_n667));
  AOI22_X1  g466(.A1(KEYINPUT8), .A2(new_n667), .B1(new_n663), .B2(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n662), .A2(new_n665), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n661), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n662), .A2(new_n665), .ZN(new_n672));
  INV_X1    g471(.A(new_n661), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n666), .A4(new_n668), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(G232gat), .A2(G233gat), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n660), .A2(new_n676), .B1(KEYINPUT41), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n598), .A2(new_n675), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n602), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G190gat), .B(G218gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n678), .B(new_n683), .C1(new_n602), .C2(new_n679), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n677), .A2(KEYINPUT41), .ZN(new_n685));
  XNOR2_X1  g484(.A(G134gat), .B(G162gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AND4_X1   g486(.A1(KEYINPUT100), .A2(new_n682), .A3(new_n684), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n690), .A2(new_n687), .B1(new_n682), .B2(new_n684), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(G230gat), .A2(G233gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n637), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT10), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n671), .B(new_n674), .C1(new_n636), .C2(new_n635), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n676), .A2(new_n638), .A3(KEYINPUT10), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(new_n698), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n695), .ZN(new_n703));
  XNOR2_X1  g502(.A(G120gat), .B(G148gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(G176gat), .B(G204gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(new_n706));
  OR2_X1    g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n699), .A2(new_n700), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n694), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n695), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n659), .A2(new_n693), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n569), .A2(new_n626), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n518), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n572), .ZN(G1324gat));
  OAI21_X1  g515(.A(G8gat), .B1(new_n714), .B2(new_n311), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT102), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n714), .A2(new_n311), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT16), .B(G8gat), .Z(new_n720));
  AOI21_X1  g519(.A(KEYINPUT101), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(G1325gat));
  INV_X1    g523(.A(G15gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n564), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n714), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT103), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n714), .A2(new_n725), .A3(new_n550), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1326gat));
  OR2_X1    g529(.A1(new_n524), .A2(new_n525), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n714), .A2(KEYINPUT104), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT104), .B1(new_n714), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT43), .B(G22gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1327gat));
  INV_X1    g536(.A(new_n659), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(new_n692), .A3(new_n712), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n569), .A2(new_n626), .A3(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(G29gat), .A3(new_n518), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT45), .Z(new_n742));
  AOI21_X1  g541(.A(new_n551), .B1(new_n508), .B2(new_n515), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n693), .B1(new_n743), .B2(new_n567), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT44), .B(new_n693), .C1(new_n743), .C2(new_n567), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n626), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n738), .A2(new_n749), .A3(new_n712), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G29gat), .B1(new_n751), .B2(new_n518), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n742), .A2(new_n752), .ZN(G1328gat));
  NOR3_X1   g552(.A1(new_n740), .A2(G36gat), .A3(new_n311), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT46), .ZN(new_n755));
  OAI21_X1  g554(.A(G36gat), .B1(new_n751), .B2(new_n311), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1329gat));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n740), .B2(new_n726), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n549), .A2(G43gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n751), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(new_n759), .C1(new_n751), .C2(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1330gat));
  OAI21_X1  g564(.A(new_n594), .B1(new_n751), .B2(new_n480), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n740), .A2(new_n594), .A3(new_n732), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n748), .A2(new_n731), .A3(new_n750), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n767), .B1(new_n771), .B2(new_n594), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(KEYINPUT48), .B2(new_n772), .ZN(G1331gat));
  NAND4_X1  g572(.A1(new_n738), .A2(new_n749), .A3(new_n692), .A4(new_n712), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n553), .B2(new_n568), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n518), .B(KEYINPUT105), .Z(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g578(.A(new_n311), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT106), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n782), .B(new_n783), .Z(G1333gat));
  AOI21_X1  g583(.A(new_n629), .B1(new_n775), .B2(new_n549), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n726), .A2(G71gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n775), .A2(new_n731), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  INV_X1    g589(.A(new_n712), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n738), .A2(new_n626), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n748), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n518), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n738), .A2(new_n626), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n569), .A2(KEYINPUT51), .A3(new_n693), .A4(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  INV_X1    g596(.A(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n744), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n518), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n663), .A3(new_n712), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n794), .B1(new_n800), .B2(new_n802), .ZN(G1336gat));
  NOR3_X1   g602(.A1(new_n311), .A2(G92gat), .A3(new_n791), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT108), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n311), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n746), .A2(new_n807), .A3(new_n747), .A4(new_n792), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(new_n808), .B2(G92gat), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n796), .B2(new_n799), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT107), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n808), .A2(new_n814), .A3(G92gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n808), .B2(G92gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n810), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(G1337gat));
  OAI21_X1  g618(.A(G99gat), .B1(new_n793), .B2(new_n550), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n726), .A2(G99gat), .A3(new_n791), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n800), .B2(new_n821), .ZN(G1338gat));
  NAND2_X1  g621(.A1(new_n796), .A2(new_n799), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n480), .A2(G106gat), .A3(new_n791), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n746), .A2(new_n731), .A3(new_n747), .A4(new_n792), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n830));
  INV_X1    g629(.A(new_n480), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n746), .A2(new_n831), .A3(new_n747), .A4(new_n792), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G106gat), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n829), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(G1339gat));
  NAND3_X1  g635(.A1(new_n699), .A2(new_n700), .A3(new_n695), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n709), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n706), .B1(new_n701), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n711), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT110), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n844), .A3(new_n711), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n838), .A2(new_n840), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n843), .A2(new_n626), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n570), .B1(new_n607), .B2(new_n596), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n611), .A2(new_n614), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n620), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n625), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n712), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n692), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n843), .A2(new_n845), .A3(new_n848), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n853), .B1(new_n688), .B2(new_n691), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT111), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n693), .B1(new_n849), .B2(new_n854), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n659), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n713), .A2(new_n749), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(KEYINPUT112), .A3(new_n866), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n480), .A3(new_n548), .A4(new_n777), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n807), .ZN(new_n873));
  INV_X1    g672(.A(G113gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n874), .A3(new_n626), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n807), .A2(new_n518), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n731), .A2(new_n726), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n749), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n878), .A2(new_n883), .A3(new_n791), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n873), .A2(new_n712), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n883), .ZN(G1341gat));
  NOR3_X1   g685(.A1(new_n878), .A2(new_n649), .A3(new_n659), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n807), .A3(new_n659), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(G127gat), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(G1342gat));
  OR2_X1    g691(.A1(new_n878), .A2(new_n692), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n693), .A2(new_n311), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT115), .Z(new_n895));
  INV_X1    g694(.A(G134gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n872), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n893), .A2(G134gat), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT116), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(KEYINPUT116), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(G1343gat));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n842), .B1(new_n847), .B2(new_n846), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n909), .A2(new_n626), .B1(new_n712), .B2(new_n853), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n859), .B1(new_n693), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n911), .A2(new_n659), .B1(new_n749), .B2(new_n713), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n659), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n866), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n731), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n869), .A2(new_n831), .A3(new_n870), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n550), .A2(new_n876), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n749), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n906), .B1(new_n922), .B2(new_n314), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n919), .ZN(new_n924));
  INV_X1    g723(.A(new_n917), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n921), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n626), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n869), .A2(new_n870), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n549), .A2(new_n480), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n930), .A2(new_n807), .A3(new_n776), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n314), .A3(new_n626), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT58), .ZN(new_n936));
  NOR2_X1   g735(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n937));
  AND2_X1   g736(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n938));
  OAI221_X1 g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .C1(new_n922), .C2(new_n314), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1344gat));
  NAND2_X1  g739(.A1(new_n918), .A2(KEYINPUT57), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n912), .A2(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n912), .A2(KEYINPUT121), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n942), .A2(new_n919), .A3(new_n731), .A4(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n941), .A2(new_n712), .A3(new_n927), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G148gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n712), .A3(new_n927), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n318), .A2(KEYINPUT59), .ZN(new_n948));
  AOI22_X1  g747(.A1(KEYINPUT59), .A2(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n791), .A2(G148gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n933), .A2(KEYINPUT120), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT120), .B1(new_n933), .B2(new_n950), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT122), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n953), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n951), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n947), .A2(new_n948), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n960), .B1(new_n945), .B2(G148gat), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n955), .A2(new_n962), .ZN(G1345gat));
  NAND3_X1  g762(.A1(new_n933), .A2(new_n323), .A3(new_n738), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n920), .A2(new_n659), .A3(new_n921), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n323), .ZN(G1346gat));
  NOR3_X1   g765(.A1(new_n930), .A2(new_n776), .A3(new_n932), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(new_n324), .A3(new_n895), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n920), .A2(new_n692), .A3(new_n921), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n324), .ZN(G1347gat));
  NOR2_X1   g769(.A1(new_n777), .A2(new_n311), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n871), .A2(new_n877), .A3(new_n971), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n972), .A2(new_n245), .A3(new_n749), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n930), .A2(new_n801), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n480), .A2(new_n807), .A3(new_n548), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n626), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n973), .B1(new_n977), .B2(new_n245), .ZN(G1348gat));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n246), .A3(new_n712), .ZN(new_n979));
  OAI21_X1  g778(.A(G176gat), .B1(new_n972), .B2(new_n791), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1349gat));
  OAI21_X1  g780(.A(G183gat), .B1(new_n972), .B2(new_n659), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n659), .A2(new_n226), .A3(new_n228), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n974), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT124), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n982), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n986), .A2(new_n990), .A3(KEYINPUT60), .A4(new_n988), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1350gat));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n249), .A3(new_n693), .ZN(new_n995));
  OAI21_X1  g794(.A(G190gat), .B1(new_n972), .B2(new_n692), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n999), .B(G190gat), .C1(new_n972), .C2(new_n692), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n998), .B1(new_n997), .B2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(G1351gat));
  NAND3_X1  g802(.A1(new_n974), .A2(new_n807), .A3(new_n931), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n1005));
  OR2_X1    g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1006), .A2(new_n626), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n941), .A2(new_n944), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n971), .A2(new_n550), .ZN(new_n1010));
  XOR2_X1   g809(.A(new_n1010), .B(KEYINPUT127), .Z(new_n1011));
  NOR2_X1   g810(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n749), .A2(new_n210), .ZN(new_n1013));
  AOI22_X1  g812(.A1(new_n1008), .A2(new_n210), .B1(new_n1012), .B2(new_n1013), .ZN(G1352gat));
  NAND2_X1  g813(.A1(new_n712), .A2(new_n211), .ZN(new_n1015));
  OR3_X1    g814(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n941), .A2(new_n712), .A3(new_n944), .ZN(new_n1017));
  OAI21_X1  g816(.A(G204gat), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1018));
  OAI21_X1  g817(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1015), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(G1353gat));
  NOR2_X1   g819(.A1(new_n659), .A2(G211gat), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n1007), .A3(new_n1021), .ZN(new_n1022));
  OR3_X1    g821(.A1(new_n1009), .A2(new_n659), .A3(new_n1010), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1023), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1023), .B2(G211gat), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G1354gat));
  NAND3_X1  g825(.A1(new_n1006), .A2(new_n693), .A3(new_n1007), .ZN(new_n1027));
  INV_X1    g826(.A(G218gat), .ZN(new_n1028));
  NOR2_X1   g827(.A1(new_n692), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g828(.A1(new_n1027), .A2(new_n1028), .B1(new_n1012), .B2(new_n1029), .ZN(G1355gat));
endmodule


