

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U558 ( .A(n543), .B(n542), .ZN(n664) );
  XNOR2_X1 U559 ( .A(n536), .B(n535), .ZN(n537) );
  NOR2_X2 U560 ( .A1(n802), .A2(n801), .ZN(n803) );
  AND2_X2 U561 ( .A1(n826), .A2(n526), .ZN(n828) );
  OR2_X2 U562 ( .A1(n664), .A2(n548), .ZN(n544) );
  NOR2_X1 U563 ( .A1(n747), .A2(n746), .ZN(n754) );
  AND2_X1 U564 ( .A1(n754), .A2(n1029), .ZN(n748) );
  AND2_X1 U565 ( .A1(n815), .A2(n795), .ZN(n794) );
  INV_X1 U566 ( .A(G2105), .ZN(n533) );
  XNOR2_X1 U567 ( .A(KEYINPUT68), .B(G543), .ZN(n543) );
  OR2_X1 U568 ( .A1(n824), .A2(n823), .ZN(n525) );
  AND2_X1 U569 ( .A1(n825), .A2(n525), .ZN(n526) );
  INV_X1 U570 ( .A(KEYINPUT29), .ZN(n770) );
  XNOR2_X1 U571 ( .A(n770), .B(KEYINPUT102), .ZN(n771) );
  BUF_X1 U572 ( .A(n742), .Z(n778) );
  NOR2_X1 U573 ( .A1(G1966), .A2(n824), .ZN(n788) );
  NOR2_X1 U574 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U575 ( .A1(n742), .A2(G8), .ZN(n824) );
  INV_X1 U576 ( .A(KEYINPUT109), .ZN(n827) );
  INV_X1 U577 ( .A(KEYINPUT23), .ZN(n534) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n527) );
  XNOR2_X1 U579 ( .A(n534), .B(KEYINPUT66), .ZN(n535) );
  NOR2_X1 U580 ( .A1(n830), .A2(n829), .ZN(n832) );
  INV_X1 U581 ( .A(KEYINPUT0), .ZN(n542) );
  NOR2_X1 U582 ( .A1(n540), .A2(n539), .ZN(n694) );
  BUF_X1 U583 ( .A(n694), .Z(G160) );
  NOR2_X2 U584 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U585 ( .A(n528), .B(n527), .ZN(n897) );
  NAND2_X1 U586 ( .A1(n897), .A2(G137), .ZN(n531) );
  INV_X1 U587 ( .A(G2105), .ZN(n529) );
  NOR2_X2 U588 ( .A1(G2104), .A2(n529), .ZN(n893) );
  NAND2_X1 U589 ( .A1(G125), .A2(n893), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n531), .A2(n530), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XNOR2_X2 U592 ( .A(n532), .B(KEYINPUT67), .ZN(n892) );
  NAND2_X1 U593 ( .A1(G113), .A2(n892), .ZN(n538) );
  AND2_X4 U594 ( .A1(n533), .A2(G2104), .ZN(n896) );
  NAND2_X1 U595 ( .A1(G101), .A2(n896), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n650) );
  NAND2_X1 U598 ( .A1(n650), .A2(G89), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n541), .B(KEYINPUT4), .ZN(n546) );
  INV_X1 U600 ( .A(G651), .ZN(n548) );
  XNOR2_X2 U601 ( .A(KEYINPUT69), .B(n544), .ZN(n655) );
  NAND2_X1 U602 ( .A1(G76), .A2(n655), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U604 ( .A(KEYINPUT5), .B(n547), .ZN(n555) );
  NOR2_X1 U605 ( .A1(G543), .A2(n548), .ZN(n549) );
  XOR2_X2 U606 ( .A(KEYINPUT1), .B(n549), .Z(n662) );
  NAND2_X1 U607 ( .A1(n662), .A2(G63), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT75), .B(n550), .Z(n552) );
  NOR2_X2 U609 ( .A1(G651), .A2(n664), .ZN(n658) );
  NAND2_X1 U610 ( .A1(n658), .A2(G51), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n556), .ZN(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U616 ( .A1(G102), .A2(n896), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G138), .A2(n897), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G114), .A2(n892), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G126), .A2(n893), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G52), .A2(n658), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G64), .A2(n662), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G90), .A2(n650), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G77), .A2(n655), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U630 ( .A1(n569), .A2(n568), .ZN(G171) );
  AND2_X1 U631 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U632 ( .A(G132), .ZN(G219) );
  INV_X1 U633 ( .A(G82), .ZN(G220) );
  INV_X1 U634 ( .A(G57), .ZN(G237) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n849) );
  NAND2_X1 U638 ( .A1(n849), .A2(G567), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n571), .B(KEYINPUT71), .ZN(n572) );
  XNOR2_X1 U640 ( .A(KEYINPUT11), .B(n572), .ZN(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n662), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT14), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G43), .A2(n658), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT72), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n650), .A2(G81), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G68), .A2(n655), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X2 U651 ( .A1(n582), .A2(n581), .ZN(n1034) );
  NAND2_X1 U652 ( .A1(n1034), .A2(G860), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G54), .A2(n658), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT74), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G92), .A2(n650), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G79), .A2(n655), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G66), .A2(n662), .ZN(n586) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n586), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X2 U664 ( .A(KEYINPUT15), .B(n591), .ZN(n1029) );
  INV_X1 U665 ( .A(n1029), .ZN(n608) );
  INV_X1 U666 ( .A(G868), .ZN(n676) );
  NAND2_X1 U667 ( .A1(n608), .A2(n676), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G53), .A2(n658), .ZN(n595) );
  NAND2_X1 U670 ( .A1(G65), .A2(n662), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U672 ( .A(KEYINPUT70), .B(n596), .Z(n600) );
  NAND2_X1 U673 ( .A1(G91), .A2(n650), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G78), .A2(n655), .ZN(n597) );
  AND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(G299) );
  XNOR2_X1 U677 ( .A(KEYINPUT76), .B(n676), .ZN(n601) );
  NOR2_X1 U678 ( .A1(G286), .A2(n601), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT77), .B(n602), .Z(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(G297) );
  INV_X1 U682 ( .A(G860), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n606), .A2(n1029), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(n608), .A2(n676), .ZN(n609) );
  XOR2_X1 U687 ( .A(KEYINPUT78), .B(n609), .Z(n610) );
  NOR2_X1 U688 ( .A1(G559), .A2(n610), .ZN(n612) );
  AND2_X1 U689 ( .A1(n676), .A2(n1034), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U691 ( .A(KEYINPUT79), .B(n613), .Z(G282) );
  NAND2_X1 U692 ( .A1(G123), .A2(n893), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT18), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G99), .A2(n896), .ZN(n615) );
  XNOR2_X1 U695 ( .A(n615), .B(KEYINPUT80), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G111), .A2(n892), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G135), .A2(n897), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n948) );
  XNOR2_X1 U701 ( .A(G2096), .B(n948), .ZN(n623) );
  INV_X1 U702 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G67), .A2(n662), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G93), .A2(n650), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G80), .A2(n655), .ZN(n626) );
  XNOR2_X1 U708 ( .A(KEYINPUT81), .B(n626), .ZN(n627) );
  NOR2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n658), .A2(G55), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n675) );
  NAND2_X1 U712 ( .A1(G559), .A2(n1029), .ZN(n631) );
  XOR2_X1 U713 ( .A(n1034), .B(n631), .Z(n673) );
  NOR2_X1 U714 ( .A1(G860), .A2(n673), .ZN(n632) );
  XOR2_X1 U715 ( .A(n675), .B(n632), .Z(G145) );
  NAND2_X1 U716 ( .A1(G50), .A2(n658), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G62), .A2(n662), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G88), .A2(n650), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G75), .A2(n655), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT86), .B(n639), .Z(G303) );
  NAND2_X1 U724 ( .A1(n655), .A2(G73), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n640) );
  XNOR2_X1 U726 ( .A(KEYINPUT84), .B(n640), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n642), .B(n641), .ZN(n649) );
  NAND2_X1 U728 ( .A1(G48), .A2(n658), .ZN(n644) );
  NAND2_X1 U729 ( .A1(G61), .A2(n662), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G86), .A2(n650), .ZN(n645) );
  XNOR2_X1 U732 ( .A(KEYINPUT83), .B(n645), .ZN(n646) );
  NOR2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(G305) );
  AND2_X1 U735 ( .A1(n662), .A2(G60), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G47), .A2(n658), .ZN(n652) );
  NAND2_X1 U737 ( .A1(G85), .A2(n650), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n655), .A2(G72), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n657), .A2(n656), .ZN(G290) );
  NAND2_X1 U742 ( .A1(G49), .A2(n658), .ZN(n660) );
  NAND2_X1 U743 ( .A1(G74), .A2(G651), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n663), .B(KEYINPUT82), .ZN(n666) );
  NAND2_X1 U747 ( .A1(G87), .A2(n664), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n666), .A2(n665), .ZN(G288) );
  XNOR2_X1 U749 ( .A(G303), .B(G305), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n667), .B(n675), .ZN(n668) );
  XNOR2_X1 U751 ( .A(KEYINPUT87), .B(n668), .ZN(n670) );
  XNOR2_X1 U752 ( .A(G290), .B(KEYINPUT19), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U754 ( .A(n671), .B(G299), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(G288), .ZN(n917) );
  XNOR2_X1 U756 ( .A(n673), .B(n917), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G868), .ZN(n678) );
  NAND2_X1 U758 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2084), .A2(G2078), .ZN(n679) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U764 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U766 ( .A1(G108), .A2(G120), .ZN(n683) );
  NOR2_X1 U767 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G69), .A2(n684), .ZN(n856) );
  NAND2_X1 U769 ( .A1(G567), .A2(n856), .ZN(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT88), .ZN(n690) );
  NOR2_X1 U771 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U772 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U773 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G96), .A2(n688), .ZN(n857) );
  NAND2_X1 U775 ( .A1(G2106), .A2(n857), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(n691), .ZN(G319) );
  INV_X1 U778 ( .A(G319), .ZN(n693) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n855) );
  NAND2_X1 U781 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(n694), .A2(G40), .ZN(n696) );
  INV_X1 U783 ( .A(KEYINPUT90), .ZN(n695) );
  XNOR2_X2 U784 ( .A(n696), .B(n695), .ZN(n728) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n727) );
  INV_X1 U786 ( .A(n727), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n728), .A2(n697), .ZN(n725) );
  INV_X1 U788 ( .A(n725), .ZN(n843) );
  XNOR2_X1 U789 ( .A(G2067), .B(KEYINPUT37), .ZN(n841) );
  NAND2_X1 U790 ( .A1(G104), .A2(n896), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G140), .A2(n897), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U793 ( .A(KEYINPUT34), .B(n700), .ZN(n705) );
  NAND2_X1 U794 ( .A1(G116), .A2(n892), .ZN(n702) );
  NAND2_X1 U795 ( .A1(G128), .A2(n893), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U797 ( .A(KEYINPUT35), .B(n703), .Z(n704) );
  NOR2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U799 ( .A(KEYINPUT36), .B(n706), .ZN(n910) );
  NOR2_X1 U800 ( .A1(n841), .A2(n910), .ZN(n952) );
  NAND2_X1 U801 ( .A1(n843), .A2(n952), .ZN(n839) );
  NAND2_X1 U802 ( .A1(G95), .A2(n896), .ZN(n708) );
  NAND2_X1 U803 ( .A1(G131), .A2(n897), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U805 ( .A(KEYINPUT92), .B(n709), .Z(n711) );
  NAND2_X1 U806 ( .A1(n893), .A2(G119), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U808 ( .A1(G107), .A2(n892), .ZN(n712) );
  XNOR2_X1 U809 ( .A(KEYINPUT91), .B(n712), .ZN(n713) );
  NOR2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n906) );
  INV_X1 U811 ( .A(G1991), .ZN(n970) );
  NOR2_X1 U812 ( .A1(n906), .A2(n970), .ZN(n724) );
  NAND2_X1 U813 ( .A1(G105), .A2(n896), .ZN(n715) );
  XNOR2_X1 U814 ( .A(n715), .B(KEYINPUT38), .ZN(n722) );
  NAND2_X1 U815 ( .A1(G117), .A2(n892), .ZN(n717) );
  NAND2_X1 U816 ( .A1(G129), .A2(n893), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U818 ( .A1(G141), .A2(n897), .ZN(n718) );
  XNOR2_X1 U819 ( .A(KEYINPUT93), .B(n718), .ZN(n719) );
  NOR2_X1 U820 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U821 ( .A1(n722), .A2(n721), .ZN(n909) );
  AND2_X1 U822 ( .A1(n909), .A2(G1996), .ZN(n723) );
  NOR2_X1 U823 ( .A1(n724), .A2(n723), .ZN(n954) );
  NOR2_X1 U824 ( .A1(n954), .A2(n725), .ZN(n835) );
  INV_X1 U825 ( .A(n835), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n839), .A2(n726), .ZN(n830) );
  NAND2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X2 U828 ( .A(n729), .B(KEYINPUT64), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n778), .A2(G2084), .ZN(n790) );
  NOR2_X1 U830 ( .A1(n788), .A2(n790), .ZN(n730) );
  NAND2_X1 U831 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U832 ( .A(n731), .B(KEYINPUT30), .ZN(n732) );
  NOR2_X1 U833 ( .A1(G168), .A2(n732), .ZN(n733) );
  XNOR2_X1 U834 ( .A(n733), .B(KEYINPUT103), .ZN(n738) );
  XOR2_X1 U835 ( .A(G1961), .B(KEYINPUT94), .Z(n988) );
  NAND2_X1 U836 ( .A1(n778), .A2(n988), .ZN(n735) );
  XNOR2_X1 U837 ( .A(n742), .B(KEYINPUT95), .ZN(n760) );
  XNOR2_X1 U838 ( .A(KEYINPUT25), .B(G2078), .ZN(n973) );
  NAND2_X1 U839 ( .A1(n760), .A2(n973), .ZN(n734) );
  NAND2_X1 U840 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U841 ( .A(KEYINPUT96), .B(n736), .ZN(n773) );
  OR2_X1 U842 ( .A1(n773), .A2(G171), .ZN(n737) );
  NAND2_X1 U843 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U844 ( .A(n739), .B(KEYINPUT31), .ZN(n777) );
  NAND2_X1 U845 ( .A1(n742), .A2(G1341), .ZN(n740) );
  XNOR2_X1 U846 ( .A(n740), .B(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U847 ( .A1(n741), .A2(n1034), .ZN(n747) );
  INV_X1 U848 ( .A(KEYINPUT26), .ZN(n745) );
  INV_X1 U849 ( .A(n742), .ZN(n743) );
  NAND2_X1 U850 ( .A1(n743), .A2(G1996), .ZN(n744) );
  XNOR2_X1 U851 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U852 ( .A(n748), .B(KEYINPUT99), .ZN(n753) );
  NAND2_X1 U853 ( .A1(G2067), .A2(n760), .ZN(n749) );
  XNOR2_X1 U854 ( .A(n749), .B(KEYINPUT100), .ZN(n751) );
  NAND2_X1 U855 ( .A1(G1348), .A2(n778), .ZN(n750) );
  NAND2_X1 U856 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U857 ( .A1(n753), .A2(n752), .ZN(n757) );
  NOR2_X1 U858 ( .A1(n1029), .A2(n754), .ZN(n755) );
  XNOR2_X1 U859 ( .A(n755), .B(KEYINPUT101), .ZN(n756) );
  NAND2_X1 U860 ( .A1(n757), .A2(n756), .ZN(n764) );
  INV_X1 U861 ( .A(G299), .ZN(n1026) );
  NAND2_X1 U862 ( .A1(G2072), .A2(n760), .ZN(n758) );
  XNOR2_X1 U863 ( .A(n758), .B(KEYINPUT27), .ZN(n762) );
  INV_X1 U864 ( .A(G1956), .ZN(n759) );
  NOR2_X1 U865 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U866 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U867 ( .A1(n1026), .A2(n765), .ZN(n763) );
  NAND2_X1 U868 ( .A1(n764), .A2(n763), .ZN(n769) );
  NOR2_X1 U869 ( .A1(n1026), .A2(n765), .ZN(n767) );
  XNOR2_X1 U870 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n766) );
  XNOR2_X1 U871 ( .A(n767), .B(n766), .ZN(n768) );
  NAND2_X1 U872 ( .A1(n769), .A2(n768), .ZN(n772) );
  XNOR2_X1 U873 ( .A(n772), .B(n771), .ZN(n775) );
  NAND2_X1 U874 ( .A1(n773), .A2(G171), .ZN(n774) );
  NAND2_X1 U875 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U876 ( .A1(n777), .A2(n776), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n787), .A2(G286), .ZN(n783) );
  NOR2_X1 U878 ( .A1(G1971), .A2(n824), .ZN(n780) );
  NOR2_X1 U879 ( .A1(n778), .A2(G2090), .ZN(n779) );
  NOR2_X1 U880 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U881 ( .A1(n781), .A2(G303), .ZN(n782) );
  NAND2_X1 U882 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U883 ( .A1(n784), .A2(G8), .ZN(n785) );
  XNOR2_X1 U884 ( .A(KEYINPUT32), .B(n785), .ZN(n814) );
  INV_X1 U885 ( .A(KEYINPUT104), .ZN(n786) );
  XNOR2_X1 U886 ( .A(n787), .B(n786), .ZN(n789) );
  NAND2_X1 U887 ( .A1(G8), .A2(n790), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n815) );
  INV_X1 U889 ( .A(n824), .ZN(n793) );
  NAND2_X1 U890 ( .A1(G1976), .A2(G288), .ZN(n1022) );
  AND2_X1 U891 ( .A1(n793), .A2(n1022), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n814), .A2(n794), .ZN(n799) );
  INV_X1 U893 ( .A(n795), .ZN(n797) );
  NOR2_X1 U894 ( .A1(G1976), .A2(G288), .ZN(n806) );
  NOR2_X1 U895 ( .A1(G303), .A2(G1971), .ZN(n796) );
  NOR2_X1 U896 ( .A1(n806), .A2(n796), .ZN(n1023) );
  OR2_X1 U897 ( .A1(n797), .A2(n1023), .ZN(n798) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U899 ( .A(n800), .B(KEYINPUT65), .ZN(n802) );
  INV_X1 U900 ( .A(KEYINPUT105), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n824), .A2(n805), .ZN(n801) );
  NOR2_X1 U902 ( .A1(KEYINPUT33), .A2(n803), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n806), .A2(KEYINPUT33), .ZN(n804) );
  NAND2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n806), .A2(KEYINPUT105), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n824), .A2(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n813) );
  XOR2_X1 U909 ( .A(G1981), .B(KEYINPUT106), .Z(n812) );
  XNOR2_X1 U910 ( .A(G305), .B(n812), .ZN(n1037) );
  NAND2_X1 U911 ( .A1(n813), .A2(n1037), .ZN(n826) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n819) );
  NOR2_X1 U913 ( .A1(G303), .A2(G2090), .ZN(n816) );
  XOR2_X1 U914 ( .A(KEYINPUT107), .B(n816), .Z(n817) );
  NAND2_X1 U915 ( .A1(G8), .A2(n817), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n820), .B(KEYINPUT108), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n821), .A2(n824), .ZN(n825) );
  NOR2_X1 U919 ( .A1(G1981), .A2(G305), .ZN(n822) );
  XOR2_X1 U920 ( .A(n822), .B(KEYINPUT24), .Z(n823) );
  XNOR2_X1 U921 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(G1986), .B(G290), .ZN(n1025) );
  NAND2_X1 U923 ( .A1(n1025), .A2(n843), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n846) );
  NOR2_X1 U925 ( .A1(G1996), .A2(n909), .ZN(n940) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n833) );
  AND2_X1 U927 ( .A1(n970), .A2(n906), .ZN(n949) );
  NOR2_X1 U928 ( .A1(n833), .A2(n949), .ZN(n834) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT110), .ZN(n837) );
  NOR2_X1 U931 ( .A1(n940), .A2(n837), .ZN(n838) );
  XNOR2_X1 U932 ( .A(n838), .B(KEYINPUT39), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n842) );
  NAND2_X1 U934 ( .A1(n841), .A2(n910), .ZN(n958) );
  NAND2_X1 U935 ( .A1(n842), .A2(n958), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n844), .A2(n843), .ZN(n845) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(n848) );
  XOR2_X1 U938 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n847) );
  XNOR2_X1 U939 ( .A(n848), .B(n847), .ZN(G329) );
  NAND2_X1 U940 ( .A1(n849), .A2(G2106), .ZN(n850) );
  XNOR2_X1 U941 ( .A(n850), .B(KEYINPUT112), .ZN(G217) );
  NAND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n851) );
  XNOR2_X1 U943 ( .A(KEYINPUT113), .B(n851), .ZN(n852) );
  NAND2_X1 U944 ( .A1(n852), .A2(G661), .ZN(n853) );
  XNOR2_X1 U945 ( .A(KEYINPUT114), .B(n853), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n855), .A2(n854), .ZN(G188) );
  XNOR2_X1 U948 ( .A(G120), .B(KEYINPUT115), .ZN(G236) );
  INV_X1 U950 ( .A(G108), .ZN(G238) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  NOR2_X1 U952 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(G2096), .B(KEYINPUT43), .Z(n859) );
  XNOR2_X1 U955 ( .A(G2090), .B(G2678), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(n860), .B(KEYINPUT116), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U960 ( .A(KEYINPUT42), .B(G2100), .Z(n864) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U964 ( .A(G1976), .B(G1971), .Z(n868) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1961), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(n869), .B(KEYINPUT41), .Z(n871) );
  XNOR2_X1 U968 ( .A(G1966), .B(G1981), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U970 ( .A(G2474), .B(G1956), .Z(n873) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G100), .A2(n896), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G112), .A2(n892), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n878), .B(KEYINPUT117), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G136), .A2(n897), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n893), .A2(G124), .ZN(n881) );
  XOR2_X1 U981 ( .A(KEYINPUT44), .B(n881), .Z(n882) );
  NOR2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT118), .B(n884), .ZN(G162) );
  NAND2_X1 U984 ( .A1(G103), .A2(n896), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G139), .A2(n897), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G115), .A2(n892), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G127), .A2(n893), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n942) );
  NAND2_X1 U992 ( .A1(G118), .A2(n892), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U995 ( .A1(G106), .A2(n896), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G142), .A2(n897), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(KEYINPUT45), .B(n900), .Z(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n942), .B(n903), .Z(n904) );
  XNOR2_X1 U1001 ( .A(G162), .B(n904), .ZN(n905) );
  XOR2_X1 U1002 ( .A(n905), .B(n948), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G164), .B(n906), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n915) );
  XNOR2_X1 U1005 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n912) );
  XOR2_X1 U1006 ( .A(n910), .B(n909), .Z(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(G160), .B(n913), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1011 ( .A(G171), .B(n1034), .ZN(n921) );
  XOR2_X1 U1012 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n919) );
  XNOR2_X1 U1013 ( .A(n1029), .B(n917), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(n922), .B(G286), .ZN(n923) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n923), .ZN(G397) );
  XOR2_X1 U1018 ( .A(G2451), .B(G2430), .Z(n925) );
  XNOR2_X1 U1019 ( .A(G2438), .B(G2443), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n925), .B(n924), .ZN(n931) );
  XOR2_X1 U1021 ( .A(G2435), .B(G2454), .Z(n927) );
  XNOR2_X1 U1022 ( .A(G1348), .B(G1341), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n929) );
  XOR2_X1 U1024 ( .A(G2446), .B(G2427), .Z(n928) );
  XNOR2_X1 U1025 ( .A(n929), .B(n928), .ZN(n930) );
  XOR2_X1 U1026 ( .A(n931), .B(n930), .Z(n932) );
  NAND2_X1 U1027 ( .A1(G14), .A2(n932), .ZN(n938) );
  NAND2_X1 U1028 ( .A1(G319), .A2(n938), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(G227), .A2(G229), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT49), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(G395), .A2(G397), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(G225) );
  INV_X1 U1034 ( .A(G225), .ZN(G308) );
  INV_X1 U1035 ( .A(G69), .ZN(G235) );
  INV_X1 U1036 ( .A(n938), .ZN(G401) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n964) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT51), .B(n941), .Z(n947) );
  XOR2_X1 U1041 ( .A(G2072), .B(n942), .Z(n944) );
  XOR2_X1 U1042 ( .A(G164), .B(G2078), .Z(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT50), .B(n945), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n961) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT121), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G160), .B(G2084), .Z(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n957), .B(KEYINPUT122), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(KEYINPUT52), .B(n962), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n965), .A2(G29), .ZN(n1021) );
  XOR2_X1 U1058 ( .A(G2090), .B(G35), .Z(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(KEYINPUT125), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(G34), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G2084), .B(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n986) );
  XNOR2_X1 U1063 ( .A(n970), .B(G25), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n971), .A2(G28), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT123), .ZN(n983) );
  XNOR2_X1 U1066 ( .A(G27), .B(n973), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G2067), .B(G26), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G2072), .B(G33), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n981) );
  INV_X1 U1071 ( .A(G1996), .ZN(n978) );
  XOR2_X1 U1072 ( .A(G32), .B(n978), .Z(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1076 ( .A(KEYINPUT53), .B(n984), .Z(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n1013) );
  NAND2_X1 U1078 ( .A1(KEYINPUT55), .A2(n1013), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(G11), .A2(n987), .ZN(n1019) );
  XNOR2_X1 U1080 ( .A(G5), .B(n988), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n989), .B(KEYINPUT126), .ZN(n1002) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(G4), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1956), .B(G20), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G19), .B(G1341), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT127), .B(G1981), .Z(n995) );
  XNOR2_X1 U1089 ( .A(G6), .B(n995), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1091 ( .A(KEYINPUT60), .B(n998), .Z(n1000) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1971), .B(G22), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1005) );
  NAND2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(n1010), .B(KEYINPUT61), .ZN(n1012) );
  INV_X1 U1103 ( .A(G16), .ZN(n1011) );
  NAND2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1017) );
  INV_X1 U1105 ( .A(n1013), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1047) );
  XOR2_X1 U1111 ( .A(KEYINPUT56), .B(G16), .Z(n1045) );
  NAND2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1033) );
  XNOR2_X1 U1114 ( .A(n1026), .B(G1956), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(G1971), .A2(G303), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(G1348), .B(n1029), .Z(n1030) );
  NOR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1043) );
  XOR2_X1 U1120 ( .A(n1034), .B(G1341), .Z(n1036) );
  XOR2_X1 U1121 ( .A(G171), .B(G1961), .Z(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1041) );
  XNOR2_X1 U1123 ( .A(G1966), .B(G168), .ZN(n1038) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1125 ( .A(n1039), .B(KEYINPUT57), .ZN(n1040) );
  NAND2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NOR2_X1 U1127 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NOR2_X1 U1128 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NOR2_X1 U1129 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1130 ( .A(n1048), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1131 ( .A(G311), .ZN(G150) );
  INV_X1 U1132 ( .A(G303), .ZN(G166) );
endmodule

