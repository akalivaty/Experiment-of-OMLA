

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G2104), .A2(n552), .ZN(n880) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n522), .Z(n877) );
  AND2_X1 U553 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X1 U554 ( .A1(n920), .A2(n814), .ZN(n519) );
  NOR2_X1 U555 ( .A1(n802), .A2(n519), .ZN(n520) );
  XNOR2_X1 U556 ( .A(KEYINPUT99), .B(n769), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n688), .A2(n771), .ZN(n730) );
  NAND2_X1 U558 ( .A1(G8), .A2(n730), .ZN(n763) );
  OR2_X1 U559 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U560 ( .A(n535), .B(KEYINPUT65), .ZN(G160) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  NAND2_X1 U562 ( .A1(G137), .A2(n877), .ZN(n525) );
  NAND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X1 U564 ( .A(KEYINPUT68), .B(n523), .Z(n881) );
  NAND2_X1 U565 ( .A1(G113), .A2(n881), .ZN(n524) );
  NAND2_X1 U566 ( .A1(n525), .A2(n524), .ZN(n534) );
  INV_X1 U567 ( .A(G2105), .ZN(n552) );
  NAND2_X1 U568 ( .A1(G125), .A2(n880), .ZN(n530) );
  AND2_X1 U569 ( .A1(G2104), .A2(G101), .ZN(n526) );
  NAND2_X1 U570 ( .A1(n526), .A2(n552), .ZN(n527) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n527), .Z(n528) );
  XNOR2_X1 U572 ( .A(n528), .B(KEYINPUT66), .ZN(n529) );
  NAND2_X1 U573 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U574 ( .A(KEYINPUT67), .ZN(n531) );
  XNOR2_X1 U575 ( .A(n532), .B(n531), .ZN(n533) );
  AND2_X1 U576 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U577 ( .A(G57), .ZN(G237) );
  INV_X1 U578 ( .A(G69), .ZN(G235) );
  INV_X1 U579 ( .A(G108), .ZN(G238) );
  INV_X1 U580 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U581 ( .A(G651), .B(KEYINPUT69), .ZN(n543) );
  NOR2_X1 U582 ( .A1(G543), .A2(n543), .ZN(n536) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n536), .Z(n648) );
  NAND2_X1 U584 ( .A1(n648), .A2(G63), .ZN(n537) );
  XNOR2_X1 U585 ( .A(n537), .B(KEYINPUT78), .ZN(n540) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  NOR2_X1 U587 ( .A1(G651), .A2(n636), .ZN(n538) );
  XNOR2_X1 U588 ( .A(KEYINPUT64), .B(n538), .ZN(n649) );
  NAND2_X1 U589 ( .A1(G51), .A2(n649), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U591 ( .A(KEYINPUT6), .B(n541), .ZN(n550) );
  NOR2_X1 U592 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U593 ( .A1(n644), .A2(G89), .ZN(n542) );
  XNOR2_X1 U594 ( .A(n542), .B(KEYINPUT4), .ZN(n546) );
  NOR2_X1 U595 ( .A1(n636), .A2(n543), .ZN(n544) );
  XNOR2_X1 U596 ( .A(KEYINPUT70), .B(n544), .ZN(n645) );
  NAND2_X1 U597 ( .A1(G76), .A2(n645), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U599 ( .A(KEYINPUT5), .B(n547), .ZN(n548) );
  XNOR2_X1 U600 ( .A(KEYINPUT77), .B(n548), .ZN(n549) );
  NOR2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U602 ( .A(KEYINPUT7), .B(n551), .Z(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U604 ( .A1(n552), .A2(G2104), .ZN(n876) );
  NAND2_X1 U605 ( .A1(G102), .A2(n876), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G138), .A2(n877), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U608 ( .A1(G126), .A2(n880), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G114), .A2(n881), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U611 ( .A1(n558), .A2(n557), .ZN(G164) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U614 ( .A(G223), .ZN(n819) );
  NAND2_X1 U615 ( .A1(n819), .A2(G567), .ZN(n560) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  XOR2_X1 U617 ( .A(G860), .B(KEYINPUT76), .Z(n599) );
  NAND2_X1 U618 ( .A1(n644), .A2(G81), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G68), .A2(n645), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT13), .B(n564), .Z(n568) );
  NAND2_X1 U623 ( .A1(G56), .A2(n648), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT75), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT14), .ZN(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G43), .A2(n649), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n915) );
  OR2_X1 U629 ( .A1(n599), .A2(n915), .ZN(G153) );
  NAND2_X1 U630 ( .A1(G90), .A2(n644), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G77), .A2(n645), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT9), .B(KEYINPUT72), .Z(n573) );
  XNOR2_X1 U634 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G64), .A2(n648), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G52), .A2(n649), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U638 ( .A(KEYINPUT71), .B(n577), .Z(n578) );
  NOR2_X1 U639 ( .A1(n579), .A2(n578), .ZN(G171) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U642 ( .A1(G66), .A2(n648), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G54), .A2(n649), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G92), .A2(n644), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G79), .A2(n645), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U649 ( .A(n586), .B(KEYINPUT15), .ZN(n914) );
  INV_X1 U650 ( .A(G868), .ZN(n663) );
  NAND2_X1 U651 ( .A1(n914), .A2(n663), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U653 ( .A1(n649), .A2(G53), .ZN(n595) );
  NAND2_X1 U654 ( .A1(G91), .A2(n644), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G65), .A2(n648), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G78), .A2(n645), .ZN(n591) );
  XNOR2_X1 U658 ( .A(KEYINPUT73), .B(n591), .ZN(n592) );
  NOR2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n596), .B(KEYINPUT74), .ZN(G299) );
  NOR2_X1 U662 ( .A1(G286), .A2(n663), .ZN(n598) );
  NOR2_X1 U663 ( .A1(G299), .A2(G868), .ZN(n597) );
  NOR2_X1 U664 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U666 ( .A(n914), .ZN(n642) );
  NAND2_X1 U667 ( .A1(n600), .A2(n642), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n915), .ZN(n604) );
  NAND2_X1 U670 ( .A1(n642), .A2(G868), .ZN(n602) );
  NOR2_X1 U671 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U672 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G99), .A2(n876), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT80), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n881), .A2(G111), .ZN(n606) );
  XOR2_X1 U676 ( .A(KEYINPUT79), .B(n606), .Z(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G123), .A2(n880), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n877), .A2(G135), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n983) );
  XNOR2_X1 U683 ( .A(G2096), .B(n983), .ZN(n615) );
  INV_X1 U684 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G86), .A2(n644), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G61), .A2(n648), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n645), .A2(G73), .ZN(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT2), .B(n618), .Z(n619) );
  NOR2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G48), .A2(n649), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(G305) );
  NAND2_X1 U694 ( .A1(G88), .A2(n644), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G50), .A2(n649), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n648), .A2(G62), .ZN(n625) );
  XOR2_X1 U698 ( .A(KEYINPUT82), .B(n625), .Z(n626) );
  NOR2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G75), .A2(n645), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(G303) );
  INV_X1 U702 ( .A(G303), .ZN(G166) );
  AND2_X1 U703 ( .A1(G72), .A2(n645), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G85), .A2(n644), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G47), .A2(n649), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n648), .A2(G60), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U710 ( .A1(G87), .A2(n636), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n648), .A2(n639), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G49), .A2(n649), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G559), .A2(n642), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n915), .B(n643), .ZN(n829) );
  NAND2_X1 U718 ( .A1(G93), .A2(n644), .ZN(n647) );
  NAND2_X1 U719 ( .A1(G80), .A2(n645), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n653) );
  NAND2_X1 U721 ( .A1(G67), .A2(n648), .ZN(n651) );
  NAND2_X1 U722 ( .A1(G55), .A2(n649), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U725 ( .A(KEYINPUT81), .B(n654), .ZN(n831) );
  XOR2_X1 U726 ( .A(G305), .B(n831), .Z(n656) );
  XNOR2_X1 U727 ( .A(G299), .B(G166), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(G290), .ZN(n660) );
  XNOR2_X1 U730 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n893) );
  XOR2_X1 U733 ( .A(n893), .B(KEYINPUT84), .Z(n661) );
  XOR2_X1 U734 ( .A(n829), .B(n661), .Z(n662) );
  NAND2_X1 U735 ( .A1(n662), .A2(G868), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n663), .A2(n831), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U744 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n671) );
  NAND2_X1 U745 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n672), .A2(G218), .ZN(n673) );
  NAND2_X1 U748 ( .A1(G96), .A2(n673), .ZN(n827) );
  NAND2_X1 U749 ( .A1(n827), .A2(G2106), .ZN(n678) );
  NOR2_X1 U750 ( .A1(G236), .A2(G238), .ZN(n675) );
  NOR2_X1 U751 ( .A1(G235), .A2(G237), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U753 ( .A(KEYINPUT86), .B(n676), .ZN(n826) );
  NAND2_X1 U754 ( .A1(n826), .A2(G567), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n832) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U757 ( .A1(n832), .A2(n679), .ZN(n823) );
  NAND2_X1 U758 ( .A1(n823), .A2(G36), .ZN(G176) );
  NOR2_X1 U759 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X1 U760 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U761 ( .A(n770), .ZN(n688) );
  AND2_X1 U762 ( .A1(n771), .A2(n688), .ZN(n705) );
  NAND2_X1 U763 ( .A1(n705), .A2(G2072), .ZN(n680) );
  XNOR2_X1 U764 ( .A(n680), .B(KEYINPUT27), .ZN(n682) );
  INV_X1 U765 ( .A(G1956), .ZN(n947) );
  NOR2_X1 U766 ( .A1(n947), .A2(n705), .ZN(n681) );
  NOR2_X1 U767 ( .A1(n682), .A2(n681), .ZN(n684) );
  INV_X1 U768 ( .A(G299), .ZN(n921) );
  NOR2_X1 U769 ( .A1(n684), .A2(n921), .ZN(n683) );
  XOR2_X1 U770 ( .A(n683), .B(KEYINPUT28), .Z(n703) );
  NAND2_X1 U771 ( .A1(n684), .A2(n921), .ZN(n701) );
  AND2_X1 U772 ( .A1(n771), .A2(G1996), .ZN(n685) );
  AND2_X1 U773 ( .A1(n685), .A2(n688), .ZN(n687) );
  XOR2_X1 U774 ( .A(KEYINPUT26), .B(KEYINPUT92), .Z(n686) );
  XNOR2_X1 U775 ( .A(n687), .B(n686), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n730), .A2(G1341), .ZN(n689) );
  NAND2_X1 U777 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U778 ( .A(n691), .B(KEYINPUT93), .ZN(n696) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n730), .ZN(n693) );
  NAND2_X1 U780 ( .A1(G2067), .A2(n705), .ZN(n692) );
  NAND2_X1 U781 ( .A1(n693), .A2(n692), .ZN(n697) );
  AND2_X1 U782 ( .A1(n697), .A2(n914), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n915), .A2(n694), .ZN(n695) );
  AND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U785 ( .A1(n697), .A2(n914), .ZN(n698) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U787 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U789 ( .A(n704), .B(KEYINPUT29), .ZN(n709) );
  NAND2_X1 U790 ( .A1(G1961), .A2(n730), .ZN(n707) );
  XOR2_X1 U791 ( .A(G2078), .B(KEYINPUT25), .Z(n1015) );
  NAND2_X1 U792 ( .A1(n705), .A2(n1015), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U794 ( .A1(G301), .A2(n710), .ZN(n708) );
  NOR2_X1 U795 ( .A1(n709), .A2(n708), .ZN(n721) );
  AND2_X1 U796 ( .A1(G301), .A2(n710), .ZN(n718) );
  NOR2_X1 U797 ( .A1(n763), .A2(G1966), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(KEYINPUT91), .ZN(n723) );
  INV_X1 U799 ( .A(G8), .ZN(n712) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n730), .ZN(n724) );
  NOR2_X1 U801 ( .A1(n712), .A2(n724), .ZN(n713) );
  AND2_X1 U802 ( .A1(n723), .A2(n713), .ZN(n715) );
  XOR2_X1 U803 ( .A(KEYINPUT94), .B(KEYINPUT30), .Z(n714) );
  XNOR2_X1 U804 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U805 ( .A1(G168), .A2(n716), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U807 ( .A(n719), .B(KEYINPUT31), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U809 ( .A(n722), .B(KEYINPUT95), .ZN(n729) );
  AND2_X1 U810 ( .A1(n729), .A2(n723), .ZN(n726) );
  NAND2_X1 U811 ( .A1(G8), .A2(n724), .ZN(n725) );
  NAND2_X1 U812 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U813 ( .A(n727), .B(KEYINPUT96), .ZN(n740) );
  AND2_X1 U814 ( .A1(G286), .A2(G8), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n737) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n730), .ZN(n731) );
  XNOR2_X1 U817 ( .A(KEYINPUT97), .B(n731), .ZN(n734) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n763), .ZN(n732) );
  NOR2_X1 U819 ( .A1(G166), .A2(n732), .ZN(n733) );
  NAND2_X1 U820 ( .A1(n734), .A2(n733), .ZN(n735) );
  OR2_X1 U821 ( .A1(n712), .A2(n735), .ZN(n736) );
  AND2_X1 U822 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U823 ( .A(n738), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U824 ( .A1(n740), .A2(n739), .ZN(n762) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n742) );
  NOR2_X1 U826 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n925) );
  NAND2_X1 U828 ( .A1(n742), .A2(KEYINPUT33), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n743), .A2(n763), .ZN(n745) );
  XOR2_X1 U830 ( .A(G1981), .B(G305), .Z(n932) );
  INV_X1 U831 ( .A(n932), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n749) );
  AND2_X1 U833 ( .A1(n749), .A2(KEYINPUT33), .ZN(n752) );
  INV_X1 U834 ( .A(n752), .ZN(n746) );
  AND2_X1 U835 ( .A1(n925), .A2(n746), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n762), .A2(n747), .ZN(n754) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n924) );
  INV_X1 U838 ( .A(n924), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n763), .A2(n748), .ZN(n750) );
  AND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  OR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n768) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U844 ( .A1(G8), .A2(n755), .ZN(n756) );
  XNOR2_X1 U845 ( .A(n756), .B(KEYINPUT98), .ZN(n760) );
  NOR2_X1 U846 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XOR2_X1 U847 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  NOR2_X1 U848 ( .A1(n763), .A2(n758), .ZN(n764) );
  INV_X1 U849 ( .A(n764), .ZN(n759) );
  AND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n766) );
  OR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n771), .A2(n770), .ZN(n814) );
  NAND2_X1 U855 ( .A1(G104), .A2(n876), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G140), .A2(n877), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U858 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U859 ( .A1(G128), .A2(n880), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G116), .A2(n881), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U862 ( .A(n777), .B(KEYINPUT35), .Z(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U864 ( .A(KEYINPUT36), .B(n780), .Z(n781) );
  XNOR2_X1 U865 ( .A(KEYINPUT88), .B(n781), .ZN(n887) );
  XOR2_X1 U866 ( .A(KEYINPUT37), .B(G2067), .Z(n811) );
  AND2_X1 U867 ( .A1(n887), .A2(n811), .ZN(n989) );
  NAND2_X1 U868 ( .A1(n814), .A2(n989), .ZN(n809) );
  NAND2_X1 U869 ( .A1(n881), .A2(G107), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n782), .B(KEYINPUT90), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G95), .A2(n876), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G131), .A2(n877), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G119), .A2(n880), .ZN(n785) );
  XNOR2_X1 U875 ( .A(KEYINPUT89), .B(n785), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n863) );
  AND2_X1 U878 ( .A1(n863), .A2(G1991), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G129), .A2(n880), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G117), .A2(n881), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n876), .A2(G105), .ZN(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n877), .A2(G141), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n864) );
  AND2_X1 U887 ( .A1(n864), .A2(G1996), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n981) );
  INV_X1 U889 ( .A(n814), .ZN(n799) );
  NOR2_X1 U890 ( .A1(n981), .A2(n799), .ZN(n806) );
  INV_X1 U891 ( .A(n806), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n809), .A2(n800), .ZN(n802) );
  XOR2_X1 U893 ( .A(G1986), .B(KEYINPUT87), .Z(n801) );
  XNOR2_X1 U894 ( .A(G290), .B(n801), .ZN(n920) );
  NAND2_X1 U895 ( .A1(n521), .A2(n520), .ZN(n817) );
  NOR2_X1 U896 ( .A1(n864), .A2(G1996), .ZN(n803) );
  XNOR2_X1 U897 ( .A(n803), .B(KEYINPUT100), .ZN(n978) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n863), .ZN(n984) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n984), .A2(n804), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n978), .A2(n807), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n887), .A2(n811), .ZN(n812) );
  XNOR2_X1 U906 ( .A(n812), .B(KEYINPUT101), .ZN(n992) );
  NAND2_X1 U907 ( .A1(n813), .A2(n992), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n819), .ZN(G217) );
  NAND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n821) );
  INV_X1 U913 ( .A(G661), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G1), .A2(G3), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n825), .B(KEYINPUT104), .ZN(G188) );
  INV_X1 U920 ( .A(G132), .ZN(G219) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G82), .ZN(G220) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n828), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U925 ( .A(G261), .ZN(G325) );
  NOR2_X1 U926 ( .A1(G860), .A2(n829), .ZN(n830) );
  XOR2_X1 U927 ( .A(n831), .B(n830), .Z(G145) );
  INV_X1 U928 ( .A(n832), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT108), .B(G2678), .Z(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT43), .B(G2096), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(n835), .B(KEYINPUT107), .Z(n837) );
  XNOR2_X1 U933 ( .A(G2078), .B(G2072), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(G2100), .B(G2090), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2084), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1981), .B(G1956), .Z(n845) );
  XNOR2_X1 U942 ( .A(G1966), .B(G1961), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n846), .B(G2474), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1971), .B(G1976), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(KEYINPUT41), .B(G1986), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U951 ( .A1(n880), .A2(G124), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G112), .A2(n881), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G100), .A2(n876), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G136), .A2(n877), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n861) );
  XNOR2_X1 U960 ( .A(G164), .B(n983), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U962 ( .A(n862), .B(G162), .Z(n866) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n875) );
  NAND2_X1 U965 ( .A1(G130), .A2(n880), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G118), .A2(n881), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U968 ( .A1(G106), .A2(n876), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G142), .A2(n877), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(KEYINPUT45), .B(n871), .Z(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U973 ( .A(n875), .B(n874), .Z(n889) );
  NAND2_X1 U974 ( .A1(G103), .A2(n876), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G139), .A2(n877), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U977 ( .A1(G127), .A2(n880), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G115), .A2(n881), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n972) );
  XOR2_X1 U982 ( .A(n887), .B(n972), .Z(n888) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U984 ( .A(G160), .B(n890), .Z(n891) );
  NOR2_X1 U985 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U986 ( .A(G286), .B(n914), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n892), .B(n915), .ZN(n895) );
  XOR2_X1 U988 ( .A(G301), .B(n893), .Z(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U991 ( .A(KEYINPUT102), .B(G2446), .Z(n898) );
  XNOR2_X1 U992 ( .A(G2443), .B(G2454), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(n899), .B(G2451), .Z(n901) );
  XNOR2_X1 U995 ( .A(G1348), .B(G1341), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U997 ( .A(G2435), .B(G2427), .Z(n903) );
  XNOR2_X1 U998 ( .A(G2430), .B(G2438), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n906), .ZN(n912) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n912), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(n912), .ZN(G401) );
  XNOR2_X1 U1010 ( .A(G16), .B(KEYINPUT56), .ZN(n939) );
  XOR2_X1 U1011 ( .A(G1348), .B(KEYINPUT119), .Z(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(G1341), .B(n915), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n937) );
  XNOR2_X1 U1015 ( .A(G1961), .B(KEYINPUT120), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(G301), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n929) );
  XNOR2_X1 U1018 ( .A(n921), .B(G1956), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(G1971), .A2(G303), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n935) );
  XNOR2_X1 U1024 ( .A(G1966), .B(G168), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(n930), .B(KEYINPUT118), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1027 ( .A(KEYINPUT57), .B(n933), .Z(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n970) );
  INV_X1 U1031 ( .A(G16), .ZN(n968) );
  XNOR2_X1 U1032 ( .A(G1986), .B(G24), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(G1971), .B(G22), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(G1976), .B(G23), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT125), .B(n942), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT126), .B(n945), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(n946), .B(KEYINPUT58), .ZN(n962) );
  XNOR2_X1 U1040 ( .A(G20), .B(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(G1981), .B(G6), .Z(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G19), .B(G1341), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(KEYINPUT122), .B(n952), .ZN(n956) );
  XOR2_X1 U1046 ( .A(KEYINPUT123), .B(G4), .Z(n954) );
  XNOR2_X1 U1047 ( .A(G1348), .B(KEYINPUT59), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n954), .B(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT60), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G1966), .B(KEYINPUT124), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G21), .B(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1055 ( .A(KEYINPUT121), .B(G1961), .Z(n963) );
  XNOR2_X1 U1056 ( .A(G5), .B(n963), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT61), .B(n966), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n971), .B(KEYINPUT127), .ZN(n1003) );
  XOR2_X1 U1062 ( .A(G2072), .B(n972), .Z(n974) );
  XOR2_X1 U1063 ( .A(G164), .B(G2078), .Z(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(n975), .B(KEYINPUT113), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n976), .B(KEYINPUT50), .ZN(n997) );
  XOR2_X1 U1067 ( .A(G2090), .B(G162), .Z(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n979), .B(KEYINPUT51), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n980), .B(KEYINPUT111), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n994) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1073 ( .A(KEYINPUT109), .B(n985), .Z(n987) );
  XNOR2_X1 U1074 ( .A(G160), .B(G2084), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(n990), .B(KEYINPUT110), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1080 ( .A(KEYINPUT112), .B(n995), .Z(n996) );
  NOR2_X1 U1081 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1082 ( .A(KEYINPUT52), .B(n998), .Z(n999) );
  NOR2_X1 U1083 ( .A1(KEYINPUT55), .A2(n999), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(KEYINPUT114), .B(n1000), .Z(n1001) );
  NAND2_X1 U1085 ( .A1(n1001), .A2(G29), .ZN(n1002) );
  NAND2_X1 U1086 ( .A1(n1003), .A2(n1002), .ZN(n1028) );
  XOR2_X1 U1087 ( .A(G2090), .B(G35), .Z(n1006) );
  XOR2_X1 U1088 ( .A(KEYINPUT54), .B(G34), .Z(n1004) );
  XNOR2_X1 U1089 ( .A(n1004), .B(G2084), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1021) );
  XNOR2_X1 U1091 ( .A(G2067), .B(G26), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G32), .B(G1996), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1014) );
  XOR2_X1 U1094 ( .A(G2072), .B(G33), .Z(n1009) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(G28), .ZN(n1012) );
  XOR2_X1 U1096 ( .A(G25), .B(G1991), .Z(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT115), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(G27), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT53), .B(n1018), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(KEYINPUT116), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(KEYINPUT55), .B(n1022), .ZN(n1024) );
  INV_X1 U1106 ( .A(G29), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(G11), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(KEYINPUT117), .B(n1026), .Z(n1027) );
  NOR2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1029), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

