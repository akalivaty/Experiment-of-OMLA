//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n438, new_n443, new_n444, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n651,
    new_n652, new_n653, new_n656, new_n658, new_n659, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G96), .Z(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  AND2_X1   g017(.A1(KEYINPUT66), .A2(G108), .ZN(new_n443));
  NOR2_X1   g018(.A1(KEYINPUT66), .A2(G108), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(G238));
  NAND4_X1  g020(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g028(.A1(G237), .A2(G235), .A3(G236), .ZN(new_n454));
  OAI21_X1  g029(.A(new_n454), .B1(new_n444), .B2(new_n443), .ZN(new_n455));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g033(.A1(new_n436), .A2(new_n438), .A3(G44), .A4(G132), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT2), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  AND3_X1   g037(.A1(new_n460), .A2(KEYINPUT68), .A3(G2106), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n458), .A2(G567), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT68), .B1(new_n460), .B2(G2106), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NOR3_X1   g054(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT69), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  OR2_X1    g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(new_n467), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(KEYINPUT70), .A3(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n485), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G136), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  NAND2_X1  g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n482), .B2(new_n483), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n467), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n505), .B(new_n507), .C1(new_n469), .C2(new_n468), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT3), .B(G2104), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n510), .B2(new_n505), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n503), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(G88), .B1(new_n520), .B2(G50), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT72), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n514), .B2(new_n515), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(KEYINPUT73), .B(G651), .C1(new_n524), .C2(new_n526), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n522), .B1(new_n529), .B2(new_n530), .ZN(G166));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n514), .A2(new_n515), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n520), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT76), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n542), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT7), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n546), .A3(new_n543), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n539), .A2(KEYINPUT75), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(KEYINPUT5), .A2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(KEYINPUT5), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n538), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(KEYINPUT6), .A2(G651), .ZN(new_n552));
  NOR2_X1   g127(.A1(KEYINPUT6), .A2(G651), .ZN(new_n553));
  OAI21_X1  g128(.A(G543), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(G51), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(new_n557), .B1(G89), .B2(new_n518), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n548), .A2(new_n558), .ZN(G286));
  INV_X1    g134(.A(G286), .ZN(G168));
  OAI22_X1  g135(.A1(new_n550), .A2(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n561));
  INV_X1    g136(.A(G90), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT77), .B(G52), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n561), .A2(new_n562), .B1(new_n554), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G651), .ZN(new_n565));
  OAI21_X1  g140(.A(G64), .B1(new_n549), .B2(new_n550), .ZN(new_n566));
  NAND2_X1  g141(.A1(G77), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n564), .A2(new_n568), .ZN(G171));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  INV_X1    g145(.A(G56), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n514), .B2(new_n515), .ZN(new_n572));
  NAND2_X1  g147(.A1(G68), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n549), .A2(new_n550), .ZN(new_n576));
  OAI211_X1 g151(.A(KEYINPUT78), .B(new_n573), .C1(new_n576), .C2(new_n571), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(G651), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n518), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G860), .ZN(G153));
  NAND4_X1  g157(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g158(.A1(G1), .A2(G3), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT8), .ZN(new_n585));
  NAND4_X1  g160(.A1(G319), .A2(G483), .A3(G661), .A4(new_n585), .ZN(G188));
  INV_X1    g161(.A(G78), .ZN(new_n587));
  OR3_X1    g162(.A1(new_n587), .A2(new_n519), .A3(KEYINPUT79), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT79), .B1(new_n587), .B2(new_n519), .ZN(new_n589));
  INV_X1    g164(.A(G65), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n576), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G91), .B2(new_n518), .ZN(new_n592));
  INV_X1    g167(.A(G53), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n554), .A2(KEYINPUT9), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT9), .B1(new_n554), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(G299));
  NAND2_X1  g172(.A1(new_n516), .A2(new_n517), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n537), .A2(new_n598), .A3(G90), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT77), .B(G52), .Z(new_n600));
  NAND2_X1  g175(.A1(new_n520), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n567), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n537), .B2(G64), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n599), .B(new_n601), .C1(new_n603), .C2(new_n565), .ZN(G301));
  NAND2_X1  g179(.A1(new_n529), .A2(new_n530), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n521), .ZN(G303));
  NOR3_X1   g181(.A1(new_n549), .A2(new_n550), .A3(G74), .ZN(new_n607));
  INV_X1    g182(.A(G49), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n607), .A2(new_n565), .B1(new_n554), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G87), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n561), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT80), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n537), .B2(G74), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n520), .A2(G49), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n537), .A2(new_n598), .A3(G87), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(G288));
  INV_X1    g194(.A(G86), .ZN(new_n620));
  INV_X1    g195(.A(G48), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n561), .A2(new_n620), .B1(new_n554), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n624));
  OAI21_X1  g199(.A(G61), .B1(new_n549), .B2(new_n550), .ZN(new_n625));
  NAND2_X1  g200(.A1(G73), .A2(G543), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n627), .B2(G651), .ZN(new_n628));
  AOI211_X1 g203(.A(KEYINPUT81), .B(new_n565), .C1(new_n625), .C2(new_n626), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(G305));
  AOI22_X1  g205(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(new_n565), .ZN(new_n632));
  INV_X1    g207(.A(G85), .ZN(new_n633));
  INV_X1    g208(.A(G47), .ZN(new_n634));
  OAI22_X1  g209(.A1(new_n561), .A2(new_n633), .B1(new_n554), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G290));
  NAND2_X1  g212(.A1(G301), .A2(G868), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT10), .ZN(new_n640));
  INV_X1    g215(.A(G92), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n561), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(G79), .A2(G543), .ZN(new_n644));
  INV_X1    g219(.A(G66), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n576), .B2(new_n645), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n646), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n638), .B1(new_n648), .B2(G868), .ZN(G284));
  OAI21_X1  g224(.A(new_n638), .B1(new_n648), .B2(G868), .ZN(G321));
  INV_X1    g225(.A(G868), .ZN(new_n651));
  NOR2_X1   g226(.A1(G286), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G299), .B(KEYINPUT82), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n651), .ZN(G297));
  AOI21_X1  g229(.A(new_n652), .B1(new_n653), .B2(new_n651), .ZN(G280));
  INV_X1    g230(.A(G559), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n648), .B1(new_n656), .B2(G860), .ZN(G148));
  NAND2_X1  g232(.A1(new_n648), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G868), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(G868), .B2(new_n581), .ZN(G323));
  XNOR2_X1  g235(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g236(.A1(new_n510), .A2(new_n474), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT13), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n494), .A2(G135), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n486), .A2(G123), .ZN(new_n667));
  OR2_X1    g242(.A1(G99), .A2(G2105), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n668), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G2096), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(G2096), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n665), .A2(new_n673), .A3(new_n674), .ZN(G156));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT15), .B(G2435), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(G2438), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2427), .B(G2430), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n682), .A3(new_n680), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(KEYINPUT14), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1341), .B(G1348), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2451), .B(G2454), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT16), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(KEYINPUT16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(new_n687), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n686), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G2443), .B(G2446), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n681), .B2(new_n683), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n695), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n701), .A3(new_n685), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n697), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G14), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n698), .B1(new_n697), .B2(new_n702), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n676), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n697), .A2(new_n702), .ZN(new_n707));
  INV_X1    g282(.A(new_n698), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n709), .A2(KEYINPUT84), .A3(G14), .A4(new_n703), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(G401));
  XOR2_X1   g286(.A(G2072), .B(G2078), .Z(new_n712));
  XOR2_X1   g287(.A(G2084), .B(G2090), .Z(new_n713));
  XNOR2_X1  g288(.A(G2067), .B(G2678), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n712), .B1(new_n715), .B2(KEYINPUT18), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(new_n672), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(KEYINPUT17), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n713), .A2(new_n714), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2100), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(G2100), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n724), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n716), .B(G2096), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(new_n727), .A3(new_n722), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(G227));
  XNOR2_X1  g305(.A(G1981), .B(G1986), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(G1956), .B(G2474), .ZN(new_n735));
  XNOR2_X1  g310(.A(G1961), .B(G1966), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1971), .ZN(new_n740));
  INV_X1    g315(.A(G1976), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G1971), .A2(G1976), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT19), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n742), .A2(KEYINPUT19), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n739), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n748), .A2(new_n737), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n748), .B2(new_n737), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n748), .A2(new_n755), .A3(new_n738), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n748), .B2(new_n738), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n734), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n748), .A2(new_n737), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(KEYINPUT85), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n748), .A2(new_n737), .A3(new_n751), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n748), .A2(new_n738), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT20), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n748), .A2(new_n755), .A3(new_n738), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n763), .A2(new_n767), .A3(new_n750), .A4(new_n733), .ZN(new_n768));
  XOR2_X1   g343(.A(G1991), .B(G1996), .Z(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n759), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n759), .B2(new_n768), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n732), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n759), .A2(new_n768), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(new_n769), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n759), .A2(new_n768), .A3(new_n770), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n775), .A2(new_n731), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(G229));
  AOI22_X1  g354(.A1(new_n537), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT81), .B1(new_n780), .B2(new_n565), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n627), .A2(new_n624), .A3(G651), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n622), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G16), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G6), .B2(new_n784), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(G22), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT86), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n784), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1971), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G1971), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n784), .A2(G23), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n795), .B1(new_n797), .B2(new_n784), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n786), .B2(new_n787), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n494), .A2(G131), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n486), .A2(G119), .ZN(new_n805));
  OR2_X1    g380(.A1(G95), .A2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n806), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G25), .B2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n784), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n636), .B2(new_n784), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1986), .Z(new_n817));
  NAND4_X1  g392(.A1(new_n803), .A2(new_n813), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G4), .A2(G16), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n648), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT87), .B(G1348), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n581), .A2(new_n784), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n784), .B2(G19), .ZN(new_n827));
  INV_X1    g402(.A(G1341), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n824), .A2(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT27), .B(G1996), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT93), .ZN(new_n831));
  OAI211_X1 g406(.A(G141), .B(new_n467), .C1(new_n480), .C2(new_n484), .ZN(new_n832));
  OAI211_X1 g407(.A(G129), .B(G2105), .C1(new_n480), .C2(new_n484), .ZN(new_n833));
  NAND3_X1  g408(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT26), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n836), .A2(new_n837), .B1(G105), .B2(new_n474), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n832), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G29), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(G32), .ZN(new_n843));
  OAI221_X1 g418(.A(new_n829), .B1(new_n828), .B2(new_n827), .C1(new_n831), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(G171), .A2(new_n784), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G5), .B2(new_n784), .ZN(new_n846));
  INV_X1    g421(.A(G1961), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT24), .ZN(new_n848));
  INV_X1    g423(.A(G34), .ZN(new_n849));
  AOI21_X1  g424(.A(G29), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G160), .B2(new_n841), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n846), .A2(new_n847), .B1(G2084), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(new_n847), .ZN(new_n854));
  INV_X1    g429(.A(G2078), .ZN(new_n855));
  NOR2_X1   g430(.A1(G164), .A2(new_n841), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G27), .B2(new_n841), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G1966), .ZN(new_n859));
  NAND2_X1  g434(.A1(G286), .A2(G16), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n784), .A2(G21), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI211_X1 g437(.A(new_n853), .B(new_n858), .C1(new_n859), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n784), .A2(G20), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT23), .Z(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G299), .B2(G16), .ZN(new_n866));
  INV_X1    g441(.A(G1956), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n862), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(G1966), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n857), .A2(new_n855), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n670), .A2(new_n841), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT95), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT31), .B(G11), .Z(new_n874));
  INV_X1    g449(.A(G28), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(KEYINPUT30), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT96), .Z(new_n877));
  AOI21_X1  g452(.A(G29), .B1(new_n875), .B2(KEYINPUT30), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n841), .A2(G26), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(G140), .B(new_n467), .C1(new_n480), .C2(new_n484), .ZN(new_n884));
  OAI211_X1 g459(.A(G128), .B(G2105), .C1(new_n480), .C2(new_n484), .ZN(new_n885));
  OR2_X1    g460(.A1(G104), .A2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n883), .B1(new_n888), .B2(G29), .ZN(new_n889));
  INV_X1    g464(.A(G2067), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n872), .A2(KEYINPUT95), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n880), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n863), .A2(new_n870), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n841), .A2(G35), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT97), .Z(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G162), .B2(new_n841), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT29), .ZN(new_n898));
  AOI211_X1 g473(.A(new_n844), .B(new_n894), .C1(G2090), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(G115), .A2(G2104), .ZN(new_n900));
  INV_X1    g475(.A(G127), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n476), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G2105), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(KEYINPUT91), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(KEYINPUT91), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g481(.A(G139), .B(new_n467), .C1(new_n480), .C2(new_n484), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(KEYINPUT25), .Z(new_n909));
  AOI21_X1  g484(.A(KEYINPUT90), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(KEYINPUT90), .A3(new_n909), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT92), .A4(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT92), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n904), .A2(new_n912), .A3(new_n905), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(G29), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(G29), .A2(G33), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT89), .Z(new_n919));
  AND2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n920), .A2(G2072), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(G2072), .A3(new_n919), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n843), .A2(new_n831), .B1(G2084), .B2(new_n852), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT94), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n898), .A2(G2090), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT98), .Z(new_n928));
  OR2_X1    g503(.A1(new_n924), .A2(new_n925), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n899), .A2(new_n926), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n820), .A2(new_n930), .ZN(G311));
  OR2_X1    g506(.A1(new_n820), .A2(new_n930), .ZN(G150));
  NAND2_X1  g507(.A1(new_n648), .A2(G559), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT99), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT38), .ZN(new_n935));
  OAI211_X1 g510(.A(G55), .B(G543), .C1(new_n552), .C2(new_n553), .ZN(new_n936));
  INV_X1    g511(.A(G93), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n561), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(G67), .B1(new_n549), .B2(new_n550), .ZN(new_n939));
  NAND2_X1  g514(.A1(G80), .A2(G543), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n565), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n580), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n578), .A3(new_n579), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n935), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT39), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT100), .ZN(new_n949));
  AOI21_X1  g524(.A(G860), .B1(new_n947), .B2(KEYINPUT39), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n943), .A2(G860), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT102), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n955), .ZN(G145));
  OAI21_X1  g531(.A(KEYINPUT103), .B1(new_n509), .B2(new_n511), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n505), .B1(new_n468), .B2(new_n469), .ZN(new_n958));
  INV_X1    g533(.A(new_n507), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n508), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT104), .B1(new_n499), .B2(new_n502), .ZN(new_n963));
  INV_X1    g538(.A(new_n498), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n468), .B2(new_n469), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n965), .B(new_n966), .C1(new_n500), .C2(new_n501), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n957), .A2(new_n962), .A3(new_n963), .A4(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n963), .A2(new_n967), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n888), .A2(new_n971), .A3(new_n957), .A4(new_n962), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n970), .A2(new_n840), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n840), .B1(new_n970), .B2(new_n972), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n916), .B(new_n913), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n976));
  INV_X1    g551(.A(G118), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(G2105), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n486), .B2(G130), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n480), .A2(new_n484), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(G142), .A3(new_n467), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n663), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n663), .A3(new_n981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n809), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n663), .B1(new_n979), .B2(new_n981), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(G130), .A3(G2105), .ZN(new_n988));
  INV_X1    g563(.A(new_n978), .ZN(new_n989));
  AND4_X1   g564(.A1(new_n663), .A2(new_n981), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n808), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n970), .A2(new_n972), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n839), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n970), .A2(new_n972), .A3(new_n840), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n975), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n975), .A2(new_n997), .ZN(new_n1001));
  INV_X1    g576(.A(new_n992), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n975), .A2(new_n992), .A3(new_n997), .A4(KEYINPUT105), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n496), .A2(G160), .ZN(new_n1006));
  INV_X1    g581(.A(G160), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n489), .A2(new_n495), .A3(new_n1007), .A4(new_n490), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n670), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n671), .A3(new_n1008), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT106), .B(G37), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n998), .A2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n1003), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g595(.A(KEYINPUT108), .B1(new_n942), .B2(G868), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n643), .A2(new_n647), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G299), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n592), .A2(new_n596), .A3(new_n643), .A4(new_n647), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT41), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(KEYINPUT41), .A3(new_n1024), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n946), .B(new_n658), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT42), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1035), .A3(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(new_n636), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G166), .A2(G290), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n797), .A2(KEYINPUT107), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT107), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n796), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(G305), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n796), .A2(new_n1041), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n796), .A2(new_n1041), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n783), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND4_X1   g621(.A1(new_n1038), .A2(new_n1039), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1038), .A2(new_n1039), .B1(new_n1046), .B2(new_n1043), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1037), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1034), .A2(new_n1036), .A3(new_n1049), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(G868), .A3(new_n1052), .ZN(new_n1053));
  MUX2_X1   g628(.A(KEYINPUT108), .B(new_n1021), .S(new_n1053), .Z(G295));
  MUX2_X1   g629(.A(KEYINPUT108), .B(new_n1021), .S(new_n1053), .Z(G331));
  INV_X1    g630(.A(new_n1025), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n518), .A2(G89), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n539), .B2(KEYINPUT75), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n541), .A2(new_n546), .A3(new_n543), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n546), .B1(new_n541), .B2(new_n543), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n556), .A2(new_n557), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(G301), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n548), .A2(G171), .A3(new_n558), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n944), .A2(new_n1062), .A3(new_n1063), .A4(new_n945), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1058), .A2(new_n1061), .A3(G301), .ZN(new_n1065));
  AOI21_X1  g640(.A(G171), .B1(new_n548), .B2(new_n558), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n942), .A2(new_n578), .A3(new_n579), .ZN(new_n1067));
  INV_X1    g642(.A(new_n941), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n518), .A2(G93), .B1(new_n520), .B2(G55), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n578), .A2(new_n579), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1065), .A2(new_n1066), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1056), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1064), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(KEYINPUT109), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n946), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1049), .B(new_n1072), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G37), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n946), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1076), .B1(new_n946), .B2(new_n1075), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1064), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1029), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1049), .B1(new_n1086), .B2(new_n1072), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT43), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1025), .B(new_n1073), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1079), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1050), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT43), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1080), .A3(new_n1092), .A4(new_n1015), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(KEYINPUT44), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1082), .A2(new_n1087), .A3(KEYINPUT43), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT110), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1091), .A2(new_n1015), .A3(new_n1080), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n1092), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1095), .B1(new_n1101), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g677(.A(new_n808), .B(new_n812), .Z(new_n1103));
  INV_X1    g678(.A(G1996), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n839), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n888), .B(new_n890), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n636), .B(G1986), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1384), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n962), .A2(new_n963), .A3(new_n967), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n961), .B1(new_n960), .B2(new_n508), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT45), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G160), .A2(G40), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1110), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n612), .A2(new_n741), .A3(new_n617), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G40), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n472), .A2(new_n478), .A3(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1111), .B(new_n1124), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n797), .A2(G1976), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1122), .A2(G8), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(G8), .A3(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT52), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n780), .A2(new_n565), .ZN(new_n1132));
  OAI21_X1  g707(.A(G1981), .B1(new_n1132), .B2(new_n622), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(G305), .B2(G1981), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT49), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT49), .B(new_n1133), .C1(G305), .C2(G1981), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(G8), .A3(new_n1125), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1131), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1125), .A2(G8), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1141), .A2(new_n1136), .A3(KEYINPUT113), .A4(new_n1138), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1130), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G303), .A2(G8), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT55), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT50), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n968), .B2(new_n1111), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n512), .A2(new_n1111), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1124), .B1(new_n1148), .B2(KEYINPUT50), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT112), .B(G2090), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1117), .B1(new_n1148), .B2(new_n1115), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1115), .A2(G1384), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n968), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1150), .A2(new_n1151), .B1(new_n740), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G8), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1145), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT55), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1144), .B(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1153), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n962), .A2(new_n963), .A3(new_n967), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(new_n957), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n960), .A2(new_n508), .ZN(new_n1164));
  AOI21_X1  g739(.A(G1384), .B1(new_n1164), .B2(new_n503), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1124), .B1(new_n1165), .B2(KEYINPUT45), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT111), .B(new_n740), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n968), .A2(new_n1146), .A3(new_n1111), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1117), .B1(new_n1148), .B2(KEYINPUT50), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(new_n1169), .A3(new_n1151), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT111), .B1(new_n1155), .B2(new_n740), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1160), .B(G8), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1143), .A2(new_n1158), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT114), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1124), .B1(G164), .B2(new_n1161), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1116), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1178), .B2(new_n859), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT45), .B1(new_n968), .B2(new_n1111), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1175), .B(new_n859), .C1(new_n1180), .C2(new_n1176), .ZN(new_n1181));
  INV_X1    g756(.A(G2084), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1168), .A2(new_n1169), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(G8), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(G286), .A2(G8), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT117), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT51), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1176), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT114), .B1(new_n1190), .B2(G1966), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(new_n1183), .A3(new_n1181), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1187), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1185), .A2(new_n1189), .A3(new_n1187), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1174), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n867), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT57), .ZN(new_n1199));
  XNOR2_X1  g774(.A(G299), .B(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT56), .B(G2072), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1152), .A2(new_n1154), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1198), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1205));
  INV_X1    g780(.A(G1348), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1125), .A2(G2067), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n648), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1200), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1204), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1207), .A2(new_n1208), .A3(KEYINPUT60), .A4(new_n1022), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT59), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1152), .A2(new_n1154), .A3(new_n1104), .ZN(new_n1217));
  XOR2_X1   g792(.A(KEYINPUT58), .B(G1341), .Z(new_n1218));
  NAND2_X1  g793(.A1(new_n1125), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n580), .A2(KEYINPUT116), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1216), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1221), .ZN(new_n1223));
  AOI211_X1 g798(.A(KEYINPUT59), .B(new_n1223), .C1(new_n1217), .C2(new_n1219), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1215), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1203), .A2(KEYINPUT61), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1198), .A2(new_n1227), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT60), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1209), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1207), .A2(KEYINPUT60), .A3(new_n1208), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(new_n648), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g809(.A(new_n1214), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g810(.A1(new_n1197), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1152), .A2(new_n1154), .A3(new_n855), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT53), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g814(.A1(new_n1238), .A2(G2078), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1240), .ZN(new_n1241));
  NOR3_X1   g816(.A1(new_n1180), .A2(new_n1241), .A3(new_n1176), .ZN(new_n1242));
  AOI21_X1  g817(.A(G1961), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1243));
  INV_X1    g818(.A(KEYINPUT119), .ZN(new_n1244));
  NOR3_X1   g819(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1205), .A2(new_n847), .ZN(new_n1246));
  NAND3_X1  g821(.A1(new_n1116), .A2(new_n1240), .A3(new_n1177), .ZN(new_n1247));
  AOI21_X1  g822(.A(KEYINPUT119), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1239), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g824(.A(KEYINPUT54), .B1(new_n1249), .B2(G171), .ZN(new_n1250));
  INV_X1    g825(.A(new_n478), .ZN(new_n1251));
  OR2_X1    g826(.A1(new_n1251), .A2(KEYINPUT120), .ZN(new_n1252));
  NOR3_X1   g827(.A1(new_n472), .A2(new_n1123), .A3(new_n1241), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1251), .A2(KEYINPUT120), .ZN(new_n1254));
  AND3_X1   g829(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g830(.A1(new_n1116), .A2(new_n1154), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g831(.A1(new_n1239), .A2(new_n1246), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g832(.A(KEYINPUT122), .ZN(new_n1258));
  AND3_X1   g833(.A1(new_n1257), .A2(new_n1258), .A3(G171), .ZN(new_n1259));
  AOI21_X1  g834(.A(new_n1258), .B1(new_n1257), .B2(G171), .ZN(new_n1260));
  NOR2_X1   g835(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g836(.A(KEYINPUT123), .B1(new_n1250), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g837(.A(new_n1260), .ZN(new_n1263));
  NAND3_X1  g838(.A1(new_n1257), .A2(new_n1258), .A3(G171), .ZN(new_n1264));
  NAND2_X1  g839(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g840(.A(KEYINPUT123), .ZN(new_n1266));
  OAI21_X1  g841(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1267));
  NAND3_X1  g842(.A1(new_n1246), .A2(new_n1247), .A3(KEYINPUT119), .ZN(new_n1268));
  AOI22_X1  g843(.A1(new_n1267), .A2(new_n1268), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1269));
  NAND2_X1  g844(.A1(new_n1269), .A2(G301), .ZN(new_n1270));
  NAND4_X1  g845(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT54), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g846(.A1(new_n1262), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g847(.A1(new_n1257), .A2(G171), .ZN(new_n1273));
  AOI21_X1  g848(.A(new_n1273), .B1(new_n1249), .B2(G171), .ZN(new_n1274));
  XNOR2_X1  g849(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n1275));
  OAI21_X1  g850(.A(KEYINPUT121), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g851(.A(KEYINPUT121), .ZN(new_n1277));
  INV_X1    g852(.A(new_n1275), .ZN(new_n1278));
  NOR2_X1   g853(.A1(new_n1269), .A2(G301), .ZN(new_n1279));
  OAI211_X1 g854(.A(new_n1277), .B(new_n1278), .C1(new_n1279), .C2(new_n1273), .ZN(new_n1280));
  NAND2_X1  g855(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  AND3_X1   g856(.A1(new_n1236), .A2(new_n1272), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g857(.A(KEYINPUT115), .ZN(new_n1283));
  OAI21_X1  g858(.A(G8), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1284));
  NAND2_X1  g859(.A1(new_n1284), .A2(new_n1145), .ZN(new_n1285));
  NAND4_X1  g860(.A1(new_n1285), .A2(new_n1143), .A3(KEYINPUT63), .A4(new_n1173), .ZN(new_n1286));
  NAND3_X1  g861(.A1(new_n1192), .A2(G8), .A3(G168), .ZN(new_n1287));
  OAI21_X1  g862(.A(new_n1283), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g863(.A(new_n740), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1289));
  INV_X1    g864(.A(KEYINPUT111), .ZN(new_n1290));
  NAND2_X1  g865(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g866(.A1(new_n1291), .A2(new_n1170), .A3(new_n1167), .ZN(new_n1292));
  AOI21_X1  g867(.A(new_n1160), .B1(new_n1292), .B2(G8), .ZN(new_n1293));
  NAND2_X1  g868(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1294));
  INV_X1    g869(.A(new_n1130), .ZN(new_n1295));
  NAND2_X1  g870(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g871(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  AND2_X1   g872(.A1(new_n1173), .A2(KEYINPUT63), .ZN(new_n1298));
  INV_X1    g873(.A(new_n1287), .ZN(new_n1299));
  NAND4_X1  g874(.A1(new_n1297), .A2(KEYINPUT115), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  INV_X1    g875(.A(KEYINPUT63), .ZN(new_n1301));
  NAND3_X1  g876(.A1(new_n1143), .A2(new_n1158), .A3(new_n1173), .ZN(new_n1302));
  OAI21_X1  g877(.A(new_n1301), .B1(new_n1302), .B2(new_n1287), .ZN(new_n1303));
  NAND3_X1  g878(.A1(new_n1288), .A2(new_n1300), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g879(.A(new_n1193), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1305));
  NAND2_X1  g880(.A1(new_n1305), .A2(KEYINPUT51), .ZN(new_n1306));
  AOI21_X1  g881(.A(new_n1193), .B1(new_n1192), .B2(G8), .ZN(new_n1307));
  OAI21_X1  g882(.A(new_n1196), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g883(.A(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g884(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g885(.A1(new_n1195), .A2(KEYINPUT62), .A3(new_n1196), .ZN(new_n1311));
  NOR3_X1   g886(.A1(new_n1302), .A2(G301), .A3(new_n1269), .ZN(new_n1312));
  NAND3_X1  g887(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  NOR2_X1   g888(.A1(new_n1296), .A2(new_n1173), .ZN(new_n1314));
  NAND3_X1  g889(.A1(new_n1294), .A2(new_n741), .A3(new_n618), .ZN(new_n1315));
  OAI21_X1  g890(.A(new_n1315), .B1(G1981), .B2(G305), .ZN(new_n1316));
  AOI21_X1  g891(.A(new_n1314), .B1(new_n1316), .B2(new_n1141), .ZN(new_n1317));
  NAND3_X1  g892(.A1(new_n1304), .A2(new_n1313), .A3(new_n1317), .ZN(new_n1318));
  OAI21_X1  g893(.A(new_n1119), .B1(new_n1282), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g894(.A1(new_n1118), .A2(new_n1104), .ZN(new_n1320));
  INV_X1    g895(.A(KEYINPUT46), .ZN(new_n1321));
  NOR2_X1   g896(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  XOR2_X1   g897(.A(new_n1322), .B(KEYINPUT124), .Z(new_n1323));
  NAND2_X1  g898(.A1(new_n1106), .A2(new_n840), .ZN(new_n1324));
  AOI22_X1  g899(.A1(new_n1320), .A2(new_n1321), .B1(new_n1118), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g900(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  XNOR2_X1  g901(.A(new_n1326), .B(KEYINPUT47), .ZN(new_n1327));
  INV_X1    g902(.A(new_n1118), .ZN(new_n1328));
  OR3_X1    g903(.A1(new_n1328), .A2(G1986), .A3(G290), .ZN(new_n1329));
  INV_X1    g904(.A(KEYINPUT48), .ZN(new_n1330));
  OR2_X1    g905(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g906(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1332));
  OAI211_X1 g907(.A(new_n1331), .B(new_n1332), .C1(new_n1328), .C2(new_n1108), .ZN(new_n1333));
  NAND2_X1  g908(.A1(new_n809), .A2(new_n812), .ZN(new_n1334));
  OAI22_X1  g909(.A1(new_n1107), .A2(new_n1334), .B1(G2067), .B2(new_n888), .ZN(new_n1335));
  NAND2_X1  g910(.A1(new_n1335), .A2(new_n1118), .ZN(new_n1336));
  AND3_X1   g911(.A1(new_n1327), .A2(new_n1333), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g912(.A1(new_n1319), .A2(new_n1337), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g913(.A(KEYINPUT127), .ZN(new_n1340));
  INV_X1    g914(.A(KEYINPUT126), .ZN(new_n1341));
  NAND2_X1  g915(.A1(G319), .A2(new_n729), .ZN(new_n1342));
  AOI21_X1  g916(.A(new_n1342), .B1(new_n706), .B2(new_n710), .ZN(new_n1343));
  NAND2_X1  g917(.A1(new_n1343), .A2(new_n778), .ZN(new_n1344));
  NAND2_X1  g918(.A1(new_n1344), .A2(KEYINPUT125), .ZN(new_n1345));
  INV_X1    g919(.A(KEYINPUT125), .ZN(new_n1346));
  NAND3_X1  g920(.A1(new_n1343), .A2(new_n778), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g921(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  AND4_X1   g922(.A1(new_n1341), .A2(new_n1094), .A3(new_n1019), .A4(new_n1348), .ZN(new_n1349));
  AOI22_X1  g923(.A1(new_n1014), .A2(new_n1018), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1350));
  AOI21_X1  g924(.A(new_n1341), .B1(new_n1350), .B2(new_n1094), .ZN(new_n1351));
  OAI21_X1  g925(.A(new_n1340), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g926(.A1(new_n1019), .A2(new_n1348), .ZN(new_n1353));
  AND2_X1   g927(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1354));
  OAI21_X1  g928(.A(KEYINPUT126), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g929(.A1(new_n1350), .A2(new_n1341), .A3(new_n1094), .ZN(new_n1356));
  NAND3_X1  g930(.A1(new_n1355), .A2(KEYINPUT127), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g931(.A1(new_n1352), .A2(new_n1357), .ZN(G308));
  NAND2_X1  g932(.A1(new_n1355), .A2(new_n1356), .ZN(G225));
endmodule


