//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT65), .B(G77), .Z(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT66), .B(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(G50), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n209), .A3(new_n230), .ZN(new_n231));
  NOR4_X1   g0031(.A1(new_n215), .A2(new_n227), .A3(new_n228), .A4(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G222), .A2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G223), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n257), .B(new_n258), .C1(new_n216), .C2(new_n253), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n250), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n260), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT68), .B(G226), .Z(new_n267));
  OAI211_X1 g0067(.A(new_n259), .B(new_n263), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI211_X1 g0070(.A(KEYINPUT71), .B(new_n270), .C1(G200), .C2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n230), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(new_n208), .B2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n279), .B2(new_n274), .ZN(new_n280));
  OAI21_X1  g0080(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n209), .A2(G33), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n281), .B1(new_n282), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n280), .B1(new_n289), .B2(new_n277), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(KEYINPUT9), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n271), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n268), .A2(G179), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT70), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n290), .B1(new_n297), .B2(new_n268), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G238), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n263), .B1(new_n266), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(G1698), .B1(new_n251), .B2(new_n252), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G226), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT72), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G33), .A3(G97), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n304), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n302), .B1(new_n311), .B2(new_n258), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n312), .A2(new_n313), .ZN(new_n316));
  OAI21_X1  g0116(.A(G169), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT14), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n312), .B(new_n313), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(G169), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n316), .A2(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(KEYINPUT73), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(new_n314), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n318), .B(new_n321), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n288), .A2(new_n327), .B1(new_n209), .B2(G68), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(KEYINPUT74), .B1(new_n274), .B2(new_n284), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n277), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT12), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n273), .A2(KEYINPUT75), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n333), .B2(KEYINPUT75), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n272), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n273), .A2(new_n277), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n334), .B1(new_n208), .B2(G20), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n335), .A2(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n322), .A2(G190), .A3(new_n323), .A4(new_n314), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(G200), .B2(new_n319), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n326), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n277), .ZN(new_n346));
  INV_X1    g0146(.A(new_n285), .ZN(new_n347));
  INV_X1    g0147(.A(G87), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT15), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT15), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G87), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n288), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n347), .A2(new_n283), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n216), .A2(G20), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n346), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n279), .A2(new_n327), .B1(new_n216), .B2(new_n272), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n253), .A2(G232), .A3(new_n255), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n205), .C2(new_n253), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n258), .ZN(new_n363));
  INV_X1    g0163(.A(new_n266), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n262), .B1(new_n364), .B2(new_n217), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n359), .B1(new_n367), .B2(G190), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n367), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n358), .B1(new_n366), .B2(new_n297), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n325), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n300), .A2(new_n345), .A3(new_n370), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n251), .A2(new_n209), .A3(new_n252), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT7), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n251), .A2(new_n377), .A3(new_n209), .A4(new_n252), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(G68), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n376), .A2(KEYINPUT76), .A3(G68), .A4(new_n378), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G58), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n334), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n201), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT77), .B(G20), .C1(new_n385), .C2(new_n201), .ZN(new_n389));
  INV_X1    g0189(.A(G159), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n284), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(new_n379), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n393), .A2(new_n396), .A3(new_n277), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n285), .B(KEYINPUT69), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n278), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n272), .B2(new_n398), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n399), .B(KEYINPUT78), .C1(new_n272), .C2(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n263), .B1(new_n266), .B2(new_n234), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n255), .A2(G226), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G223), .B2(G1698), .ZN(new_n408));
  AND2_X1   g0208(.A1(KEYINPUT3), .A2(G33), .ZN(new_n409));
  NOR2_X1   g0209(.A1(KEYINPUT3), .A2(G33), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n408), .A2(new_n411), .B1(new_n250), .B2(new_n348), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n412), .B2(new_n258), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G179), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n297), .B2(new_n413), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT18), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n269), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G200), .B2(new_n413), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n397), .A2(new_n404), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT79), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n397), .A2(new_n404), .A3(KEYINPUT79), .A4(new_n419), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n422), .A2(KEYINPUT80), .A3(KEYINPUT17), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n397), .A2(new_n404), .A3(new_n429), .A4(new_n419), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT81), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n417), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n374), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  NOR2_X1   g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n438), .A2(new_n265), .A3(G274), .A4(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n436), .B2(new_n437), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n265), .ZN(new_n443));
  INV_X1    g0243(.A(G270), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n411), .A2(G303), .ZN(new_n446));
  OAI211_X1 g0246(.A(G264), .B(G1698), .C1(new_n409), .C2(new_n410), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(new_n255), .C1(new_n409), .C2(new_n410), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n265), .B1(new_n449), .B2(KEYINPUT89), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT89), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n446), .A2(new_n451), .A3(new_n447), .A4(new_n448), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n445), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(KEYINPUT84), .A2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT84), .A2(G116), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(G20), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n458), .A3(new_n277), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT20), .A4(new_n277), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n208), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n272), .A2(new_n464), .A3(new_n230), .A4(new_n276), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n454), .A2(new_n455), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n466), .A2(G116), .B1(new_n273), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n453), .A2(G179), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT90), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT90), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n453), .A2(new_n473), .A3(G179), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n449), .A2(KEYINPUT89), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n258), .A3(new_n452), .ZN(new_n476));
  INV_X1    g0276(.A(new_n445), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n297), .B1(new_n463), .B2(new_n469), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(KEYINPUT21), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n472), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n481), .A2(KEYINPUT91), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(KEYINPUT91), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n479), .ZN(new_n484));
  XOR2_X1   g0284(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n470), .B1(new_n478), .B2(G200), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n269), .B2(new_n478), .ZN(new_n488));
  AND4_X1   g0288(.A1(new_n482), .A2(new_n483), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n376), .A2(G107), .A3(new_n378), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n283), .A2(G77), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT82), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT6), .B1(new_n206), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n490), .B(new_n492), .C1(new_n209), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n277), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n272), .A2(G97), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n466), .B2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G250), .A2(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n255), .A2(G244), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n253), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n457), .ZN(new_n507));
  OAI211_X1 g0307(.A(G244), .B(new_n255), .C1(new_n409), .C2(new_n410), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n508), .A2(new_n504), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n258), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n442), .A2(G257), .A3(new_n265), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n441), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n297), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n501), .B(new_n513), .C1(G179), .C2(new_n512), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(G200), .ZN(new_n515));
  INV_X1    g0315(.A(new_n500), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n497), .B2(new_n277), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n517), .C1(new_n269), .C2(new_n512), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n253), .A2(G244), .A3(G1698), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n253), .A2(G238), .A3(new_n255), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n467), .A2(G33), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n258), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n208), .A2(G45), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G250), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n258), .A2(new_n527), .B1(new_n261), .B2(new_n526), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n325), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n524), .B2(new_n258), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(G169), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n352), .A2(new_n272), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT85), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT85), .B1(new_n349), .B2(new_n351), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n535), .A2(new_n465), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n348), .A2(new_n204), .A3(new_n205), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n307), .B2(new_n309), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(G20), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n209), .B(G68), .C1(new_n409), .C2(new_n410), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n288), .B2(new_n204), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n534), .B(new_n538), .C1(new_n546), .C2(new_n346), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT86), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n346), .B1(new_n542), .B2(new_n545), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n533), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n538), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n532), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n531), .A2(G190), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n369), .B2(new_n531), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n466), .A2(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n553), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI211_X1 g0360(.A(G179), .B(new_n528), .C1(new_n524), .C2(new_n258), .ZN(new_n561));
  INV_X1    g0361(.A(new_n531), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n297), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n551), .B1(new_n550), .B2(new_n538), .ZN(new_n564));
  NOR4_X1   g0364(.A1(new_n549), .A2(KEYINPUT86), .A3(new_n537), .A4(new_n533), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(G200), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(new_n550), .A3(new_n556), .A4(new_n554), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT87), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n520), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT88), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n209), .B(G87), .C1(new_n409), .C2(new_n410), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n253), .A2(new_n575), .A3(new_n209), .A4(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n205), .A3(G20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n250), .B1(new_n454), .B2(new_n455), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(new_n209), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n577), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n578), .B1(new_n577), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n277), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT25), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n272), .B2(G107), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n272), .A2(new_n589), .A3(G107), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n591), .A2(new_n592), .B1(new_n205), .B2(new_n465), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n442), .A2(new_n258), .A3(new_n261), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n442), .A2(G264), .A3(new_n265), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT95), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n442), .A2(KEYINPUT95), .A3(G264), .A4(new_n265), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G250), .B(new_n255), .C1(new_n409), .C2(new_n410), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT93), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n253), .A2(KEYINPUT93), .A3(G250), .A4(new_n255), .ZN(new_n605));
  XNOR2_X1  g0405(.A(KEYINPUT94), .B(G294), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G33), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n604), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n258), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n441), .A2(new_n597), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n609), .B2(new_n258), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n611), .A2(new_n325), .B1(new_n613), .B2(new_n297), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n595), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g0415(.A(G190), .B(new_n612), .C1(new_n258), .C2(new_n609), .ZN(new_n616));
  AOI21_X1  g0416(.A(G200), .B1(new_n601), .B2(new_n610), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n588), .B(new_n594), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n559), .B1(new_n553), .B2(new_n558), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n566), .A2(KEYINPUT87), .A3(new_n568), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n519), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(KEYINPUT88), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n435), .A2(new_n489), .A3(new_n572), .A4(new_n623), .ZN(G372));
  AND2_X1   g0424(.A1(new_n480), .A2(new_n474), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n625), .A2(new_n615), .A3(new_n472), .A4(new_n486), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n514), .A2(new_n618), .A3(new_n518), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n553), .A2(new_n558), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n505), .A2(new_n253), .B1(G33), .B2(G283), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n508), .A2(new_n504), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n265), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n511), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(G169), .B1(new_n634), .B2(new_n441), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n632), .A2(G179), .A3(new_n633), .A4(new_n596), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(new_n517), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n566), .A2(new_n637), .A3(new_n638), .A4(new_n568), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n566), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n514), .B1(new_n620), .B2(new_n621), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n629), .B(new_n640), .C1(new_n641), .C2(new_n638), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n435), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n417), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n431), .B1(new_n426), .B2(new_n427), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n373), .B1(new_n344), .B2(new_n343), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n342), .B2(new_n326), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n643), .A2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(G213), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n470), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n489), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(KEYINPUT96), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(KEYINPUT96), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n656), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n588), .B2(new_n594), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n619), .A2(new_n667), .B1(new_n615), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n483), .A2(new_n486), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n656), .B1(new_n670), .B2(new_n482), .ZN(new_n671));
  INV_X1    g0471(.A(new_n619), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n595), .A2(new_n614), .A3(new_n666), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT97), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n212), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n539), .A2(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n229), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n670), .A2(new_n482), .A3(new_n615), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n628), .A3(new_n627), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n641), .A2(new_n638), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n628), .A2(new_n637), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n553), .B1(new_n689), .B2(KEYINPUT26), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n685), .B1(new_n691), .B2(new_n666), .ZN(new_n692));
  INV_X1    g0492(.A(G330), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n623), .A2(new_n489), .A3(new_n572), .A4(new_n666), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n478), .A2(new_n325), .ZN(new_n695));
  INV_X1    g0495(.A(new_n611), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n634), .A2(new_n531), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n696), .A4(new_n697), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n531), .A2(G179), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n478), .A2(new_n702), .A3(new_n611), .A4(new_n512), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n656), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT31), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n693), .B1(new_n694), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n642), .A2(new_n666), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n692), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n684), .B1(new_n710), .B2(G1), .ZN(G364));
  OR2_X1    g0511(.A1(new_n660), .A2(G330), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(KEYINPUT98), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(KEYINPUT98), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n209), .A2(G13), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT99), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G45), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G1), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n679), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n713), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n665), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n660), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n212), .A2(new_n253), .ZN(new_n727));
  INV_X1    g0527(.A(G355), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n727), .A2(new_n728), .B1(G116), .B2(new_n212), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n678), .A2(new_n253), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n229), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n439), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n244), .A2(new_n439), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n230), .B1(G20), .B2(new_n297), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n719), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n209), .A2(new_n269), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n325), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n209), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n325), .A3(G200), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G58), .A2(new_n742), .B1(new_n745), .B2(new_n216), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n744), .A2(G179), .A3(new_n369), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n205), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT102), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n741), .A2(new_n369), .A3(G179), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n411), .B1(new_n751), .B2(G87), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n752), .A2(new_n750), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n325), .A2(new_n369), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT100), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(KEYINPUT100), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n755), .A2(new_n743), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT103), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(KEYINPUT103), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G50), .A2(new_n761), .B1(new_n767), .B2(G68), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n743), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n770), .A2(new_n771), .A3(new_n390), .ZN(new_n772));
  INV_X1    g0572(.A(new_n771), .ZN(new_n773));
  INV_X1    g0573(.A(new_n770), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(G159), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n209), .B1(new_n769), .B2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n772), .B(new_n775), .C1(G97), .C2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n753), .A2(new_n754), .A3(new_n768), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n745), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n411), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n747), .A2(G283), .B1(G329), .B2(new_n774), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  INV_X1    g0584(.A(new_n751), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n782), .B(new_n786), .C1(new_n606), .C2(new_n777), .ZN(new_n787));
  INV_X1    g0587(.A(G326), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n760), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n742), .A2(G322), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT33), .B(G317), .Z(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n766), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT104), .Z(new_n793));
  OAI21_X1  g0593(.A(new_n779), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT105), .ZN(new_n795));
  INV_X1    g0595(.A(new_n736), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n794), .B2(KEYINPUT105), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n739), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n720), .A2(new_n721), .B1(new_n726), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  INV_X1    g0600(.A(new_n719), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n736), .A2(new_n722), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n327), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT106), .B(G283), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n760), .A2(new_n784), .B1(new_n766), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n742), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n806), .A2(new_n807), .B1(new_n780), .B2(new_n468), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n785), .A2(new_n205), .B1(new_n748), .B2(new_n348), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n411), .B1(new_n776), .B2(new_n204), .C1(new_n781), .C2(new_n770), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n805), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n748), .A2(new_n334), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n411), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n751), .A2(G50), .B1(G132), .B2(new_n774), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n384), .C2(new_n776), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G143), .A2(new_n742), .B1(new_n745), .B2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n766), .B2(new_n282), .C1(new_n817), .C2(new_n760), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n815), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n811), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n373), .A2(new_n656), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n370), .B1(new_n358), .B2(new_n666), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n373), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n803), .B1(new_n796), .B2(new_n822), .C1(new_n825), .C2(new_n723), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n708), .B(new_n825), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n707), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n719), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(new_n496), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT35), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(KEYINPUT35), .ZN(new_n836));
  INV_X1    g0636(.A(G116), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n230), .A2(new_n209), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT36), .Z(new_n840));
  OAI211_X1 g0640(.A(new_n732), .B(new_n216), .C1(new_n384), .C2(new_n334), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n274), .A2(G68), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n208), .B(G13), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n326), .A2(new_n342), .A3(new_n666), .ZN(new_n845));
  INV_X1    g0645(.A(new_n405), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n416), .B1(new_n846), .B2(new_n654), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n422), .A3(new_n423), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n393), .A2(new_n277), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n383), .B2(new_n392), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n399), .B1(new_n272), .B2(new_n398), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n654), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n415), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n422), .A3(new_n423), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n853), .ZN(new_n858));
  OAI211_X1 g0658(.A(KEYINPUT38), .B(new_n857), .C1(new_n433), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT107), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n858), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n645), .B2(new_n417), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n863), .A2(KEYINPUT107), .A3(KEYINPUT38), .A4(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n857), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n861), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n857), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n846), .A2(new_n654), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n645), .B2(new_n417), .ZN(new_n872));
  INV_X1    g0672(.A(new_n420), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n847), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n849), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n870), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n845), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n666), .B1(new_n332), .B2(new_n341), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n326), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n881), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n345), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n642), .A2(new_n666), .A3(new_n825), .ZN(new_n885));
  INV_X1    g0685(.A(new_n823), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n868), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n644), .A2(new_n853), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT108), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n868), .B2(new_n887), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n880), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n435), .B1(new_n692), .B2(new_n709), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n649), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n896), .B(new_n898), .Z(new_n899));
  INV_X1    g0699(.A(new_n825), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n694), .B2(new_n706), .ZN(new_n901));
  INV_X1    g0701(.A(new_n884), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n868), .A2(new_n904), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n900), .B(new_n884), .C1(new_n694), .C2(new_n706), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n870), .B2(new_n876), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n434), .B(new_n374), .C1(new_n694), .C2(new_n706), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n693), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n208), .B2(new_n716), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n899), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n844), .B1(new_n914), .B2(new_n915), .ZN(G367));
  INV_X1    g0716(.A(new_n669), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n637), .A2(new_n656), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT112), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n520), .B1(new_n517), .B2(new_n666), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n675), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n671), .A2(new_n672), .A3(new_n921), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n926), .A2(KEYINPUT42), .B1(new_n637), .B2(new_n666), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n557), .A2(new_n656), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n628), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT109), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n553), .A2(new_n557), .A3(new_n656), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n925), .A2(new_n927), .B1(KEYINPUT43), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT113), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n933), .A2(KEYINPUT110), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(KEYINPUT110), .ZN(new_n938));
  XNOR2_X1  g0738(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n935), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n936), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n923), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n923), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n679), .B(KEYINPUT41), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n676), .A2(new_n921), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT45), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n676), .A2(new_n921), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n917), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n952), .A3(new_n669), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n673), .B1(new_n668), .B2(new_n671), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n665), .B(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n710), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n948), .B1(new_n958), .B2(new_n710), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n947), .B1(new_n959), .B2(new_n718), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n933), .A2(new_n724), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n738), .B1(new_n678), .B2(new_n352), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n731), .B2(new_n240), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n719), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n253), .B(new_n965), .C1(G107), .C2(new_n777), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n748), .A2(new_n204), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G303), .B2(new_n742), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n774), .A2(G317), .ZN(new_n969));
  INV_X1    g0769(.A(new_n804), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n745), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n966), .A2(new_n968), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G311), .A2(new_n761), .B1(new_n767), .B2(new_n606), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT46), .B1(new_n751), .B2(new_n467), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT114), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G58), .A2(new_n751), .B1(new_n747), .B2(new_n216), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n742), .A2(G150), .B1(G137), .B2(new_n774), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n777), .A2(G68), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n411), .B1(new_n745), .B2(G50), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G143), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n760), .A2(new_n982), .B1(new_n766), .B2(new_n390), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n972), .A2(new_n976), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n964), .B1(new_n985), .B2(new_n736), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n961), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n960), .A2(new_n987), .ZN(G387));
  OR2_X1    g0788(.A1(new_n668), .A2(new_n725), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n727), .A2(new_n681), .B1(G107), .B2(new_n212), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n285), .A2(G50), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT115), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g0794(.A(G45), .B1(G68), .B2(G77), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n993), .A2(new_n681), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n731), .B1(new_n237), .B2(G45), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n719), .B1(new_n998), .B2(new_n738), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n806), .A2(new_n274), .B1(new_n780), .B2(new_n334), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n751), .A2(new_n216), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n282), .B2(new_n770), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n1000), .A2(new_n1002), .A3(new_n411), .A4(new_n967), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n535), .A2(new_n536), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n777), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G159), .A2(new_n761), .B1(new_n767), .B2(new_n398), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n253), .B1(new_n774), .B2(G326), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G317), .A2(new_n742), .B1(new_n745), .B2(G303), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT116), .B(G322), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n766), .B2(new_n781), .C1(new_n760), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n751), .A2(new_n606), .B1(new_n777), .B2(new_n970), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1008), .B1(new_n468), .B2(new_n748), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1007), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n999), .B1(new_n1020), .B2(new_n736), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n957), .A2(new_n718), .B1(new_n989), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n957), .A2(new_n710), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(KEYINPUT117), .A3(new_n679), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n710), .B2(new_n957), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT117), .B1(new_n1023), .B2(new_n679), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(G393));
  INV_X1    g0827(.A(new_n955), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n669), .B1(new_n950), .B2(new_n952), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1023), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n958), .A3(new_n679), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n730), .A2(new_n247), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n737), .C1(new_n204), .C2(new_n212), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n719), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n921), .A2(new_n725), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n760), .A2(new_n282), .B1(new_n390), .B2(new_n806), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n767), .A2(G50), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n780), .A2(new_n285), .B1(new_n770), .B2(new_n982), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G68), .B2(new_n751), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n776), .A2(new_n327), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n411), .B(new_n1041), .C1(G87), .C2(new_n747), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n780), .A2(new_n807), .B1(new_n770), .B2(new_n1010), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n411), .B1(new_n468), .B2(new_n776), .C1(new_n748), .C2(new_n205), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n751), .C2(new_n970), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n761), .A2(G317), .B1(G311), .B2(new_n742), .ZN(new_n1047));
  XOR2_X1   g0847(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1046), .B(new_n1049), .C1(new_n784), .C2(new_n766), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1034), .B(new_n1035), .C1(new_n736), .C2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n718), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1031), .A2(new_n1055), .ZN(G390));
  NAND2_X1  g0856(.A1(new_n435), .A2(new_n707), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n897), .A2(new_n649), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n901), .A2(G330), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n884), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n901), .A2(G330), .A3(new_n902), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n885), .A2(new_n886), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n824), .A2(new_n373), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n691), .A2(new_n666), .A3(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1066), .A2(new_n886), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1058), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT119), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1063), .A2(new_n902), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n845), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n845), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n887), .A2(KEYINPUT119), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n869), .A2(new_n1076), .A3(new_n878), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n845), .B1(new_n870), .B2(new_n876), .C1(new_n1067), .C2(new_n884), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n1061), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1061), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1070), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1061), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n1079), .A3(new_n1069), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n679), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n877), .B1(KEYINPUT39), .B2(new_n868), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n722), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G283), .A2(new_n761), .B1(new_n767), .B2(G107), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n812), .B1(G97), .B2(new_n745), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n742), .A2(G116), .B1(G294), .B2(new_n774), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n253), .B(new_n1041), .C1(new_n751), .C2(G87), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n785), .B2(new_n282), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n751), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n767), .A2(G137), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G132), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n806), .A2(new_n1099), .B1(new_n770), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G50), .B2(new_n747), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n253), .B1(new_n780), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G159), .B2(new_n777), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n761), .A2(G128), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1098), .A2(new_n1102), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n796), .B1(new_n1094), .B2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n801), .B(new_n1108), .C1(new_n287), .C2(new_n802), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1089), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT120), .B1(new_n1111), .B2(new_n718), .ZN(new_n1112));
  AND4_X1   g0912(.A1(KEYINPUT120), .A2(new_n1085), .A3(new_n718), .A4(new_n1079), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1087), .B(new_n1110), .C1(new_n1112), .C2(new_n1113), .ZN(G378));
  INV_X1    g0914(.A(new_n1058), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1086), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n894), .B1(new_n888), .B2(new_n890), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n879), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n294), .A2(new_n299), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n290), .A2(new_n654), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1122), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n300), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(new_n1123), .A3(new_n1119), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n909), .A2(G330), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n868), .A2(new_n904), .B1(new_n907), .B2(KEYINPUT40), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1130), .B1(new_n1133), .B2(new_n693), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1118), .A2(new_n895), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1131), .B1(new_n909), .B2(G330), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n693), .B(new_n1130), .C1(new_n905), .C2(new_n908), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1088), .A2(new_n845), .B1(new_n893), .B2(new_n894), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n893), .A2(new_n894), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1116), .A2(new_n1141), .A3(KEYINPUT57), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n679), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT125), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT57), .B1(new_n1116), .B2(new_n1141), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT125), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1147), .A3(new_n679), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT124), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1134), .A2(new_n1132), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n896), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1118), .A2(new_n895), .B1(new_n1134), .B2(new_n1132), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n718), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1130), .A2(new_n722), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n802), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n719), .B1(G50), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n761), .A2(G116), .B1(new_n1004), .B2(new_n745), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n204), .B2(new_n766), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n774), .A2(G283), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n748), .B2(new_n384), .C1(new_n205), .C2(new_n806), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1001), .A2(new_n264), .A3(new_n411), .A4(new_n979), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT58), .Z(new_n1164));
  OAI21_X1  g0964(.A(new_n274), .B1(new_n409), .B2(G41), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n806), .A2(new_n1166), .B1(new_n780), .B2(new_n817), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n785), .A2(new_n1103), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT121), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G150), .C2(new_n777), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n1100), .B2(new_n760), .C1(new_n1099), .C2(new_n766), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n747), .C2(G159), .ZN(new_n1174));
  INV_X1    g0974(.A(G124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n770), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1164), .B(new_n1165), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT123), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n796), .B1(new_n1177), .B2(KEYINPUT123), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1157), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1155), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1150), .B1(new_n1154), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n718), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1181), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1184), .A2(KEYINPUT124), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1149), .A2(new_n1188), .ZN(G375));
  NAND2_X1  g0989(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n884), .A2(new_n722), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n719), .B1(G68), .B2(new_n1156), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT126), .Z(new_n1193));
  OAI221_X1 g0993(.A(new_n253), .B1(new_n776), .B2(new_n274), .C1(new_n748), .C2(new_n384), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n806), .A2(new_n817), .B1(new_n780), .B2(new_n282), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n785), .A2(new_n390), .B1(new_n770), .B2(new_n1166), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n760), .A2(new_n1099), .B1(new_n766), .B2(new_n1103), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1005), .B1(new_n766), .B2(new_n468), .C1(new_n807), .C2(new_n760), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G283), .A2(new_n742), .B1(new_n747), .B2(G77), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n253), .B1(new_n751), .B2(G97), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n745), .A2(G107), .B1(G303), .B2(new_n774), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1197), .A2(new_n1198), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1193), .B1(new_n736), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1190), .A2(new_n718), .B1(new_n1191), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n948), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1070), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1190), .A2(new_n1115), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  INV_X1    g1011(.A(G384), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1213), .A2(G387), .A3(G381), .A4(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(G407));
  AOI21_X1  g1017(.A(new_n1145), .B1(new_n1143), .B2(KEYINPUT125), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1187), .B1(new_n1218), .B2(new_n1148), .ZN(new_n1219));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1221), .ZN(G409));
  NAND3_X1  g1022(.A1(new_n1070), .A2(new_n1209), .A3(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n679), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1209), .B1(new_n1070), .B2(KEYINPUT60), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1206), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(new_n1212), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1212), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n655), .A2(G213), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT127), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1115), .A2(new_n1086), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n1207), .ZN(new_n1235));
  AND4_X1   g1035(.A1(new_n1233), .A2(new_n1116), .A3(new_n1141), .A4(new_n1207), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1154), .A2(new_n1181), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G378), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1232), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1230), .B(new_n1240), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT62), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1142), .A2(new_n1147), .A3(new_n679), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1147), .B1(new_n1142), .B2(new_n679), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1145), .ZN(new_n1245));
  OAI21_X1  g1045(.A(G378), .B1(new_n1245), .B2(new_n1187), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1230), .A4(new_n1240), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1232), .A2(G2897), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1227), .A2(new_n1228), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1220), .B1(new_n1149), .B2(new_n1188), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1240), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1242), .A2(new_n1248), .A3(new_n1249), .A4(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n947), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1028), .A2(new_n1029), .A3(new_n1023), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n710), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1207), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1261), .B2(new_n1183), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n987), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1211), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G393), .B(new_n799), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n960), .A2(new_n987), .A3(G390), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1257), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1246), .A2(new_n1240), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1253), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1230), .A4(new_n1240), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1241), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1274), .A3(new_n1269), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1271), .A2(new_n1277), .ZN(G405));
  OAI21_X1  g1078(.A(new_n1230), .B1(new_n1216), .B2(new_n1254), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1246), .A2(new_n1221), .A3(new_n1229), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1279), .A2(new_n1269), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1269), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


