//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  AND2_X1   g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n213), .A2(G20), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n215), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  INV_X1    g0044(.A(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n242), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT69), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(new_n205), .B2(G20), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n206), .A2(KEYINPUT69), .A3(G1), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n243), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n255), .A2(new_n261), .B1(new_n243), .B2(new_n257), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n206), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n206), .A2(new_n266), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n263), .A2(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G58), .A2(G68), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n206), .B1(new_n269), .B2(new_n243), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n260), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G223), .A3(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G77), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(new_n274), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n214), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n205), .A2(new_n286), .B1(new_n214), .B2(new_n280), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n291), .A3(new_n285), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n214), .B2(new_n280), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n294), .A3(new_n205), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n273), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G179), .B2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n272), .B(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(new_n298), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n298), .A2(G200), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n303), .A2(new_n309), .A3(new_n305), .A4(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n206), .A2(G33), .A3(G77), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n245), .A2(G20), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n267), .C2(new_n243), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT72), .A3(new_n260), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT72), .B1(new_n314), .B2(new_n260), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT11), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT11), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n315), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n254), .A2(new_n245), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT12), .B1(new_n256), .B2(G68), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n256), .A2(KEYINPUT12), .A3(G68), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(new_n261), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n318), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n286), .A2(new_n205), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(G238), .A3(new_n281), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n295), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G226), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n275), .ZN(new_n334));
  INV_X1    g0134(.A(G232), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G1698), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n334), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n281), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n329), .B1(new_n332), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n340), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n282), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(new_n295), .A3(new_n328), .A4(new_n331), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(G169), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n332), .A2(new_n341), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n345), .B(G179), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n346), .B2(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n327), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n346), .A2(G200), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n345), .B(G190), .C1(new_n349), .C2(new_n350), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n326), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(KEYINPUT73), .A3(new_n357), .ZN(new_n361));
  INV_X1    g0161(.A(G244), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n330), .A2(new_n281), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n295), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n274), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n282), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n295), .B(new_n371), .C1(new_n362), .C2(new_n363), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n299), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n261), .B(G77), .C1(new_n253), .C2(new_n252), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G77), .B2(new_n256), .ZN(new_n376));
  INV_X1    g0176(.A(new_n260), .ZN(new_n377));
  INV_X1    g0177(.A(new_n263), .ZN(new_n378));
  NOR2_X1   g0178(.A1(G20), .A2(G33), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n378), .A2(new_n379), .B1(G20), .B2(G77), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(new_n264), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n377), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G179), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n365), .A2(new_n370), .A3(new_n386), .A4(new_n372), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n374), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n373), .A2(G200), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n365), .A2(new_n370), .A3(G190), .A4(new_n372), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n384), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n311), .A2(new_n360), .A3(new_n361), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n337), .A2(new_n338), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(new_n206), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n266), .ZN(new_n398));
  NAND2_X1  g0198(.A1(KEYINPUT3), .A2(G33), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n245), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n269), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n379), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n377), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n398), .A2(new_n206), .A3(new_n399), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n400), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT74), .B1(new_n415), .B2(G68), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT74), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n417), .B(new_n245), .C1(new_n414), .C2(new_n400), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n407), .A2(new_n410), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT75), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n402), .A2(new_n417), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(KEYINPUT74), .A3(G68), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT75), .A4(new_n420), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n411), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n261), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n254), .A2(new_n263), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(KEYINPUT76), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n430), .A2(new_n432), .B1(new_n257), .B2(new_n263), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n333), .A2(G1698), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(G223), .B2(G1698), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n435), .A2(new_n395), .B1(new_n266), .B2(new_n217), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n282), .B1(G232), .B2(new_n287), .ZN(new_n437));
  AOI21_X1  g0237(.A(G200), .B1(new_n437), .B2(new_n295), .ZN(new_n438));
  INV_X1    g0238(.A(G190), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n437), .A2(new_n295), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n426), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n433), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n422), .A2(new_n423), .A3(new_n420), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT75), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n424), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n450), .B2(new_n411), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n437), .A2(new_n295), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G169), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n386), .B2(new_n452), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT18), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n409), .A2(new_n410), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n260), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n449), .B2(new_n424), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n457), .B(new_n454), .C1(new_n460), .C2(new_n446), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n451), .A2(KEYINPUT17), .A3(new_n442), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n445), .A2(new_n456), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n394), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT5), .B1(new_n289), .B2(new_n291), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n205), .B(G45), .C1(new_n466), .C2(G41), .ZN(new_n467));
  OAI211_X1 g0267(.A(G270), .B(new_n281), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n469));
  INV_X1    g0269(.A(new_n467), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT68), .B(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(KEYINPUT5), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT81), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(G270), .A4(new_n281), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G303), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n398), .A2(new_n476), .A3(new_n399), .ZN(new_n477));
  MUX2_X1   g0277(.A(G257), .B(G264), .S(G1698), .Z(new_n478));
  OAI211_X1 g0278(.A(new_n282), .B(new_n477), .C1(new_n478), .C2(new_n395), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n470), .B(new_n294), .C1(KEYINPUT5), .C2(new_n471), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n257), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n205), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n256), .A2(new_n486), .A3(new_n259), .A4(new_n258), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(new_n484), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n258), .A2(new_n259), .B1(G20), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(new_n206), .C1(G33), .C2(new_n219), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT20), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n299), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n483), .A2(new_n496), .A3(KEYINPUT21), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n481), .B1(new_n469), .B2(new_n474), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n492), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n502), .B2(new_n488), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT82), .A3(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n483), .A2(new_n496), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT83), .B1(new_n500), .B2(new_n503), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n483), .A2(new_n386), .ZN(new_n512));
  INV_X1    g0312(.A(new_n495), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n483), .B2(G200), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n439), .B2(new_n483), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n506), .A2(new_n511), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n257), .A2(new_n219), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n487), .B2(new_n219), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT78), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n396), .B2(new_n401), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT6), .ZN(new_n523));
  AND2_X1   g0323(.A1(G97), .A2(G107), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n202), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n368), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT77), .B1(new_n267), .B2(new_n278), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT77), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n379), .A2(new_n529), .A3(G77), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n527), .A2(G20), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n521), .B1(new_n532), .B2(new_n260), .ZN(new_n533));
  AOI211_X1 g0333(.A(KEYINPUT78), .B(new_n377), .C1(new_n522), .C2(new_n531), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n520), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(new_n275), .C1(new_n337), .C2(new_n338), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n490), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n282), .ZN(new_n542));
  OAI211_X1 g0342(.A(G257), .B(new_n281), .C1(new_n465), .C2(new_n467), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(new_n480), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n542), .A2(new_n386), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(G169), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n535), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n368), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT25), .B1(new_n257), .B2(new_n368), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n368), .B2(new_n487), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G116), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(G20), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n206), .B2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n368), .A2(KEYINPUT23), .A3(G20), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n206), .B(G87), .C1(new_n337), .C2(new_n338), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n558), .A2(KEYINPUT22), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(KEYINPUT22), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT24), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(new_n557), .C1(new_n559), .C2(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n551), .B1(new_n565), .B2(new_n260), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n289), .A2(new_n291), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n466), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n282), .B1(new_n568), .B2(new_n470), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n218), .A2(new_n275), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n220), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n337), .C2(new_n338), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n569), .A2(G264), .B1(new_n282), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(KEYINPUT85), .A3(new_n439), .A4(new_n480), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT85), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n282), .ZN(new_n578));
  OAI211_X1 g0378(.A(G264), .B(new_n281), .C1(new_n465), .C2(new_n467), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n480), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G200), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(G190), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n576), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n566), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n528), .A2(new_n530), .ZN(new_n586));
  XNOR2_X1  g0386(.A(G97), .B(G107), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n523), .A2(new_n219), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n523), .B1(new_n368), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n589), .B2(new_n206), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n368), .B1(new_n414), .B2(new_n400), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n260), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n532), .A2(new_n521), .A3(new_n260), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n519), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n542), .A2(new_n439), .A3(new_n544), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n543), .A2(new_n480), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n282), .B2(new_n541), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n598), .B2(G200), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n548), .A2(new_n585), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n602), .A3(G169), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n386), .B2(new_n580), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n580), .B2(G169), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n377), .B1(new_n562), .B2(new_n564), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n551), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n206), .B1(new_n340), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G87), .B2(new_n203), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n206), .B(G68), .C1(new_n337), .C2(new_n338), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n608), .B1(new_n264), .B2(new_n219), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n260), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n381), .A2(new_n257), .ZN(new_n615));
  INV_X1    g0415(.A(new_n487), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G87), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n205), .A2(new_n293), .A3(G45), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n218), .B1(new_n285), .B2(G1), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n281), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(G244), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n623));
  OAI211_X1 g0423(.A(G238), .B(new_n275), .C1(new_n337), .C2(new_n338), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n552), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT79), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n281), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT79), .A4(new_n552), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n618), .B1(new_n629), .B2(G190), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(new_n626), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n282), .A3(new_n628), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n621), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G200), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n381), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n616), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n614), .A2(new_n615), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT80), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n614), .A2(KEYINPUT80), .A3(new_n615), .A4(new_n637), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n386), .B(new_n622), .C1(new_n627), .C2(new_n628), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n299), .B1(new_n632), .B2(new_n621), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n607), .A2(new_n635), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n517), .A2(new_n601), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n464), .A2(new_n646), .ZN(G372));
  AND2_X1   g0447(.A1(new_n456), .A2(new_n461), .ZN(new_n648));
  INV_X1    g0448(.A(new_n388), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n357), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n354), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n445), .A2(new_n462), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n653), .A2(new_n654), .B1(new_n308), .B2(new_n310), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n302), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n464), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT88), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n542), .A2(new_n386), .A3(new_n544), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n598), .B2(G169), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n595), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n535), .A2(new_n547), .A3(KEYINPUT88), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n632), .A2(G179), .A3(new_n621), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n299), .B2(new_n629), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n665), .A2(new_n638), .B1(new_n630), .B2(new_n634), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n662), .A2(new_n663), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n644), .A2(new_n635), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT26), .B1(new_n669), .B2(new_n548), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n665), .A2(new_n671), .A3(new_n638), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n665), .B2(new_n638), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n668), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT82), .B1(new_n504), .B2(KEYINPUT21), .ZN(new_n677));
  NOR4_X1   g0477(.A1(new_n500), .A2(new_n503), .A3(new_n498), .A4(new_n510), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n511), .B(new_n514), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n666), .A2(new_n548), .A3(new_n600), .A4(new_n585), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n680), .A2(new_n607), .B1(new_n681), .B2(KEYINPUT86), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n593), .A2(new_n594), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n599), .A2(new_n683), .A3(new_n520), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n595), .A2(new_n661), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT86), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(new_n585), .A4(new_n666), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n676), .B1(new_n682), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n657), .B1(new_n658), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT90), .ZN(G369));
  NAND3_X1  g0491(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n566), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n585), .A3(new_n607), .ZN(new_n701));
  INV_X1    g0501(.A(new_n607), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n697), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n698), .A2(new_n495), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n679), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n517), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n679), .A2(new_n698), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n701), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n702), .A2(new_n698), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0516(.A(new_n209), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n567), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n213), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n719), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  INV_X1    g0524(.A(G330), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n632), .A2(new_n575), .A3(new_n621), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n629), .A2(new_n728), .A3(new_n575), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n512), .A2(new_n727), .A3(new_n598), .A4(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n542), .A2(new_n544), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n483), .A2(new_n733), .A3(new_n386), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(KEYINPUT30), .A3(new_n729), .A4(new_n727), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n580), .A2(new_n386), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n483), .A3(new_n633), .A4(new_n733), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n697), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n646), .A2(new_n698), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n725), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n685), .A2(new_n667), .A3(new_n635), .A4(new_n644), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n675), .B(new_n745), .C1(new_n746), .C2(new_n667), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n681), .B1(new_n680), .B2(new_n607), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT29), .B(new_n698), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n506), .A2(new_n511), .A3(new_n514), .A4(new_n607), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n681), .A2(KEYINPUT86), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n688), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n668), .A2(new_n670), .A3(new_n675), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n697), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n749), .B1(new_n754), .B2(KEYINPUT29), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n744), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n724), .B1(new_n757), .B2(G1), .ZN(G364));
  AND2_X1   g0558(.A1(new_n206), .A2(G13), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n205), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n718), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n708), .B2(G330), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G330), .B2(new_n708), .ZN(new_n764));
  INV_X1    g0564(.A(new_n762), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n206), .B1(KEYINPUT96), .B2(new_n299), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n299), .A2(KEYINPUT96), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n259), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n206), .A2(new_n386), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n439), .A3(new_n581), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n274), .B1(new_n771), .B2(new_n278), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n581), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n243), .A2(new_n775), .B1(new_n777), .B2(new_n403), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n206), .A2(new_n386), .A3(new_n581), .A4(G190), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n772), .B(new_n778), .C1(G68), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n206), .B1(new_n781), .B2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n219), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n206), .A2(new_n581), .A3(G179), .A4(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n368), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n206), .A2(new_n439), .A3(new_n581), .A4(G179), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n783), .B(new_n786), .C1(G87), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n781), .A2(G20), .A3(new_n439), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT97), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  OR3_X1    g0593(.A1(new_n792), .A2(KEYINPUT32), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT32), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n780), .A2(new_n788), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n771), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n274), .B1(new_n797), .B2(G311), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  INV_X1    g0599(.A(new_n779), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n792), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G329), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G303), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n776), .A2(G322), .B1(G283), .B2(new_n784), .ZN(new_n809));
  INV_X1    g0609(.A(new_n782), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n774), .A2(G326), .B1(G294), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n803), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n769), .B1(new_n796), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G13), .A2(G33), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G20), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT95), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n768), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n717), .A2(new_n395), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT94), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G355), .B1(new_n484), .B2(new_n717), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n249), .A2(new_n285), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n717), .A2(new_n274), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n722), .B2(G45), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n765), .B(new_n813), .C1(new_n819), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n708), .B2(new_n817), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n764), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n385), .A2(new_n697), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n388), .A2(new_n391), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT101), .A4(new_n831), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n649), .A2(new_n697), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n698), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n754), .A2(new_n837), .B1(new_n689), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n762), .B1(new_n744), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n744), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n768), .A2(new_n814), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n762), .B1(new_n844), .B2(G77), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n395), .B1(new_n806), .B2(new_n368), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT99), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n785), .A2(new_n217), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n775), .A2(new_n476), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(G294), .C2(new_n776), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n800), .A2(new_n851), .B1(new_n771), .B2(new_n484), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n783), .B(new_n852), .C1(G311), .C2(new_n802), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n847), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n274), .B1(new_n792), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT100), .Z(new_n857));
  AOI22_X1  g0657(.A1(new_n797), .A2(G159), .B1(new_n779), .B2(G150), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n776), .A2(G143), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n775), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n785), .A2(new_n245), .B1(new_n403), .B2(new_n782), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n807), .B2(G50), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n854), .B1(new_n857), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n845), .B1(new_n868), .B2(new_n768), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n815), .B2(new_n837), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n842), .A2(new_n870), .ZN(G384));
  NAND2_X1  g0671(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n259), .A2(new_n206), .A3(new_n484), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n527), .B2(KEYINPUT35), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT102), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT36), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n213), .B(G77), .C1(new_n403), .C2(new_n245), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n205), .B(G13), .C1(new_n879), .C2(new_n244), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT103), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n839), .B1(new_n752), .B2(new_n753), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n388), .A2(new_n697), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n884), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT103), .B(new_n886), .C1(new_n689), .C2(new_n839), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n422), .A2(new_n423), .A3(new_n408), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n377), .B1(new_n889), .B2(new_n410), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n446), .B1(new_n450), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n443), .B1(new_n455), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n695), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n695), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n460), .A2(new_n446), .B1(new_n454), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n443), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n463), .A2(new_n893), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n326), .A2(new_n698), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n354), .A2(new_n357), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n354), .A2(new_n910), .A3(new_n357), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n353), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n357), .A2(new_n913), .A3(new_n351), .A4(new_n348), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n906), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(KEYINPUT105), .A3(new_n906), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n888), .A2(new_n905), .A3(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n648), .A2(new_n895), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n354), .A2(new_n697), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n899), .B2(new_n900), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT39), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n904), .A2(KEYINPUT108), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n899), .A2(new_n900), .A3(new_n931), .A4(KEYINPUT38), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT107), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT106), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n451), .B2(new_n442), .ZN(new_n936));
  NOR4_X1   g0736(.A1(new_n460), .A2(KEYINPUT106), .A3(new_n446), .A4(new_n441), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n426), .A2(new_n433), .B1(new_n455), .B2(new_n695), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n934), .B1(new_n939), .B2(new_n897), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n443), .A2(KEYINPUT106), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n896), .ZN(new_n942));
  OAI211_X1 g0742(.A(KEYINPUT107), .B(KEYINPUT37), .C1(new_n942), .C2(new_n937), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n898), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n895), .B1(new_n460), .B2(new_n446), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n463), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n928), .B1(new_n933), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n923), .B1(new_n925), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n464), .B(new_n749), .C1(new_n754), .C2(KEYINPUT29), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n657), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n950), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n837), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n912), .B2(new_n919), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n739), .A2(new_n740), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n601), .A2(new_n645), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n957), .A2(new_n680), .A3(new_n516), .A4(new_n698), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n958), .A3(new_n742), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT109), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(KEYINPUT40), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n955), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT109), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n929), .A2(new_n932), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n962), .B(new_n964), .C1(new_n965), .C2(new_n948), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT40), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n926), .A2(new_n927), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n963), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n464), .A2(new_n959), .ZN(new_n971));
  OAI21_X1  g0771(.A(G330), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n953), .A2(new_n973), .B1(new_n205), .B2(new_n759), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n953), .A2(new_n973), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n881), .B1(new_n974), .B2(new_n975), .ZN(G367));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n712), .A2(new_n713), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n686), .B1(new_n595), .B2(new_n698), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n685), .A2(new_n697), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n977), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n981), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n714), .B2(new_n983), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT111), .B1(new_n710), .B2(KEYINPUT112), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(KEYINPUT111), .A3(new_n989), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT112), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n710), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n711), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n712), .B1(new_n704), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(new_n709), .Z(new_n1000));
  AOI21_X1  g0800(.A(new_n756), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n718), .B(KEYINPUT41), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n760), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n981), .B(KEYINPUT110), .Z(new_n1004));
  AOI21_X1  g0804(.A(new_n685), .B1(new_n1004), .B2(new_n702), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(new_n697), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n712), .A2(new_n983), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT42), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n618), .A2(new_n697), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n675), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n666), .A2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n1009), .A2(KEYINPUT43), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1009), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1004), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n996), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1020), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1003), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n819), .B1(new_n209), .B2(new_n381), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n824), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n236), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n762), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n782), .A2(new_n245), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n274), .B1(new_n243), .B2(new_n771), .C1(new_n800), .C2(new_n793), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G143), .C2(new_n774), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n777), .A2(new_n265), .B1(new_n278), .B2(new_n785), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G58), .B2(new_n787), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT113), .B(G137), .Z(new_n1034));
  OAI211_X1 g0834(.A(new_n1031), .B(new_n1033), .C1(new_n792), .C2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT114), .Z(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT46), .B1(new_n787), .B2(G116), .ZN(new_n1037));
  INV_X1    g0837(.A(G294), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n395), .B1(new_n851), .B2(new_n771), .C1(new_n800), .C2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(G317), .C2(new_n802), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n774), .A2(G311), .B1(G107), .B2(new_n810), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n776), .A2(G303), .B1(G97), .B2(new_n784), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1036), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT47), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1028), .B1(new_n1046), .B2(new_n768), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n817), .B2(new_n1014), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT115), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1024), .A2(new_n1050), .ZN(G387));
  NOR2_X1   g0851(.A1(new_n233), .A2(new_n285), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n378), .A2(new_n243), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n720), .B(new_n285), .C1(new_n245), .C2(new_n278), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n824), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(KEYINPUT116), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(KEYINPUT116), .B2(new_n1056), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n821), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(G107), .B2(new_n209), .C1(new_n720), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n819), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n787), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n775), .A2(new_n793), .B1(new_n278), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n636), .B2(new_n810), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n802), .A2(G150), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n274), .B1(new_n245), .B2(new_n771), .C1(new_n800), .C2(new_n263), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n776), .A2(G50), .B1(G97), .B2(new_n784), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n802), .A2(G326), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n274), .B1(new_n784), .B2(G116), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1062), .A2(new_n1038), .B1(new_n851), .B2(new_n782), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n797), .A2(G303), .B1(new_n779), .B2(G311), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n776), .A2(G317), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n774), .A2(G322), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1070), .B(new_n1071), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1069), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n768), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1061), .A2(new_n762), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n705), .B2(new_n818), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n1000), .B2(new_n761), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1000), .A2(new_n757), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n718), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1000), .A2(new_n757), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  AOI22_X1  g0891(.A1(G311), .A2(new_n776), .B1(new_n774), .B2(G317), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  NOR2_X1   g0893(.A1(new_n782), .A2(new_n484), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1094), .B(new_n786), .C1(G283), .C2(new_n787), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n802), .A2(G322), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n395), .B1(new_n771), .B2(new_n1038), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G303), .B2(new_n779), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G150), .A2(new_n774), .B1(new_n776), .B2(G159), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT51), .Z(new_n1101));
  NOR2_X1   g0901(.A1(new_n782), .A2(new_n278), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1102), .B(new_n848), .C1(G68), .C2(new_n787), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n802), .A2(G143), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n274), .B1(new_n771), .B2(new_n263), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G50), .B2(new_n779), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n769), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n242), .A2(new_n1026), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n819), .B1(new_n219), .B2(new_n209), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n762), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1108), .B(new_n1111), .C1(new_n1021), .C2(new_n818), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n990), .B(new_n710), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n760), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1088), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n997), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n719), .B1(new_n1114), .B2(new_n1088), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(G390));
  INV_X1    g0920(.A(new_n920), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n885), .B2(new_n887), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n928), .B1(new_n933), .B2(new_n948), .C1(new_n1122), .C2(new_n925), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n959), .A2(G330), .A3(new_n837), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n747), .A2(new_n748), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n886), .B1(new_n1127), .B2(new_n839), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n925), .B1(new_n1128), .B2(new_n920), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n965), .B2(new_n948), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n925), .B1(new_n888), .B2(new_n920), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n949), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1126), .A2(new_n1124), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n743), .A2(new_n837), .A3(new_n920), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT117), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n949), .A2(new_n815), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n762), .B1(new_n844), .B2(new_n378), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n484), .A2(new_n777), .B1(new_n775), .B2(new_n851), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1102), .B(new_n1141), .C1(G68), .C2(new_n784), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n395), .B1(new_n219), .B2(new_n771), .C1(new_n800), .C2(new_n368), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G294), .B2(new_n802), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n217), .C2(new_n806), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT118), .Z(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n775), .A2(new_n1147), .B1(new_n243), .B2(new_n785), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n777), .A2(new_n855), .B1(new_n782), .B2(new_n793), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n802), .A2(G125), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n787), .A2(G150), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT53), .Z(new_n1153));
  OAI21_X1  g0953(.A(new_n274), .B1(new_n800), .B2(new_n1034), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n797), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .A4(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT119), .B1(new_n1146), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n769), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1146), .A2(KEYINPUT119), .A3(new_n1158), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1140), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1138), .A2(new_n761), .B1(new_n1139), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n743), .A2(new_n464), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n657), .A2(new_n951), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n920), .B1(new_n743), .B2(new_n837), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n888), .B1(new_n1166), .B2(new_n1126), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1128), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1135), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1165), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n718), .B1(new_n1138), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1163), .B1(new_n1172), .B2(new_n1174), .ZN(G378));
  OAI21_X1  g0975(.A(new_n762), .B1(new_n844), .B2(G50), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n273), .A2(new_n695), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n311), .B(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1178), .B(new_n1179), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n815), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n777), .A2(new_n368), .B1(new_n403), .B2(new_n785), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n395), .B(new_n471), .C1(new_n800), .C2(new_n219), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n636), .B2(new_n797), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1029), .B1(G77), .B2(new_n787), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n851), .C2(new_n792), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1183), .B(new_n1187), .C1(G116), .C2(new_n774), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n800), .A2(new_n855), .B1(new_n771), .B2(new_n860), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n774), .A2(G125), .B1(G150), .B2(new_n810), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1147), .B2(new_n777), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n787), .C2(new_n1156), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n802), .A2(G124), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n784), .C2(G159), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n243), .B1(G33), .B2(G41), .C1(new_n567), .C2(new_n274), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1189), .A2(new_n1199), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1176), .B(new_n1182), .C1(new_n768), .C2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n965), .A2(new_n948), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n964), .A2(KEYINPUT40), .A3(new_n961), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n969), .B(G330), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1180), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n966), .A2(G330), .A3(new_n969), .A4(new_n1181), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n950), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n950), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1204), .B1(new_n1214), .B2(new_n761), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n950), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n949), .A2(new_n925), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n923), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1208), .A2(new_n1209), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1174), .A2(new_n1165), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n718), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1134), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1171), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1165), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1214), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1215), .B1(new_n1222), .B2(new_n1228), .ZN(G375));
  INV_X1    g1029(.A(new_n1170), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1135), .A2(new_n1169), .B1(new_n885), .B2(new_n887), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n761), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n274), .B1(new_n779), .B2(G116), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n368), .B2(new_n771), .C1(new_n792), .C2(new_n476), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n806), .A2(new_n219), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n785), .A2(new_n278), .B1(new_n381), .B2(new_n782), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n851), .A2(new_n777), .B1(new_n775), .B2(new_n1038), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n395), .B1(new_n797), .B2(G150), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n800), .B2(new_n1155), .C1(new_n792), .C2(new_n1147), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n806), .A2(new_n793), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n777), .A2(new_n1034), .B1(new_n403), .B2(new_n785), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n775), .A2(new_n855), .B1(new_n782), .B2(new_n243), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n768), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n765), .B1(new_n843), .B2(new_n245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n920), .C2(new_n815), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1232), .A2(KEYINPUT121), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT121), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n760), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1002), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1167), .A2(new_n1165), .A3(new_n1170), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1173), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT122), .ZN(G381));
  XNOR2_X1  g1058(.A(G375), .B(KEYINPUT123), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1119), .A2(new_n1260), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(G387), .A2(G378), .A3(G381), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(G407));
  INV_X1    g1063(.A(G378), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1259), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1255), .B1(new_n1171), .B2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1167), .A2(new_n1165), .A3(KEYINPUT60), .A4(new_n1170), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n718), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n1253), .A3(G384), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1272), .B2(new_n1253), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1266), .ZN(new_n1280));
  INV_X1    g1080(.A(G2897), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1272), .A2(new_n1253), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1273), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1286), .B2(KEYINPUT124), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1277), .A3(new_n1273), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT125), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1279), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1289), .B2(new_n1279), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1215), .C1(new_n1222), .C2(new_n1228), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1215), .B1(new_n1002), .B2(new_n1220), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1264), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1266), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(new_n829), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1119), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1024), .A2(new_n1050), .A3(G390), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G390), .B1(new_n1024), .B2(new_n1050), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1049), .B(new_n1119), .C1(new_n1003), .C2(new_n1023), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1299), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1296), .A2(new_n1276), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1266), .B(new_n1286), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1298), .A2(new_n1307), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1286), .A2(KEYINPUT124), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1282), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1278), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1288), .A2(KEYINPUT125), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1317), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1279), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1314), .B1(new_n1322), .B2(new_n1296), .ZN(new_n1323));
  AND2_X1   g1123(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1311), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1308), .A2(new_n1325), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1323), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1313), .B1(new_n1329), .B2(new_n1307), .ZN(G405));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1331), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1300), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1305), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1333), .A2(new_n1334), .A3(KEYINPUT127), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(G375), .B(G378), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1286), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1336), .A2(new_n1286), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1332), .B(new_n1335), .C1(new_n1338), .C2(new_n1339), .ZN(new_n1340));
  OR2_X1    g1140(.A1(new_n1336), .A2(new_n1286), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1341), .A2(new_n1307), .A3(KEYINPUT127), .A4(new_n1337), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(G402));
endmodule


