

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XOR2_X1 U325 ( .A(n313), .B(KEYINPUT18), .Z(n293) );
  NOR2_X1 U326 ( .A1(n380), .A2(n379), .ZN(n381) );
  XNOR2_X1 U327 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n312) );
  XNOR2_X1 U328 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U329 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U330 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n343) );
  NOR2_X1 U331 ( .A1(n469), .A2(n468), .ZN(n486) );
  XNOR2_X1 U332 ( .A(n578), .B(n343), .ZN(n547) );
  XNOR2_X1 U333 ( .A(n324), .B(n323), .ZN(n530) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n449) );
  XOR2_X1 U335 ( .A(n461), .B(KEYINPUT28), .Z(n533) );
  XNOR2_X1 U336 ( .A(n491), .B(n490), .ZN(n501) );
  XNOR2_X1 U337 ( .A(n449), .B(KEYINPUT58), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(G99GAT), .B(G85GAT), .Z(n327) );
  XOR2_X1 U341 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n295) );
  XNOR2_X1 U342 ( .A(G190GAT), .B(KEYINPUT11), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U344 ( .A(n327), .B(n296), .Z(n300) );
  XOR2_X1 U345 ( .A(G29GAT), .B(G36GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n346) );
  XOR2_X1 U348 ( .A(G50GAT), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U349 ( .A(n346), .B(n404), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U351 ( .A(n301), .B(KEYINPUT9), .Z(n303) );
  XOR2_X1 U352 ( .A(G43GAT), .B(G134GAT), .Z(n320) );
  XNOR2_X1 U353 ( .A(n320), .B(G218GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U355 ( .A(G92GAT), .B(KEYINPUT65), .Z(n305) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U358 ( .A(G106GAT), .B(n306), .Z(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n541) );
  XOR2_X1 U360 ( .A(G71GAT), .B(KEYINPUT81), .Z(n310) );
  NAND2_X1 U361 ( .A1(G227GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U363 ( .A(KEYINPUT20), .B(n311), .ZN(n324) );
  XOR2_X1 U364 ( .A(G15GAT), .B(G127GAT), .Z(n362) );
  XOR2_X1 U365 ( .A(n362), .B(KEYINPUT82), .Z(n316) );
  XNOR2_X1 U366 ( .A(n312), .B(KEYINPUT19), .ZN(n313) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n293), .B(n314), .ZN(n401) );
  XNOR2_X1 U369 ( .A(n401), .B(G99GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U371 ( .A(G176GAT), .B(G120GAT), .Z(n328) );
  XOR2_X1 U372 ( .A(n317), .B(n328), .Z(n322) );
  XOR2_X1 U373 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n319) );
  XNOR2_X1 U374 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n439) );
  XNOR2_X1 U376 ( .A(n320), .B(n439), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U378 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n446) );
  XNOR2_X1 U379 ( .A(G204GAT), .B(G92GAT), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n325), .B(G64GAT), .ZN(n391) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n326), .B(KEYINPUT13), .ZN(n366) );
  XNOR2_X1 U383 ( .A(n391), .B(n366), .ZN(n342) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n330) );
  XOR2_X1 U385 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U387 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n332) );
  XNOR2_X1 U388 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n334) );
  AND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U391 ( .A(KEYINPUT69), .B(n337), .Z(n340) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n338), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U394 ( .A(n418), .B(KEYINPUT70), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n578) );
  XOR2_X1 U397 ( .A(G197GAT), .B(G22GAT), .Z(n345) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G141GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n359) );
  XOR2_X1 U400 ( .A(KEYINPUT68), .B(G1GAT), .Z(n363) );
  XOR2_X1 U401 ( .A(n363), .B(G43GAT), .Z(n348) );
  XNOR2_X1 U402 ( .A(G50GAT), .B(n346), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n350) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT67), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U409 ( .A(G113GAT), .B(G15GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n355), .B(KEYINPUT29), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n558) );
  NAND2_X1 U414 ( .A1(n547), .A2(n558), .ZN(n361) );
  XOR2_X1 U415 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n380) );
  XOR2_X1 U417 ( .A(G8GAT), .B(G211GAT), .Z(n395) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n409) );
  XOR2_X1 U419 ( .A(n395), .B(n409), .Z(n365) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U422 ( .A(n366), .B(KEYINPUT14), .Z(n368) );
  NAND2_X1 U423 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U425 ( .A(n370), .B(n369), .Z(n378) );
  XOR2_X1 U426 ( .A(KEYINPUT78), .B(G64GAT), .Z(n372) );
  XNOR2_X1 U427 ( .A(G183GAT), .B(G78GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U429 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n374) );
  XNOR2_X1 U430 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n581) );
  XOR2_X1 U434 ( .A(n581), .B(KEYINPUT115), .Z(n568) );
  NAND2_X1 U435 ( .A1(n568), .A2(n541), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n381), .B(KEYINPUT47), .ZN(n387) );
  XNOR2_X1 U437 ( .A(KEYINPUT36), .B(n541), .ZN(n584) );
  NOR2_X1 U438 ( .A1(n584), .A2(n581), .ZN(n382) );
  XNOR2_X1 U439 ( .A(KEYINPUT45), .B(n382), .ZN(n383) );
  NAND2_X1 U440 ( .A1(n383), .A2(n578), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT117), .ZN(n385) );
  INV_X1 U442 ( .A(n558), .ZN(n574) );
  NAND2_X1 U443 ( .A1(n385), .A2(n574), .ZN(n386) );
  NAND2_X1 U444 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n388), .B(KEYINPUT48), .ZN(n528) );
  XOR2_X1 U446 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n390) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n405) );
  XNOR2_X1 U449 ( .A(n405), .B(n391), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n393) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G176GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n520) );
  NAND2_X1 U458 ( .A1(n528), .A2(n520), .ZN(n403) );
  XNOR2_X1 U459 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n571) );
  XOR2_X1 U461 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U462 ( .A1(G228GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U464 ( .A(n408), .B(G204GAT), .Z(n411) );
  XNOR2_X1 U465 ( .A(n409), .B(G211GAT), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT86), .B(KEYINPUT24), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n420) );
  XOR2_X1 U471 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n417) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT85), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n438) );
  XNOR2_X1 U474 ( .A(n418), .B(n438), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n461) );
  XOR2_X1 U476 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n422) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(G57GAT), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n431) );
  XOR2_X1 U483 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n428) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT4), .B(n429), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n443) );
  XOR2_X1 U488 ( .A(G85GAT), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G29GAT), .B(G134GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U491 ( .A(G155GAT), .B(G148GAT), .Z(n435) );
  XNOR2_X1 U492 ( .A(G127GAT), .B(G120GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n518) );
  INV_X1 U498 ( .A(n518), .ZN(n570) );
  AND2_X1 U499 ( .A1(n461), .A2(n570), .ZN(n444) );
  NAND2_X1 U500 ( .A1(n571), .A2(n444), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  NOR2_X1 U502 ( .A1(n530), .A2(n447), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n448), .B(KEYINPUT123), .ZN(n567) );
  NOR2_X1 U504 ( .A1(n541), .A2(n567), .ZN(n451) );
  INV_X1 U505 ( .A(n530), .ZN(n522) );
  NOR2_X1 U506 ( .A1(n461), .A2(n522), .ZN(n453) );
  XNOR2_X1 U507 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n572) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n520), .ZN(n462) );
  NAND2_X1 U510 ( .A1(n572), .A2(n462), .ZN(n454) );
  XNOR2_X1 U511 ( .A(KEYINPUT97), .B(n454), .ZN(n459) );
  NAND2_X1 U512 ( .A1(n522), .A2(n520), .ZN(n455) );
  XNOR2_X1 U513 ( .A(KEYINPUT98), .B(n455), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n456), .A2(n461), .ZN(n457) );
  XNOR2_X1 U515 ( .A(KEYINPUT25), .B(n457), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n460), .A2(n518), .ZN(n469) );
  XNOR2_X1 U518 ( .A(n530), .B(KEYINPUT83), .ZN(n467) );
  INV_X1 U519 ( .A(n533), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n518), .A2(n462), .ZN(n463) );
  XOR2_X1 U521 ( .A(KEYINPUT94), .B(n463), .Z(n529) );
  NAND2_X1 U522 ( .A1(n464), .A2(n529), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT95), .B(n465), .Z(n466) );
  NOR2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  INV_X1 U525 ( .A(n541), .ZN(n556) );
  NOR2_X1 U526 ( .A1(n556), .A2(n581), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U528 ( .A1(n486), .A2(n471), .ZN(n506) );
  NAND2_X1 U529 ( .A1(n578), .A2(n558), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT74), .B(n472), .Z(n489) );
  AND2_X1 U531 ( .A1(n506), .A2(n489), .ZN(n482) );
  NAND2_X1 U532 ( .A1(n518), .A2(n482), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n474) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  XOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT101), .Z(n478) );
  NAND2_X1 U538 ( .A1(n482), .A2(n520), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U541 ( .A1(n482), .A2(n522), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n484) );
  NAND2_X1 U545 ( .A1(n482), .A2(n533), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n491) );
  NOR2_X1 U549 ( .A1(n486), .A2(n584), .ZN(n487) );
  NAND2_X1 U550 ( .A1(n581), .A2(n487), .ZN(n488) );
  XNOR2_X1 U551 ( .A(KEYINPUT37), .B(n488), .ZN(n515) );
  NAND2_X1 U552 ( .A1(n515), .A2(n489), .ZN(n490) );
  NAND2_X1 U553 ( .A1(n518), .A2(n501), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n493) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n520), .A2(n501), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n522), .ZN(n499) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n498) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n501), .A2(n533), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT110), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n505) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT113), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n547), .B(KEYINPUT112), .ZN(n563) );
  NAND2_X1 U571 ( .A1(n574), .A2(n563), .ZN(n516) );
  INV_X1 U572 ( .A(n506), .ZN(n507) );
  NOR2_X1 U573 ( .A1(n516), .A2(n507), .ZN(n512) );
  NAND2_X1 U574 ( .A1(n518), .A2(n512), .ZN(n508) );
  XOR2_X1 U575 ( .A(n509), .B(n508), .Z(G1332GAT) );
  NAND2_X1 U576 ( .A1(n520), .A2(n512), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n522), .A2(n512), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U581 ( .A1(n512), .A2(n533), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  INV_X1 U583 ( .A(n515), .ZN(n517) );
  NOR2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n525), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n525), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n522), .A2(n525), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(KEYINPUT114), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n525), .A2(n533), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n528), .A2(n529), .ZN(n545) );
  NOR2_X1 U596 ( .A1(n530), .A2(n545), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(n531), .Z(n532) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n558), .A2(n537), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U602 ( .A1(n537), .A2(n563), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  INV_X1 U604 ( .A(n537), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n568), .A2(n540), .ZN(n538) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n538), .Z(n539) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  INV_X1 U611 ( .A(n572), .ZN(n544) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n558), .A2(n555), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n549) );
  NAND2_X1 U616 ( .A1(n555), .A2(n547), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .Z(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(KEYINPUT120), .ZN(n554) );
  INV_X1 U621 ( .A(n581), .ZN(n552) );
  NAND2_X1 U622 ( .A1(n555), .A2(n552), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  INV_X1 U626 ( .A(n567), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n558), .A2(n564), .ZN(n559) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n561) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U631 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(n562), .Z(n566) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n574), .A2(n583), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

