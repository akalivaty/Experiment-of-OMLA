//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n208), .A2(G20), .A3(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n213), .B2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n215), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(new_n229));
  OAI211_X1 g0029(.A(new_n211), .B(new_n219), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT83), .ZN(new_n247));
  INV_X1    g0047(.A(G169), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OR2_X1    g0052(.A1(KEYINPUT5), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT5), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n210), .B2(new_n259), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n256), .A2(G270), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n263), .A2(new_n265), .A3(G264), .A4(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G303), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n266), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n249), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n248), .B1(new_n261), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G20), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n215), .A2(new_n274), .A3(G1), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n209), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n250), .A2(G33), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n276), .A2(G116), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G116), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n277), .A2(new_n209), .B1(G20), .B2(new_n282), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G283), .ZN(new_n285));
  INV_X1    g0085(.A(G97), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n274), .C1(G33), .C2(new_n286), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n284), .A2(KEYINPUT20), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT20), .B1(new_n284), .B2(new_n287), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n281), .B(new_n283), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n247), .B(KEYINPUT21), .C1(new_n273), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n261), .A2(new_n272), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G169), .A3(new_n290), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT21), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT83), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n290), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n271), .A2(new_n249), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n257), .A2(new_n260), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n255), .A2(new_n252), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G270), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(KEYINPUT21), .B(G169), .C1(new_n297), .C2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n261), .A2(new_n272), .A3(G179), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n291), .A2(new_n295), .B1(new_n306), .B2(KEYINPUT82), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n306), .A2(KEYINPUT82), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n292), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n261), .B2(new_n272), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n310), .A2(new_n290), .A3(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n307), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n263), .A2(new_n265), .A3(G226), .A4(G1698), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n263), .A2(new_n265), .A3(G223), .A4(new_n267), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n249), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n300), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G41), .ZN(new_n323));
  INV_X1    g0123(.A(G45), .ZN(new_n324));
  AOI21_X1  g0124(.A(G1), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n322), .A2(G232), .B1(new_n260), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n300), .A3(G274), .ZN(new_n329));
  INV_X1    g0129(.A(G232), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n249), .B2(new_n318), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n328), .B1(new_n332), .B2(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n263), .A2(new_n265), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT7), .B1(new_n334), .B2(new_n274), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT7), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n336), .B(G20), .C1(new_n263), .C2(new_n265), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  INV_X1    g0139(.A(G68), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n341), .B2(new_n201), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G20), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G159), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n336), .B1(new_n270), .B2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n334), .A2(KEYINPUT7), .A3(new_n274), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n351), .B2(new_n345), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n352), .A3(new_n278), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n278), .B1(new_n250), .B2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n339), .A2(KEYINPUT8), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT8), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G58), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT67), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n339), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n276), .B2(new_n361), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n333), .B1(new_n353), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT18), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n319), .A2(new_n326), .A3(new_n309), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n332), .B2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT76), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n353), .A2(new_n368), .A3(new_n369), .A4(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n353), .A2(new_n368), .A3(new_n364), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(KEYINPUT17), .C1(KEYINPUT75), .C2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n366), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n262), .A2(KEYINPUT68), .A3(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n274), .A2(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT68), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n359), .A2(new_n378), .A3(new_n360), .A4(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n343), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n279), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n275), .A2(new_n202), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n279), .B1(G1), .B2(new_n274), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n202), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G226), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n329), .B1(new_n321), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n270), .A2(G222), .A3(new_n267), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n270), .A2(G223), .A3(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n334), .A2(G77), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n394), .B2(new_n249), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n388), .B1(G169), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n395), .A2(new_n327), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(G190), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT10), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n311), .C2(new_n395), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT9), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n387), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT71), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT9), .B1(new_n383), .B2(new_n386), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT72), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n406), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT9), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT71), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT72), .A3(new_n402), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n413), .A2(new_n414), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n399), .B1(new_n311), .B2(new_n395), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT10), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n398), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT77), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n366), .A2(new_n373), .A3(new_n423), .A4(new_n375), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n275), .A2(new_n340), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT12), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(KEYINPUT12), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(KEYINPUT74), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(KEYINPUT74), .B2(new_n430), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT11), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n378), .A2(G77), .A3(new_n380), .ZN(new_n434));
  INV_X1    g0234(.A(new_n343), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n435), .A2(new_n202), .B1(new_n274), .B2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n278), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n432), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n433), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n340), .B2(new_n385), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n334), .A2(new_n330), .A3(new_n267), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n263), .A2(new_n265), .A3(G226), .A4(new_n267), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n249), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT13), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n322), .A2(G238), .B1(new_n260), .B2(new_n325), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n442), .B(G169), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT13), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n452), .B1(new_n327), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n442), .B1(new_n456), .B2(G169), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n441), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n438), .A2(new_n440), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(G200), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(new_n309), .C2(new_n456), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(new_n270), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n334), .A2(new_n330), .A3(G1698), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n249), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n220), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n322), .A2(new_n468), .B1(new_n260), .B2(new_n325), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G200), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(G190), .A3(new_n469), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT8), .B(G58), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n473), .A2(new_n435), .B1(new_n274), .B2(new_n221), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT69), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT15), .B(G87), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n474), .A2(new_n475), .B1(new_n379), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n474), .A2(new_n475), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n278), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OR3_X1    g0279(.A1(new_n276), .A2(KEYINPUT70), .A3(G77), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT70), .B1(new_n276), .B2(G77), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n480), .A2(new_n481), .B1(G77), .B2(new_n354), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n471), .A2(new_n472), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(new_n248), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n467), .A2(new_n327), .A3(new_n469), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n459), .A2(new_n462), .A3(new_n488), .ZN(new_n489));
  AND4_X1   g0289(.A1(new_n377), .A2(new_n422), .A3(new_n424), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G257), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n298), .B1(new_n301), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(new_n267), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n285), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT78), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n300), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n497), .A2(new_n285), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT78), .A3(new_n495), .A4(new_n496), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n492), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n327), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n286), .A3(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n508), .A2(new_n274), .B1(new_n221), .B2(new_n435), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n464), .B1(new_n349), .B2(new_n350), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n278), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n275), .A2(new_n286), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G97), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n504), .B(new_n516), .C1(G169), .C2(new_n503), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n503), .A2(G190), .ZN(new_n518));
  INV_X1    g0318(.A(new_n516), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n311), .C2(new_n503), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n270), .A2(G250), .A3(new_n267), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n262), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n249), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n256), .A2(G264), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n298), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n248), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(KEYINPUT84), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n270), .A2(new_n274), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n270), .A2(KEYINPUT22), .A3(new_n274), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(G20), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT23), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n274), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n464), .A2(KEYINPUT23), .A3(G20), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n534), .A2(new_n544), .A3(new_n535), .A4(new_n541), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n279), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT25), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(KEYINPUT85), .ZN(new_n548));
  AOI21_X1  g0348(.A(G107), .B1(new_n547), .B2(KEYINPUT85), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n275), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n275), .B2(new_n549), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n513), .A2(new_n464), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI221_X1 g0352(.A(new_n529), .B1(G179), .B2(new_n528), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n274), .B1(new_n445), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(G97), .A2(G107), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n530), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT81), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n270), .A2(new_n274), .A3(G68), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n554), .B1(new_n379), .B2(new_n286), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n278), .ZN(new_n564));
  INV_X1    g0364(.A(new_n476), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n276), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n514), .A2(new_n565), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(G244), .A2(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n263), .A2(new_n265), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n263), .A2(new_n265), .A3(G238), .A4(new_n267), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n263), .A2(new_n265), .A3(new_n570), .A4(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(new_n536), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n574), .A2(new_n536), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(KEYINPUT80), .A3(new_n575), .A4(new_n573), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n300), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n260), .A2(new_n252), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n300), .A2(G250), .A3(new_n251), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n248), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n578), .A2(new_n580), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n249), .ZN(new_n587));
  INV_X1    g0387(.A(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n569), .B(new_n585), .C1(new_n589), .C2(G179), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n546), .A2(new_n552), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n528), .A2(G190), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n528), .A2(new_n311), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(G190), .A3(new_n588), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n513), .A2(new_n530), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n566), .B(new_n596), .C1(new_n563), .C2(new_n278), .ZN(new_n597));
  OAI21_X1  g0397(.A(G200), .B1(new_n581), .B2(new_n584), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n553), .A2(new_n590), .A3(new_n594), .A4(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n314), .A2(new_n490), .A3(new_n521), .A4(new_n600), .ZN(G372));
  INV_X1    g0401(.A(KEYINPUT86), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n581), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n581), .A2(new_n602), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n588), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n248), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n581), .A2(new_n584), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n327), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n569), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n517), .A2(new_n520), .A3(new_n594), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n595), .A2(new_n597), .ZN(new_n613));
  INV_X1    g0413(.A(new_n605), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n584), .B1(new_n614), .B2(new_n603), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n311), .ZN(new_n616));
  INV_X1    g0416(.A(new_n291), .ZN(new_n617));
  INV_X1    g0417(.A(new_n295), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n306), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n553), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n612), .A2(new_n611), .A3(new_n616), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n606), .A2(G200), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n610), .A2(new_n607), .B1(new_n623), .B2(new_n613), .ZN(new_n624));
  INV_X1    g0424(.A(new_n517), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT26), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n590), .A2(new_n599), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n627), .A2(new_n628), .A3(new_n517), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n611), .B(new_n622), .C1(new_n626), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n490), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n487), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n462), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n459), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT17), .B1(new_n372), .B2(KEYINPUT75), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n375), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n366), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n411), .B(new_n401), .C1(new_n415), .C2(new_n407), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT72), .B1(new_n416), .B2(new_n402), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n421), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n398), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g0443(.A(new_n643), .B(KEYINPUT87), .Z(G369));
  NAND2_X1  g0444(.A1(new_n619), .A2(new_n620), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n250), .A2(new_n274), .A3(G13), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  INV_X1    g0448(.A(G213), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G343), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n290), .ZN(new_n653));
  MUX2_X1   g0453(.A(new_n645), .B(new_n314), .S(new_n653), .Z(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n594), .A2(new_n553), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n591), .B2(new_n651), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n553), .B2(new_n651), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n651), .B(KEYINPUT88), .Z(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n553), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n307), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n306), .A2(KEYINPUT82), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n652), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n657), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n660), .A2(new_n667), .ZN(G399));
  NOR2_X1   g0468(.A1(new_n557), .A2(G116), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT89), .ZN(new_n670));
  INV_X1    g0470(.A(new_n217), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n672), .A3(new_n250), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n208), .B2(new_n672), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT28), .Z(new_n675));
  NAND3_X1  g0475(.A1(new_n611), .A2(new_n616), .A3(new_n625), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n629), .B1(new_n676), .B2(new_n628), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n622), .A2(new_n611), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n661), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n611), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n611), .A2(new_n616), .A3(KEYINPUT26), .A4(new_n625), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n628), .B1(new_n627), .B2(new_n517), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT82), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n620), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n619), .A2(new_n687), .A3(new_n665), .A4(new_n553), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n664), .A2(KEYINPUT92), .A3(new_n665), .A4(new_n553), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n624), .A2(new_n690), .A3(new_n612), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .A3(new_n651), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n681), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n305), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n261), .A2(new_n272), .A3(KEYINPUT90), .A4(G179), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n526), .A2(new_n527), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n699), .A2(new_n608), .A3(new_n503), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n581), .A2(new_n700), .A3(new_n584), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n699), .A3(new_n705), .A4(new_n503), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n528), .A2(new_n327), .A3(new_n292), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n503), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n606), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n651), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT91), .B1(new_n711), .B2(KEYINPUT31), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n703), .A2(new_n706), .B1(new_n606), .B2(new_n709), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n651), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n600), .A2(new_n314), .A3(new_n521), .A4(new_n661), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n707), .A2(new_n710), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n712), .A2(new_n716), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n695), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n675), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n215), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n250), .B1(new_n725), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n672), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n656), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n654), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n209), .B1(G20), .B2(new_n248), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n274), .A2(new_n327), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G200), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G190), .ZN(new_n734));
  INV_X1    g0534(.A(G317), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT33), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(KEYINPUT33), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n309), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n274), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n274), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n738), .B1(new_n524), .B2(new_n740), .C1(new_n269), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n270), .B1(new_n746), .B2(G329), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n732), .A2(new_n744), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n732), .A2(G190), .A3(new_n311), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n747), .B1(new_n748), .B2(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n733), .A2(new_n309), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G326), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n741), .A2(new_n309), .A3(G200), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n743), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT94), .Z(new_n759));
  NAND2_X1  g0559(.A1(new_n746), .A2(G159), .ZN(new_n760));
  INV_X1    g0560(.A(new_n740), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n760), .A2(KEYINPUT32), .B1(new_n761), .B2(G97), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(KEYINPUT32), .B2(new_n760), .ZN(new_n763));
  INV_X1    g0563(.A(new_n753), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n764), .A2(new_n202), .B1(new_n742), .B2(new_n530), .ZN(new_n765));
  INV_X1    g0565(.A(new_n734), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n766), .A2(new_n340), .B1(new_n756), .B2(new_n464), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n270), .B1(new_n749), .B2(new_n221), .C1(new_n339), .C2(new_n751), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n763), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n731), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n217), .A2(G355), .A3(new_n270), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G116), .B2(new_n217), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n242), .A2(new_n324), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n217), .A2(new_n334), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n324), .B2(new_n208), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT93), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n731), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n728), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n770), .B(new_n786), .C1(new_n654), .C2(new_n780), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n730), .A2(new_n787), .ZN(G396));
  OAI22_X1  g0588(.A1(new_n740), .A2(new_n286), .B1(new_n751), .B2(new_n524), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT95), .Z(new_n790));
  OAI21_X1  g0590(.A(new_n334), .B1(new_n745), .B2(new_n748), .ZN(new_n791));
  INV_X1    g0591(.A(new_n749), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(G116), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n756), .A2(new_n530), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G303), .B2(new_n753), .ZN(new_n795));
  INV_X1    g0595(.A(new_n742), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n734), .A2(G283), .B1(new_n796), .B2(G107), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n790), .A2(new_n793), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n756), .A2(new_n340), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n334), .B1(new_n746), .B2(G132), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n339), .B2(new_n740), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n799), .B(new_n801), .C1(G50), .C2(new_n796), .ZN(new_n802));
  INV_X1    g0602(.A(new_n751), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G143), .B1(new_n792), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n764), .B2(new_n805), .C1(new_n806), .C2(new_n766), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n798), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n731), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n731), .A2(new_n777), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n785), .B1(new_n221), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n485), .A2(new_n652), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n632), .B1(new_n483), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n487), .A2(new_n652), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n813), .B(new_n815), .C1(new_n819), .C2(new_n778), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n679), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n662), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n630), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n728), .B1(new_n825), .B2(new_n721), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n721), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n820), .B1(new_n827), .B2(new_n828), .ZN(G384));
  NOR2_X1   g0629(.A1(new_n725), .A2(new_n250), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n650), .B(KEYINPUT98), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n366), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n818), .B1(new_n630), .B2(new_n823), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n459), .A2(new_n462), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n834), .A2(new_n441), .A3(new_n652), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n459), .B(new_n462), .C1(new_n460), .C2(new_n651), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n353), .A2(new_n364), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n840), .A2(new_n650), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT18), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n365), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n637), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n338), .A2(new_n346), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n279), .B1(new_n845), .B2(new_n348), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n363), .B1(new_n846), .B2(new_n347), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n372), .B1(new_n847), .B2(new_n333), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n848), .B2(new_n841), .ZN(new_n849));
  INV_X1    g0649(.A(new_n333), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n840), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n840), .A2(new_n831), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .A4(new_n372), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n849), .A2(KEYINPUT99), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT99), .B1(new_n849), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT38), .B(new_n844), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n832), .B1(new_n839), .B2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n459), .A2(new_n652), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n860), .ZN(new_n865));
  INV_X1    g0665(.A(new_n852), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n376), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n848), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n854), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT99), .ZN(new_n872));
  INV_X1    g0672(.A(new_n372), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(new_n365), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n840), .A2(new_n650), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n853), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n854), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n849), .A2(KEYINPUT99), .A3(new_n854), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT38), .A4(new_n844), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n870), .B1(new_n871), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n864), .B(new_n865), .C1(new_n883), .C2(KEYINPUT39), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n862), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n681), .A2(new_n694), .A3(new_n490), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n642), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n714), .B1(new_n715), .B2(new_n651), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n717), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n821), .B1(new_n835), .B2(new_n836), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n860), .B2(new_n859), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n892), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n894), .A2(KEYINPUT40), .B1(new_n883), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n490), .A2(new_n891), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(G330), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n830), .B1(new_n888), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n888), .B2(new_n901), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT35), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n508), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n905), .A2(G20), .A3(G116), .A4(new_n210), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT96), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n906), .A2(new_n907), .B1(new_n904), .B2(new_n508), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n207), .A2(new_n221), .A3(new_n341), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n340), .A2(G50), .ZN(new_n913));
  OAI211_X1 g0713(.A(G1), .B(new_n215), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(new_n911), .A3(new_n914), .ZN(G367));
  NOR2_X1   g0715(.A1(new_n238), .A2(new_n774), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n782), .B1(new_n217), .B2(new_n476), .ZN(new_n917));
  INV_X1    g0717(.A(G159), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n766), .A2(new_n918), .B1(new_n742), .B2(new_n339), .ZN(new_n919));
  XNOR2_X1  g0719(.A(KEYINPUT104), .B(G137), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n751), .A2(new_n806), .B1(new_n745), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n334), .B(new_n921), .C1(G50), .C2(new_n792), .ZN(new_n922));
  INV_X1    g0722(.A(new_n756), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G77), .ZN(new_n924));
  INV_X1    g0724(.A(G143), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n922), .B(new_n924), .C1(new_n925), .C2(new_n764), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n919), .B(new_n926), .C1(G68), .C2(new_n761), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT105), .Z(new_n928));
  NOR2_X1   g0728(.A1(new_n756), .A2(new_n286), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n764), .A2(new_n748), .B1(new_n464), .B2(new_n740), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(G294), .C2(new_n734), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n749), .A2(new_n755), .B1(new_n745), .B2(new_n735), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n334), .B1(new_n751), .B2(new_n269), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT46), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n796), .A2(G116), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n931), .B(new_n936), .C1(new_n934), .C2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT47), .Z(new_n939));
  INV_X1    g0739(.A(new_n731), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n728), .B1(new_n916), .B2(new_n917), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n624), .B1(new_n597), .B2(new_n651), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n611), .A2(new_n597), .A3(new_n651), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT101), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(KEYINPUT101), .B2(new_n943), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n781), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT106), .Z(new_n947));
  OAI21_X1  g0747(.A(new_n521), .B1(new_n519), .B2(new_n661), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT103), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n625), .A2(new_n662), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n667), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT45), .Z(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n667), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT44), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n660), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n666), .A2(new_n657), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n659), .B2(new_n666), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n656), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n723), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n660), .A3(new_n955), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(new_n723), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n672), .B(KEYINPUT41), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n726), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n958), .B1(new_n949), .B2(new_n950), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT42), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n517), .B1(new_n949), .B2(new_n553), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n661), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT43), .B1(new_n945), .B2(KEYINPUT102), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(KEYINPUT102), .B2(new_n945), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(new_n974), .C1(new_n975), .C2(new_n945), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n972), .B2(new_n974), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n951), .A2(new_n656), .A3(new_n659), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n977), .B(new_n978), .Z(new_n979));
  AOI21_X1  g0779(.A(new_n947), .B1(new_n967), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(G387));
  NOR2_X1   g0781(.A1(new_n659), .A2(new_n780), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n235), .A2(new_n324), .A3(new_n270), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n473), .A2(KEYINPUT50), .A3(G50), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT50), .B1(new_n473), .B2(G50), .ZN(new_n985));
  AOI21_X1  g0785(.A(G45), .B1(G68), .B2(G77), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n670), .B1(new_n987), .B2(new_n334), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n217), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n782), .C1(new_n464), .C2(new_n217), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n728), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n742), .A2(new_n221), .B1(new_n745), .B2(new_n806), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT107), .Z(new_n993));
  NOR2_X1   g0793(.A1(new_n740), .A2(new_n476), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n929), .B(new_n994), .C1(G159), .C2(new_n753), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n270), .B1(new_n749), .B2(new_n340), .C1(new_n202), .C2(new_n751), .ZN(new_n996));
  INV_X1    g0796(.A(new_n361), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n734), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n270), .B1(new_n746), .B2(G326), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n740), .A2(new_n755), .B1(new_n742), .B2(new_n524), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n803), .A2(G317), .B1(new_n792), .B2(G303), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n764), .B2(new_n750), .C1(new_n748), .C2(new_n766), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT108), .Z(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1000), .B1(new_n282), .B2(new_n756), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n999), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n982), .B(new_n991), .C1(new_n1011), .C2(new_n731), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n960), .B2(new_n727), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n961), .A2(new_n672), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n723), .A2(new_n960), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(G393));
  INV_X1    g0816(.A(KEYINPUT109), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n963), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(new_n956), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n672), .B(new_n964), .C1(new_n1019), .C2(new_n962), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n727), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G317), .A2(new_n753), .B1(new_n803), .B2(G311), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n334), .B1(new_n745), .B2(new_n750), .C1(new_n524), .C2(new_n749), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n766), .A2(new_n269), .B1(new_n756), .B2(new_n464), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n740), .A2(new_n282), .B1(new_n742), .B2(new_n755), .ZN(new_n1027));
  OR4_X1    g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n764), .A2(new_n806), .B1(new_n918), .B2(new_n751), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n270), .B1(new_n745), .B2(new_n925), .C1(new_n473), .C2(new_n749), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n766), .A2(new_n202), .B1(new_n742), .B2(new_n340), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n740), .A2(new_n221), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1033), .A2(new_n794), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1030), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n940), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n245), .A2(new_n774), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n783), .B1(G97), .B2(new_n671), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n785), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n951), .B2(new_n780), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1020), .A2(new_n1021), .A3(new_n1041), .ZN(G390));
  OAI21_X1  g0842(.A(new_n863), .B1(new_n833), .B2(new_n838), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n865), .B1(new_n883), .B2(KEYINPUT39), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n883), .A2(new_n864), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n652), .B1(new_n685), .B2(new_n692), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n817), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n818), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1046), .B1(new_n838), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n720), .A2(G330), .A3(new_n819), .A4(new_n837), .ZN(new_n1051));
  INV_X1    g0851(.A(G330), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n821), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n891), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT111), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1045), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1054), .A2(new_n838), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT111), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n398), .ZN(new_n1061));
  AND4_X1   g0861(.A1(new_n424), .A2(new_n489), .A3(new_n641), .A4(new_n1061), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n891), .A2(new_n1062), .A3(G330), .A4(new_n377), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT112), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT112), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n490), .A2(new_n1065), .A3(G330), .A4(new_n891), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1067), .A2(new_n642), .A3(new_n886), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1054), .A2(new_n838), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1049), .A2(new_n1051), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n720), .A2(G330), .A3(new_n819), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1058), .B1(new_n838), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1072), .B2(new_n833), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1057), .A2(new_n1060), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n672), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT113), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1045), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT113), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1049), .A2(new_n838), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(new_n1046), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1080), .C1(new_n1082), .C2(new_n1059), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1067), .A2(new_n886), .A3(new_n642), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n833), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1071), .A2(new_n838), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n1058), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1087), .B2(new_n1070), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1074), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1078), .A2(new_n1083), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n814), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G97), .A2(new_n792), .B1(new_n746), .B2(G294), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n282), .B2(new_n751), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n464), .A2(new_n766), .B1(new_n764), .B2(new_n755), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n799), .A4(new_n1034), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n334), .B1(new_n742), .B2(new_n530), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT116), .Z(new_n1100));
  AOI22_X1  g0900(.A1(new_n803), .A2(G132), .B1(new_n746), .B2(G125), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n270), .C1(new_n749), .C2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n766), .A2(new_n920), .B1(new_n918), .B2(new_n740), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n764), .A2(new_n1105), .B1(new_n756), .B2(new_n202), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n742), .A2(new_n806), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1098), .A2(new_n1100), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n728), .B1(new_n997), .B2(new_n1094), .C1(new_n1110), .C2(new_n940), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1044), .B2(new_n777), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n727), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1079), .B1(new_n1082), .B2(new_n1059), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT115), .B1(new_n1116), .B2(new_n726), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1112), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1093), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(KEYINPUT120), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n896), .B2(new_n1052), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n861), .A2(new_n891), .A3(new_n892), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT40), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n871), .A2(new_n882), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n870), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n895), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1130), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n422), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1132), .B(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n388), .A2(new_n650), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT118), .Z(new_n1137));
  AND2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1122), .A2(new_n1131), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n885), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n897), .A2(new_n1143), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1120), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n885), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(KEYINPUT120), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1151), .A3(new_n727), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1143), .A2(new_n777), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n334), .B2(new_n323), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n923), .A2(G58), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n764), .B2(new_n282), .C1(new_n286), .C2(new_n766), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n323), .B(new_n334), .C1(new_n745), .C2(new_n755), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n751), .A2(new_n464), .B1(new_n749), .B2(new_n476), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n740), .A2(new_n340), .B1(new_n742), .B2(new_n221), .ZN(new_n1160));
  OR4_X1    g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT58), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1155), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n742), .A2(new_n1102), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT117), .Z(new_n1165));
  OAI22_X1  g0965(.A1(new_n751), .A2(new_n1105), .B1(new_n749), .B2(new_n805), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G125), .B2(new_n753), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G150), .A2(new_n761), .B1(new_n734), .B2(G132), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n923), .A2(G159), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1163), .B1(new_n1162), .B2(new_n1161), .C1(new_n1170), .C2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n731), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n785), .B1(new_n202), .B2(new_n814), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1153), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1152), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1088), .B(new_n1079), .C1(new_n1082), .C2(new_n1059), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1182), .A2(KEYINPUT121), .A3(new_n1068), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT121), .B1(new_n1182), .B2(new_n1068), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1180), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT121), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1075), .B2(new_n1084), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1182), .A2(KEYINPUT121), .A3(new_n1068), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1145), .A2(new_n1146), .A3(new_n1180), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1076), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1179), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(G375));
  NAND2_X1  g0994(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1195), .A2(new_n966), .A3(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT122), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n838), .A2(new_n777), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n728), .B1(G68), .B2(new_n1094), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n734), .A2(G116), .B1(new_n792), .B2(G107), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT123), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n334), .B1(new_n745), .B2(new_n269), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n803), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n753), .A2(G294), .B1(new_n796), .B2(G97), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n994), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n924), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n753), .A2(G132), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n918), .B2(new_n742), .C1(new_n766), .C2(new_n1102), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n920), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n803), .A2(new_n1210), .B1(new_n792), .B2(G150), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n334), .B1(new_n746), .B2(G128), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n761), .A2(G50), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n1156), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1202), .A2(new_n1207), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1200), .B1(new_n1215), .B2(new_n731), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1073), .A2(new_n727), .B1(new_n1199), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1198), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1093), .A2(new_n1118), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n980), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1222), .A2(G375), .A3(G381), .ZN(G407));
  NOR2_X1   g1023(.A1(new_n649), .A2(G343), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1193), .A2(new_n1220), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G407), .A2(G213), .A3(new_n1225), .ZN(G409));
  NOR2_X1   g1026(.A1(new_n980), .A2(G390), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n980), .A2(G390), .ZN(new_n1229));
  XOR2_X1   g1029(.A(G393), .B(G396), .Z(new_n1230));
  NAND4_X1  g1030(.A1(new_n1228), .A2(KEYINPUT127), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT127), .B1(new_n980), .B2(G390), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1230), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1232), .A2(new_n1227), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT61), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1074), .A2(KEYINPUT60), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1196), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n672), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1238), .A2(new_n1196), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1217), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G384), .B(new_n1217), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1224), .ZN(new_n1248));
  INV_X1    g1048(.A(G2897), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1244), .A2(new_n1246), .B1(new_n1249), .B2(new_n1248), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n966), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1190), .A2(new_n1254), .A3(new_n1151), .A4(new_n1147), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1178), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n727), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G378), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1193), .B2(G378), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1260), .B2(new_n1224), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1247), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1260), .A2(new_n1224), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1237), .B(new_n1261), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1220), .B(new_n1179), .C1(new_n1186), .C2(new_n1192), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1248), .B(new_n1247), .C1(new_n1266), .C2(new_n1259), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1236), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT125), .B1(new_n1260), .B2(new_n1224), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1271), .B(new_n1248), .C1(new_n1266), .C2(new_n1259), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1272), .A3(new_n1253), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT126), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1270), .A2(new_n1272), .A3(new_n1275), .A4(new_n1253), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT63), .B1(new_n1263), .B2(KEYINPUT124), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1231), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT124), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1267), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1269), .B1(new_n1277), .B2(new_n1283), .ZN(G405));
  NOR2_X1   g1084(.A1(new_n1193), .A2(G378), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1285), .A2(new_n1266), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1262), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1236), .ZN(G402));
endmodule


