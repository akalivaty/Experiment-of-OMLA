//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G101), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT82), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n189), .A2(new_n192), .A3(new_n197), .A4(new_n193), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n200), .A3(G101), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n204));
  INV_X1    g018(.A(G113), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n206), .A2(new_n207), .B1(KEYINPUT2), .B2(G113), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G116), .B(G119), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n208), .B1(new_n211), .B2(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n195), .A2(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n188), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n191), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n198), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n223), .A2(KEYINPUT5), .A3(G119), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(new_n205), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n208), .A2(new_n210), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT86), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT6), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n232), .A3(new_n228), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n230), .A2(new_n231), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT88), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n229), .B2(KEYINPUT86), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n231), .A4(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G125), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT66), .B(G128), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(G143), .B2(new_n242), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n246), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n253), .B1(G125), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G224), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G953), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT89), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n262), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n230), .A2(new_n233), .A3(new_n235), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n217), .A2(new_n228), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n231), .B1(new_n268), .B2(new_n234), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT87), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n267), .A2(KEYINPUT87), .A3(new_n269), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n241), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G210), .B1(G237), .B2(G902), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT7), .B1(new_n263), .B2(G953), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n262), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n262), .A2(new_n275), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n198), .A2(new_n220), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n222), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n210), .A2(KEYINPUT90), .A3(KEYINPUT5), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n225), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n282), .B2(new_n227), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n227), .A2(new_n278), .A3(new_n226), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n234), .B(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n276), .B(new_n277), .C1(new_n283), .C2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n229), .A2(new_n235), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n274), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT91), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n272), .A2(new_n273), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n273), .B1(new_n272), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G221), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n296), .B2(new_n274), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT1), .B1(new_n244), .B2(G146), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n300), .A2(G128), .B1(new_n243), .B2(new_n245), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n259), .A2(new_n243), .A3(new_n245), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n303), .A2(new_n278), .A3(KEYINPUT83), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n246), .B1(new_n256), .B2(new_n258), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n260), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n221), .B2(new_n307), .ZN(new_n308));
  OAI22_X1  g122(.A1(new_n304), .A2(new_n308), .B1(new_n261), .B2(new_n221), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G134), .ZN(new_n311));
  INV_X1    g125(.A(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT11), .B1(new_n312), .B2(G137), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT11), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n310), .A3(G134), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(G137), .ZN(new_n320));
  AND4_X1   g134(.A1(KEYINPUT64), .A2(new_n319), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT64), .B1(new_n316), .B2(new_n317), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT12), .B1(new_n309), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT83), .B1(new_n303), .B2(new_n278), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n221), .A2(new_n307), .A3(new_n305), .ZN(new_n326));
  INV_X1    g140(.A(new_n261), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n278), .ZN(new_n328));
  INV_X1    g142(.A(new_n323), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT12), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n299), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G140), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G227), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n309), .A2(KEYINPUT12), .A3(new_n323), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n330), .B1(new_n328), .B2(new_n329), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT85), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n332), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n304), .B2(new_n308), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n252), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n216), .A3(new_n202), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n221), .A2(new_n261), .A3(KEYINPUT10), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(new_n350), .A3(new_n329), .A4(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n325), .A2(new_n326), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(new_n344), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n357), .A2(KEYINPUT84), .A3(new_n329), .A4(new_n350), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n350), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n354), .A2(new_n358), .B1(new_n361), .B2(new_n323), .ZN(new_n362));
  OAI22_X1  g176(.A1(new_n343), .A2(new_n360), .B1(new_n362), .B2(new_n339), .ZN(new_n363));
  INV_X1    g177(.A(G469), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n274), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n274), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n361), .A2(new_n323), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n354), .A2(new_n358), .B1(new_n340), .B2(new_n341), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n370), .B(new_n339), .C1(KEYINPUT81), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n338), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n364), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n298), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT92), .B(G143), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n334), .A3(G214), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G237), .A2(G953), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n381), .A2(G214), .B1(new_n382), .B2(G143), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT17), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(KEYINPUT92), .B2(new_n244), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n317), .C1(new_n379), .C2(new_n377), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(KEYINPUT17), .B(G131), .C1(new_n380), .C2(new_n383), .ZN(new_n389));
  INV_X1    g203(.A(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G125), .ZN(new_n391));
  INV_X1    g205(.A(G125), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G140), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n392), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G146), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT75), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G146), .B1(new_n394), .B2(new_n395), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI211_X1 g214(.A(new_n397), .B(G146), .C1(new_n394), .C2(new_n395), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n388), .B(new_n389), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G113), .B(G122), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(new_n188), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n386), .B(new_n405), .C1(new_n379), .C2(new_n377), .ZN(new_n406));
  XNOR2_X1  g220(.A(G125), .B(G140), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n242), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n408), .C1(new_n384), .C2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n402), .A2(new_n404), .A3(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n384), .A2(new_n387), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n407), .B(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n396), .B1(new_n414), .B2(G146), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n410), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n404), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(KEYINPUT93), .A3(new_n420), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(new_n421), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT20), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n411), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n404), .B1(new_n402), .B2(new_n410), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n274), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G475), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT94), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT94), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(new_n435), .A3(new_n432), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n223), .B2(G122), .ZN(new_n439));
  INV_X1    g253(.A(G122), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT95), .A3(G116), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n439), .A2(new_n441), .B1(new_n223), .B2(G122), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(new_n191), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n191), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n254), .A2(G143), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT96), .B1(new_n258), .B2(G143), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n244), .A3(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n312), .A3(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT97), .B(KEYINPUT13), .Z(new_n452));
  OAI21_X1  g266(.A(new_n446), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT98), .B1(new_n452), .B2(new_n450), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n450), .A3(KEYINPUT98), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n445), .B(new_n451), .C1(new_n457), .C2(new_n312), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n442), .B1(KEYINPUT14), .B2(new_n191), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n446), .A2(new_n312), .A3(new_n450), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n312), .B1(new_n446), .B2(new_n450), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n439), .A2(new_n441), .ZN(new_n463));
  AOI211_X1 g277(.A(new_n191), .B(new_n442), .C1(KEYINPUT14), .C2(new_n463), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G217), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n295), .A2(new_n466), .A3(G953), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n467), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n451), .B1(new_n443), .B2(new_n444), .ZN(new_n470));
  INV_X1    g284(.A(new_n453), .ZN(new_n471));
  INV_X1    g285(.A(new_n456), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n472), .B2(new_n454), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n473), .B2(G134), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n462), .A2(new_n464), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(G902), .B(new_n479), .C1(new_n468), .C2(new_n476), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n437), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n468), .A2(new_n476), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n274), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n479), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n477), .A2(new_n480), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT99), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT100), .B(G952), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G953), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(G902), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT21), .B(G898), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n434), .A2(new_n436), .A3(new_n489), .A4(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n293), .A2(new_n376), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n321), .A2(new_n322), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n320), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n310), .A2(G134), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n312), .A2(KEYINPUT65), .A3(G137), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G131), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n261), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT67), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n252), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n323), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n257), .A2(new_n260), .B1(new_n506), .B2(G131), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT67), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n512), .B(new_n513), .C1(new_n322), .C2(new_n321), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n512), .B1(new_n322), .B2(new_n321), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n349), .A2(new_n323), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n512), .B(KEYINPUT71), .C1(new_n322), .C2(new_n321), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT30), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(new_n215), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n215), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n520), .A2(new_n521), .A3(new_n525), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n381), .A2(G210), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT27), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT26), .B(G101), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n524), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n524), .A2(KEYINPUT31), .A3(new_n526), .A4(new_n530), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n530), .B(KEYINPUT72), .Z(new_n536));
  INV_X1    g350(.A(new_n526), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n518), .A2(KEYINPUT67), .B1(new_n323), .B2(new_n510), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n525), .B1(new_n538), .B2(new_n514), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT28), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n518), .A2(new_n525), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT28), .B1(new_n541), .B2(new_n521), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n536), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n535), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n521), .A2(new_n522), .ZN(new_n549));
  INV_X1    g363(.A(new_n520), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n215), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n526), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n542), .B1(new_n552), .B2(KEYINPUT28), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT29), .A3(new_n530), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n274), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT28), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n515), .A2(new_n215), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n526), .ZN(new_n558));
  INV_X1    g372(.A(new_n536), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n558), .A2(new_n559), .A3(new_n542), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n530), .B1(new_n524), .B2(new_n526), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(G472), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT32), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n544), .B1(new_n533), .B2(new_n534), .ZN(new_n565));
  INV_X1    g379(.A(new_n547), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n548), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n466), .B1(G234), .B2(new_n274), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT66), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G128), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n572), .A3(G119), .ZN(new_n573));
  INV_X1    g387(.A(G119), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G128), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT73), .ZN(new_n577));
  INV_X1    g391(.A(G110), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(KEYINPUT24), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(KEYINPUT24), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT74), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT24), .B(G110), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n573), .A2(new_n586), .A3(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT76), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n574), .B2(G128), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n591), .A2(new_n575), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(new_n578), .C1(new_n590), .C2(new_n573), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n589), .B1(new_n588), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n407), .A2(new_n242), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n396), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n401), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n577), .A2(new_n587), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n584), .A3(new_n581), .ZN(new_n601));
  INV_X1    g415(.A(new_n400), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n592), .B1(new_n590), .B2(new_n573), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G110), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT77), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n588), .A2(new_n593), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT76), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n396), .A3(new_n609), .A4(new_n596), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT77), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n601), .A2(new_n602), .A3(new_n599), .A4(new_n604), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT22), .B(G137), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n606), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n610), .A2(new_n612), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT77), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT25), .B1(new_n621), .B2(new_n274), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT25), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n623), .B(G902), .C1(new_n618), .C2(new_n620), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n569), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n569), .A2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n568), .A2(new_n628), .A3(KEYINPUT78), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT78), .B1(new_n568), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n500), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  OAI21_X1  g446(.A(G472), .B1(new_n565), .B2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n546), .A2(new_n547), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n625), .A2(new_n627), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n376), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n434), .A2(new_n436), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n484), .A2(KEYINPUT33), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n484), .A2(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(G478), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n478), .A2(new_n274), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n477), .B2(new_n478), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n638), .A2(new_n498), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n293), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n427), .A2(new_n422), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n432), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n489), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n498), .B(KEYINPUT101), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n293), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n637), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n293), .A2(new_n499), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n376), .A2(new_n635), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n662));
  INV_X1    g476(.A(new_n569), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n621), .A2(new_n274), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n623), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n621), .A2(KEYINPUT25), .A3(new_n274), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n626), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n619), .B(KEYINPUT102), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n617), .A2(KEYINPUT36), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n662), .B1(new_n667), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n619), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n626), .B1(new_n672), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n625), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n660), .A2(new_n661), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT104), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT37), .B(G110), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  NAND2_X1  g500(.A1(new_n370), .A2(new_n338), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n359), .A2(new_n332), .A3(new_n339), .A4(new_n342), .ZN(new_n688));
  AOI21_X1  g502(.A(G902), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n366), .B1(new_n689), .B2(new_n364), .ZN(new_n690));
  INV_X1    g504(.A(new_n375), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n297), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n625), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT103), .B1(new_n625), .B2(new_n680), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n692), .B(new_n568), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n493), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n696), .B1(new_n697), .B2(new_n495), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n652), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n695), .A2(new_n293), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n258), .ZN(G30));
  XNOR2_X1  g516(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n698), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n692), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT40), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n272), .A2(new_n290), .ZN(new_n707));
  INV_X1    g521(.A(new_n273), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n272), .A2(new_n290), .A3(new_n273), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT38), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n552), .A2(new_n559), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n531), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n714), .B2(G902), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n548), .A2(new_n567), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n187), .ZN(new_n717));
  INV_X1    g531(.A(new_n489), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n638), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n682), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n706), .A2(new_n712), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G143), .ZN(G45));
  AOI21_X1  g536(.A(new_n566), .B1(new_n535), .B2(new_n545), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n540), .A2(new_n543), .A3(new_n536), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT29), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n554), .B(new_n274), .C1(new_n726), .C2(new_n561), .ZN(new_n727));
  AOI22_X1  g541(.A1(KEYINPUT32), .A2(new_n723), .B1(new_n727), .B2(G472), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n676), .A2(new_n681), .B1(new_n728), .B2(new_n567), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n717), .B1(new_n709), .B2(new_n710), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n428), .A2(new_n435), .A3(new_n432), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n435), .B1(new_n428), .B2(new_n432), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n644), .B(new_n699), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n692), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(G146), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G48));
  AOI21_X1  g551(.A(new_n636), .B1(new_n728), .B2(new_n567), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n363), .A2(new_n274), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n298), .A3(new_n365), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n646), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  AND3_X1   g558(.A1(new_n741), .A2(new_n568), .A3(new_n628), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n656), .A3(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n741), .A2(new_n568), .A3(new_n628), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n711), .A2(new_n187), .A3(new_n652), .A4(new_n654), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G116), .ZN(G18));
  NAND4_X1  g566(.A1(new_n660), .A2(new_n682), .A3(new_n568), .A4(new_n741), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  OR2_X1    g568(.A1(new_n553), .A2(new_n536), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n535), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n547), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n633), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n655), .B(new_n489), .C1(new_n434), .C2(new_n436), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n628), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n730), .A2(new_n741), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n633), .A3(new_n625), .A4(new_n627), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n638), .A2(new_n718), .A3(new_n654), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n740), .A2(new_n298), .A3(new_n365), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n293), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G122), .ZN(G24));
  OAI21_X1  g585(.A(new_n758), .B1(new_n693), .B2(new_n694), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n733), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n638), .A2(KEYINPUT109), .A3(new_n644), .A4(new_n699), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n772), .A2(new_n776), .A3(new_n761), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n392), .ZN(G27));
  NAND3_X1  g592(.A1(new_n634), .A2(KEYINPUT111), .A3(new_n564), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n567), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n728), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n628), .A3(new_n774), .A4(new_n775), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n709), .A2(new_n187), .A3(new_n710), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT110), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n709), .A2(new_n786), .A3(new_n187), .A4(new_n710), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n692), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT42), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n291), .A2(new_n292), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n786), .B1(new_n790), .B2(new_n187), .ZN(new_n791));
  INV_X1    g605(.A(new_n787), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n774), .A2(new_n775), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n738), .A3(new_n795), .A4(new_n692), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n317), .ZN(G33));
  AND3_X1   g612(.A1(new_n785), .A2(new_n692), .A3(new_n787), .ZN(new_n799));
  INV_X1    g613(.A(new_n700), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n738), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND2_X1  g616(.A1(new_n372), .A2(new_n374), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT45), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(KEYINPUT45), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n804), .A2(new_n805), .A3(new_n364), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n366), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT46), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n806), .B2(new_n366), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n365), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n298), .A3(new_n704), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n785), .A2(new_n787), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n434), .A2(new_n436), .A3(new_n644), .ZN(new_n815));
  NAND2_X1  g629(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n682), .A3(new_n635), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n813), .B(new_n822), .C1(new_n821), .C2(new_n820), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NAND2_X1  g638(.A1(new_n811), .A2(new_n298), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT47), .Z(new_n826));
  NOR4_X1   g640(.A1(new_n814), .A2(new_n568), .A3(new_n628), .A4(new_n733), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NOR4_X1   g643(.A1(new_n636), .A2(new_n815), .A3(new_n297), .A4(new_n717), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT113), .Z(new_n831));
  NAND2_X1  g645(.A1(new_n740), .A2(new_n365), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT49), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n831), .A2(new_n712), .A3(new_n716), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT114), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n832), .A2(new_n298), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n819), .A2(new_n696), .ZN(new_n838));
  INV_X1    g652(.A(new_n763), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n793), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT116), .Z(new_n841));
  NOR2_X1   g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n843), .A2(new_n187), .A3(new_n712), .A4(new_n766), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT50), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n814), .A2(new_n766), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n716), .A2(new_n636), .A3(new_n493), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n848), .A2(new_n638), .A3(new_n644), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n838), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n845), .B(new_n849), .C1(new_n772), .C2(new_n850), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n481), .A2(new_n482), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n699), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n695), .A2(new_n651), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n772), .A2(new_n776), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n858), .A2(new_n793), .B1(new_n859), .B2(new_n799), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n789), .A3(new_n796), .A4(new_n801), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n638), .A2(new_n856), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n730), .A2(new_n862), .A3(new_n863), .A4(new_n654), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n692), .A2(new_n628), .A3(new_n634), .A4(new_n633), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n730), .A2(new_n654), .A3(new_n862), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(KEYINPUT115), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n864), .A2(new_n867), .B1(new_n746), .B2(new_n750), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n738), .A2(KEYINPUT78), .ZN(new_n869));
  INV_X1    g683(.A(new_n630), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n500), .B1(new_n762), .B2(new_n769), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n638), .A2(new_n644), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n293), .A2(new_n873), .A3(new_n655), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n637), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n683), .A2(new_n753), .A3(new_n875), .A4(new_n742), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n868), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n861), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n701), .A2(new_n777), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n293), .A2(new_n719), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n667), .A2(new_n675), .A3(new_n698), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n692), .A3(new_n716), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n879), .A2(new_n880), .A3(new_n735), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n695), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n730), .A3(new_n800), .ZN(new_n886));
  INV_X1    g700(.A(new_n776), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n682), .A3(new_n767), .A4(new_n758), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n888), .A3(new_n735), .A4(new_n883), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n878), .A2(KEYINPUT53), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n866), .A2(KEYINPUT115), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n637), .A3(new_n864), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT107), .B1(new_n745), .B2(new_n656), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n748), .A2(new_n749), .A3(new_n747), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n760), .A2(new_n761), .A3(KEYINPUT108), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n768), .B1(new_n765), .B2(new_n767), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n631), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n753), .A2(new_n875), .A3(new_n742), .A4(new_n683), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n859), .A2(new_n799), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n857), .A2(new_n651), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n885), .A2(new_n793), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n801), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n797), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n901), .A2(new_n906), .A3(new_n884), .A4(new_n890), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n891), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT54), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n628), .A2(new_n846), .A3(new_n782), .A4(new_n838), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT48), .ZN(new_n913));
  OAI221_X1 g727(.A(new_n491), .B1(new_n843), .B2(new_n761), .C1(new_n848), .C2(new_n873), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n854), .A2(new_n855), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n835), .B1(new_n916), .B2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n334), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n910), .A2(G902), .ZN(new_n921));
  INV_X1    g735(.A(G210), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n271), .A2(new_n270), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n237), .B2(new_n240), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n266), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n919), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n921), .B(KEYINPUT117), .Z(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n708), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n920), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT118), .B(new_n929), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT118), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n930), .B2(new_n708), .ZN(new_n935));
  INV_X1    g749(.A(new_n929), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n937), .ZN(G51));
  NAND2_X1  g752(.A1(new_n930), .A2(new_n806), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n366), .B(KEYINPUT57), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n911), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n363), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n919), .B1(new_n939), .B2(new_n942), .ZN(G54));
  NAND3_X1  g757(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n411), .A3(new_n418), .ZN(new_n945));
  INV_X1    g759(.A(new_n919), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .A4(new_n419), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G60));
  NAND2_X1  g762(.A1(new_n639), .A2(new_n640), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n642), .B(KEYINPUT59), .Z(new_n950));
  NAND3_X1  g764(.A1(new_n911), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT119), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n946), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n951), .B2(new_n946), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n949), .B1(new_n911), .B2(new_n950), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G63));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n957));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT120), .Z(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT60), .Z(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n910), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  AOI211_X1 g776(.A(KEYINPUT121), .B(new_n962), .C1(new_n891), .C2(new_n909), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n621), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n919), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n672), .A2(new_n679), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n961), .B2(new_n963), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(KEYINPUT122), .B(new_n968), .C1(new_n961), .C2(new_n963), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g787(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n973), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G66));
  OAI21_X1  g792(.A(G953), .B1(new_n496), .B2(new_n263), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n877), .B(KEYINPUT124), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n981), .B2(G953), .ZN(new_n982));
  INV_X1    g796(.A(G898), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n925), .B1(new_n983), .B2(G953), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT125), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n982), .B(new_n985), .ZN(G69));
  NAND2_X1  g800(.A1(new_n517), .A2(new_n523), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(new_n414), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n697), .B2(new_n334), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n828), .A2(new_n789), .A3(new_n796), .A4(new_n801), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n813), .A2(new_n628), .A3(new_n782), .A4(new_n881), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n879), .A2(new_n735), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n823), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n989), .B1(new_n994), .B2(new_n334), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n862), .B1(new_n638), .B2(new_n644), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n814), .A2(new_n996), .A3(new_n705), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n997), .A2(new_n871), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT126), .Z(new_n999));
  NAND3_X1  g813(.A1(new_n828), .A2(new_n823), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n992), .A2(new_n721), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(KEYINPUT62), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(KEYINPUT62), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n334), .ZN(new_n1004));
  INV_X1    g818(.A(new_n988), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n334), .B1(G227), .B2(G900), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n1005), .B2(KEYINPUT127), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(G72));
  NAND2_X1  g823(.A1(new_n524), .A2(new_n526), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n530), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1003), .A2(new_n980), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  AOI21_X1  g828(.A(new_n1011), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1014), .ZN(new_n1016));
  INV_X1    g830(.A(new_n561), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n531), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n910), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n994), .B2(new_n981), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1010), .A2(new_n530), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n946), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1015), .A2(new_n1019), .A3(new_n1022), .ZN(G57));
endmodule


