//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n212, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1168, new_n1169, new_n1171,
    new_n1172, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G87), .ZN(G355));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n203), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n217), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n206), .A2(new_n207), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n215), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n220), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT65), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n257), .B2(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G33), .A3(G41), .ZN(new_n269));
  INV_X1    g0069(.A(new_n232), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n271), .A2(new_n263), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n265), .B1(new_n272), .B2(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G190), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT74), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n232), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n208), .A2(G20), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT8), .B(G58), .Z(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n284), .A2(new_n286), .B1(G150), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n282), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n214), .A2(G20), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT67), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n282), .A2(new_n278), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n279), .B(new_n289), .C1(G50), .C2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n274), .A2(G200), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n277), .A2(new_n298), .A3(KEYINPUT10), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT10), .B1(new_n298), .B2(new_n277), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n275), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT68), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n294), .B1(new_n304), .B2(new_n274), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n299), .A2(new_n300), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n293), .A2(G77), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G77), .B2(new_n278), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n284), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n282), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT69), .B(G107), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n317), .B1(new_n319), .B2(new_n254), .C1(new_n258), .C2(new_n222), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n261), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n265), .B1(new_n272), .B2(G244), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(KEYINPUT70), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n323), .B2(G200), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n308), .A2(new_n315), .ZN(new_n330));
  AOI21_X1  g0130(.A(G169), .B1(new_n321), .B2(new_n322), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT72), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n321), .A2(new_n301), .A3(new_n322), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n238), .A2(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(G226), .B2(G1698), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n340), .A2(new_n343), .B1(new_n285), .B2(new_n210), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n265), .B1(new_n344), .B2(new_n261), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n272), .A2(G238), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G169), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n347), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n354), .A2(new_n348), .A3(G179), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n350), .A2(new_n357), .A3(G169), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n293), .A2(G68), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT77), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  INV_X1    g0162(.A(new_n287), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n207), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n287), .A2(KEYINPUT76), .A3(G50), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n286), .A2(G77), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n203), .A2(G20), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n368), .A2(new_n281), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n369), .A2(KEYINPUT11), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(KEYINPUT11), .ZN(new_n371));
  INV_X1    g0171(.A(new_n278), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n203), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n361), .A2(new_n370), .A3(new_n371), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n359), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(G200), .B2(new_n350), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n354), .A2(new_n355), .A3(new_n348), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n324), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n306), .A2(new_n338), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n204), .A2(new_n205), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n287), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n384), .B2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n341), .A2(new_n342), .A3(G20), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT78), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n254), .C2(G20), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n392), .A2(new_n395), .B1(KEYINPUT7), .B2(new_n391), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n390), .B(KEYINPUT16), .C1(new_n203), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n384), .A2(G20), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n386), .A3(new_n387), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n391), .A2(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n394), .B1(new_n254), .B2(G20), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n203), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n398), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n405), .A3(new_n281), .ZN(new_n406));
  INV_X1    g0206(.A(new_n284), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n278), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n293), .B2(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n259), .A2(new_n255), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n410), .B1(G226), .B2(new_n255), .C1(new_n341), .C2(new_n342), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT81), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n261), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n272), .A2(G232), .ZN(new_n416));
  INV_X1    g0216(.A(new_n265), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n415), .A2(new_n324), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(G200), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n406), .A2(new_n409), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(KEYINPUT17), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n406), .A2(new_n409), .A3(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT82), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT82), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n406), .A2(new_n420), .A3(new_n425), .A4(new_n409), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n427), .B2(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n419), .A2(G179), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G169), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n406), .A2(new_n409), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n382), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n254), .A2(G250), .A3(new_n255), .ZN(new_n437));
  OAI211_X1 g0237(.A(G257), .B(G1698), .C1(new_n341), .C2(new_n342), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G294), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n261), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT5), .B(G41), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n271), .A2(G274), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n443), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n271), .A3(G264), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G200), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT88), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n441), .A2(new_n447), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(KEYINPUT87), .A3(new_n324), .A4(new_n445), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT87), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n448), .B2(G190), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n448), .A2(KEYINPUT88), .A3(new_n449), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n452), .A2(new_n454), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n254), .A2(G87), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n215), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n215), .B1(new_n318), .B2(KEYINPUT23), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n254), .A2(KEYINPUT22), .A3(G87), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT24), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n459), .A2(new_n460), .B1(G20), .B2(new_n462), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n465), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n282), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT25), .B1(new_n372), .B2(new_n211), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n214), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n278), .A2(new_n478), .A3(new_n232), .A4(new_n280), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n476), .A2(new_n477), .B1(new_n211), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n458), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n446), .A2(new_n271), .A3(G257), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n445), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT85), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT85), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n445), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n261), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n255), .C1(new_n341), .C2(new_n342), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT84), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n254), .A2(new_n499), .A3(G250), .A4(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n489), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n488), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n487), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n486), .B1(new_n483), .B2(new_n445), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n498), .A2(new_n500), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n261), .B1(new_n507), .B2(new_n495), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n508), .A3(G179), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g0310(.A1(KEYINPUT83), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(KEYINPUT83), .A2(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT6), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G107), .ZN(new_n515));
  XNOR2_X1  g0315(.A(G97), .B(G107), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n513), .A2(new_n515), .B1(new_n516), .B2(new_n514), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n517), .A2(new_n215), .B1(new_n257), .B2(new_n363), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n319), .B1(new_n402), .B2(new_n403), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n281), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n278), .A2(G97), .ZN(new_n521));
  INV_X1    g0321(.A(new_n479), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n488), .A2(new_n502), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G190), .ZN(new_n527));
  INV_X1    g0327(.A(new_n524), .ZN(new_n528));
  OAI21_X1  g0328(.A(G200), .B1(new_n488), .B2(new_n502), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n254), .A2(G238), .A3(new_n255), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n254), .A2(G244), .A3(G1698), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n261), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n443), .A2(new_n224), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n271), .A2(new_n536), .B1(G274), .B2(new_n443), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n513), .A2(new_n286), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n254), .A2(new_n215), .A3(G68), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n513), .A2(new_n318), .A3(G87), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n285), .A2(new_n210), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(new_n545), .B2(KEYINPUT19), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n281), .B1(new_n372), .B2(new_n309), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n522), .A2(G87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n535), .A2(G190), .A3(new_n537), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n539), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n543), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n318), .A2(G87), .ZN(new_n553));
  INV_X1    g0353(.A(new_n513), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n546), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n281), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n309), .A2(new_n372), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n522), .A2(new_n310), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n538), .A2(new_n304), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n535), .A2(new_n301), .A3(new_n537), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n551), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n482), .A2(new_n525), .A3(new_n530), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n522), .A2(KEYINPUT86), .A3(G116), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  INV_X1    g0366(.A(G116), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n479), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(G20), .ZN(new_n570));
  INV_X1    g0370(.A(G13), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n570), .A2(G1), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(G33), .B1(new_n511), .B2(new_n512), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n494), .A2(new_n215), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n281), .A2(new_n570), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT20), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(KEYINPUT20), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n569), .B(new_n573), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n254), .A2(G257), .A3(new_n255), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n343), .A2(G303), .ZN(new_n583));
  INV_X1    g0383(.A(G264), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n258), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n261), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n446), .A2(new_n271), .A3(G270), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n445), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n304), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n588), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n301), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n590), .A2(new_n591), .B1(new_n593), .B2(new_n581), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n453), .A2(new_n301), .A3(new_n445), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n448), .A2(new_n304), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n474), .C2(new_n480), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n581), .A2(new_n589), .A3(KEYINPUT21), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n578), .A2(new_n580), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n572), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n592), .A2(G200), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n586), .A2(new_n588), .A3(G190), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n569), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n594), .A2(new_n597), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n436), .A2(new_n564), .A3(new_n604), .ZN(G372));
  INV_X1    g0405(.A(new_n336), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n379), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n376), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n428), .ZN(new_n609));
  INV_X1    g0409(.A(new_n433), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n299), .A2(new_n300), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(new_n303), .B2(new_n305), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT89), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n564), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n506), .A2(new_n508), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n524), .B1(new_n616), .B2(G200), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n527), .A2(new_n617), .B1(new_n510), .B2(new_n524), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT89), .A3(new_n482), .A4(new_n563), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n528), .B1(new_n510), .B2(KEYINPUT90), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT90), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n503), .A2(new_n509), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n563), .A4(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n528), .B1(new_n503), .B2(new_n509), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n563), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n626), .A2(new_n629), .A3(new_n562), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n613), .B1(new_n436), .B2(new_n632), .ZN(G369));
  INV_X1    g0433(.A(new_n603), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n594), .A2(new_n598), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n571), .A2(G20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n214), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT91), .Z(new_n638));
  INV_X1    g0438(.A(KEYINPUT27), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(G213), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n581), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n635), .A2(new_n645), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n634), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(KEYINPUT92), .B(G330), .Z(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n644), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n482), .B1(new_n481), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n597), .ZN(new_n654));
  INV_X1    g0454(.A(new_n597), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n644), .B1(new_n594), .B2(new_n598), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n655), .B2(new_n652), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n218), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G1), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n544), .A2(new_n567), .ZN(new_n668));
  INV_X1    g0468(.A(new_n231), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n667), .A2(new_n668), .B1(new_n669), .B2(new_n666), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n525), .A2(new_n530), .A3(new_n563), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n482), .A3(new_n620), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n622), .A2(new_n563), .A3(new_n625), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT26), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n563), .A2(new_n627), .A3(new_n623), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n562), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(KEYINPUT29), .A3(new_n652), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n632), .A2(new_n644), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(KEYINPUT29), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n564), .A2(new_n604), .A3(new_n644), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n441), .A2(new_n447), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n592), .A2(new_n538), .A3(new_n682), .A4(new_n301), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n526), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n526), .ZN(new_n687));
  AOI21_X1  g0487(.A(G179), .B1(new_n535), .B2(new_n537), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n616), .A2(new_n448), .A3(new_n592), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(new_n644), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT31), .B1(new_n681), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n644), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n649), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n680), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n671), .B1(new_n698), .B2(G1), .ZN(G364));
  AOI21_X1  g0499(.A(new_n214), .B1(new_n636), .B2(G45), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n665), .A2(KEYINPUT93), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT93), .B1(new_n665), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n648), .B2(new_n650), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n650), .B2(new_n648), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT94), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT32), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G179), .A2(G200), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(G20), .A3(new_n324), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT99), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT99), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G159), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n215), .A2(new_n301), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT97), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n449), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G190), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n711), .A2(new_n718), .B1(new_n723), .B2(G77), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n722), .A2(new_n324), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n719), .A2(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n324), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT98), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n729), .A2(KEYINPUT98), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n724), .B1(new_n202), .B2(new_n726), .C1(new_n734), .C2(new_n207), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n727), .A2(G190), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n215), .B1(new_n712), .B2(G190), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n736), .A2(G68), .B1(G97), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT100), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n215), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n223), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(new_n324), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n343), .B(new_n743), .C1(G107), .C2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n740), .B(new_n746), .C1(new_n711), .C2(new_n718), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n725), .A2(G322), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  INV_X1    g0549(.A(new_n723), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n748), .B1(new_n749), .B2(new_n750), .C1(new_n734), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n716), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G329), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n736), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n742), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G303), .B1(new_n745), .B2(G283), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n254), .B1(new_n738), .B2(G294), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n754), .A2(new_n758), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n735), .A2(new_n747), .B1(new_n752), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n232), .B1(G20), .B2(new_n304), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n704), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n764), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n664), .A2(new_n343), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G355), .B1(new_n567), .B2(new_n664), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n252), .A2(G45), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n664), .A2(new_n254), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n669), .B2(G45), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT96), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n769), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n776), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(new_n768), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n765), .B1(new_n778), .B2(new_n780), .C1(new_n648), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n709), .A2(new_n710), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT101), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  NAND2_X1  g0585(.A1(new_n644), .A2(new_n316), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n329), .A2(new_n336), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT103), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n329), .A2(new_n336), .A3(new_n789), .A4(new_n786), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n336), .A2(new_n786), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n679), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n705), .B1(new_n793), .B2(new_n697), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n697), .B2(new_n793), .ZN(new_n795));
  INV_X1    g0595(.A(new_n764), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G143), .A2(new_n725), .B1(new_n723), .B2(G159), .ZN(new_n797));
  INV_X1    g0597(.A(G150), .ZN(new_n798));
  INV_X1    g0598(.A(new_n736), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n797), .B1(new_n798), .B2(new_n799), .C1(new_n734), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n254), .B1(new_n742), .B2(new_n207), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n744), .A2(new_n203), .B1(new_n737), .B2(new_n202), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(new_n753), .C2(G132), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n343), .B1(new_n737), .B2(new_n210), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n799), .A2(new_n808), .B1(new_n211), .B2(new_n742), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n733), .C2(G303), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n716), .A2(new_n749), .B1(new_n223), .B2(new_n744), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT102), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G116), .A2(new_n723), .B1(new_n725), .B2(G294), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n796), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n764), .A2(new_n766), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n704), .B(new_n815), .C1(new_n257), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n792), .B2(new_n767), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n795), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  INV_X1    g0620(.A(new_n517), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n822), .A2(new_n823), .A3(G116), .A4(new_n233), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT36), .Z(new_n825));
  NAND3_X1  g0625(.A1(new_n231), .A2(G77), .A3(new_n383), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n207), .A2(G68), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n214), .B(G13), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n631), .A2(new_n792), .A3(new_n652), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n336), .A2(new_n644), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n375), .A2(new_n644), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n376), .A2(new_n379), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n359), .A2(new_n375), .A3(new_n644), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT104), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n642), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n390), .B1(new_n396), .B2(new_n203), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n842), .A2(new_n398), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n397), .A2(new_n281), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n409), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n434), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n427), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n429), .A2(new_n431), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n848), .B2(new_n841), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n406), .A2(new_n409), .ZN(new_n852));
  AOI211_X1 g0652(.A(KEYINPUT37), .B(new_n432), .C1(new_n852), .C2(new_n841), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n847), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n846), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n833), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n840), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n610), .A2(new_n642), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n376), .A2(new_n644), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  XOR2_X1   g0665(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n866));
  INV_X1    g0666(.A(KEYINPUT106), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n421), .B2(new_n432), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n852), .A2(new_n848), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT106), .A3(new_n423), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n852), .A2(new_n841), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT107), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n854), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n642), .B1(new_n428), .B2(new_n433), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n852), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n866), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n846), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n865), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n858), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n863), .B1(new_n864), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n435), .B(new_n678), .C1(KEYINPUT29), .C2(new_n679), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n613), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n885), .B(new_n887), .Z(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT108), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n880), .B2(new_n881), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n873), .A2(new_n874), .B1(new_n847), .B2(new_n853), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(new_n876), .B1(new_n852), .B2(new_n878), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT108), .B(new_n858), .C1(new_n893), .C2(new_n866), .ZN(new_n894));
  AND4_X1   g0694(.A1(new_n598), .A2(new_n594), .A3(new_n597), .A4(new_n603), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n672), .A2(new_n895), .A3(new_n482), .A4(new_n652), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n694), .B1(new_n896), .B2(new_n693), .ZN(new_n897));
  INV_X1    g0697(.A(new_n695), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n837), .B(new_n792), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n891), .A2(new_n894), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n899), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n881), .B2(new_n856), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n692), .A2(new_n695), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n435), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n906), .A2(new_n908), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n910), .A2(new_n911), .A3(new_n649), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n889), .A2(new_n912), .B1(new_n214), .B2(new_n636), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n889), .A2(new_n912), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n829), .B1(new_n913), .B2(new_n914), .ZN(G367));
  OAI21_X1  g0715(.A(new_n618), .B1(new_n528), .B2(new_n652), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n622), .A2(new_n625), .A3(new_n644), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n661), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT42), .Z(new_n920));
  AOI21_X1  g0720(.A(new_n597), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n652), .B1(new_n921), .B2(new_n627), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n548), .A2(new_n549), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n644), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n563), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n562), .B2(new_n924), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n920), .A2(new_n922), .B1(KEYINPUT43), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n658), .A2(new_n918), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n929), .B(new_n930), .Z(new_n931));
  XOR2_X1   g0731(.A(new_n665), .B(KEYINPUT41), .Z(new_n932));
  NAND2_X1  g0732(.A1(new_n662), .A2(new_n918), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT109), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT109), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n662), .A2(new_n935), .A3(new_n918), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n662), .A2(new_n918), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT44), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n658), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n939), .A2(new_n941), .A3(new_n659), .A4(new_n942), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n657), .B(new_n660), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n651), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n944), .A2(new_n698), .A3(new_n945), .A4(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n932), .B1(new_n948), .B2(new_n698), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n931), .B1(new_n701), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n774), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n769), .B1(new_n218), .B2(new_n309), .C1(new_n951), .C2(new_n244), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(KEYINPUT110), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(KEYINPUT110), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n953), .A2(new_n954), .A3(new_n704), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n726), .A2(new_n798), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n744), .A2(new_n257), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n343), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT112), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n734), .B2(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n750), .A2(new_n207), .B1(KEYINPUT112), .B2(new_n958), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n759), .A2(G58), .B1(new_n738), .B2(G68), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n799), .B2(new_n717), .C1(new_n800), .C2(new_n716), .ZN(new_n964));
  OR4_X1    g0764(.A1(new_n956), .A2(new_n961), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n733), .A2(G311), .B1(G283), .B2(new_n723), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n742), .A2(new_n567), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT111), .B(G317), .Z(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n753), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n343), .B1(new_n554), .B2(new_n744), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n736), .A2(G294), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n319), .B2(new_n737), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(G303), .C2(new_n725), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n966), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n965), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n955), .B1(new_n781), .B2(new_n926), .C1(new_n978), .C2(new_n796), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n950), .A2(new_n979), .ZN(G387));
  XNOR2_X1  g0780(.A(new_n665), .B(KEYINPUT117), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n698), .B2(new_n947), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n698), .B2(new_n947), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n241), .A2(new_n442), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n985), .A2(new_n774), .B1(new_n668), .B2(new_n770), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n407), .A2(G50), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT50), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n442), .B1(new_n203), .B2(new_n257), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n668), .B(new_n989), .C1(new_n988), .C2(new_n987), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n986), .A2(new_n990), .B1(G107), .B2(new_n218), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n704), .B1(new_n991), .B2(new_n769), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n733), .A2(G159), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT115), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n742), .A2(new_n257), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n343), .B(new_n995), .C1(G97), .C2(new_n745), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n798), .B2(new_n716), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT114), .Z(new_n998));
  AOI22_X1  g0798(.A1(new_n736), .A2(new_n284), .B1(new_n310), .B2(new_n738), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n750), .B2(new_n203), .C1(new_n207), .C2(new_n726), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n994), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n759), .A2(G294), .B1(new_n738), .B2(G283), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G303), .A2(new_n723), .B1(new_n725), .B2(new_n969), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT116), .B(G322), .Z(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n749), .B2(new_n799), .C1(new_n734), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT48), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n343), .B1(new_n567), .B2(new_n744), .C1(new_n716), .C2(new_n751), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n1008), .B2(KEYINPUT49), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1001), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n992), .B1(new_n1012), .B2(new_n796), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n657), .B2(new_n768), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n947), .B2(new_n701), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n984), .A2(new_n1015), .ZN(G393));
  NAND2_X1  g0816(.A1(new_n944), .A2(new_n945), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n698), .A2(new_n947), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n948), .A3(new_n981), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n944), .A2(new_n701), .A3(new_n945), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n769), .B1(new_n218), .B2(new_n554), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n249), .B2(new_n774), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n704), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n733), .A2(G317), .B1(G311), .B2(new_n725), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n736), .A2(G303), .B1(G116), .B2(new_n738), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n808), .B2(new_n742), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n343), .B1(new_n211), .B2(new_n744), .C1(new_n716), .C2(new_n1004), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G294), .C2(new_n723), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n733), .A2(G150), .B1(G159), .B2(new_n725), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT51), .Z(new_n1032));
  AOI22_X1  g0832(.A1(new_n736), .A2(G50), .B1(G77), .B2(new_n738), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n203), .B2(new_n742), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n254), .B1(new_n223), .B2(new_n744), .C1(new_n716), .C2(new_n960), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n284), .C2(new_n723), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1026), .A2(new_n1030), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1024), .B1(new_n918), .B2(new_n781), .C1(new_n1037), .C2(new_n796), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1021), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1020), .A2(new_n1039), .ZN(G390));
  OAI211_X1 g0840(.A(G330), .B(new_n792), .C1(new_n897), .C2(new_n898), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n837), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n792), .A2(new_n677), .A3(new_n652), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n832), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n864), .B1(new_n1045), .B2(new_n837), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n891), .A2(new_n894), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n864), .B1(new_n833), .B2(new_n837), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n882), .B2(new_n883), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1043), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT118), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n1043), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n891), .A2(new_n894), .A3(new_n1046), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n696), .A2(new_n792), .A3(new_n837), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n884), .C2(new_n1048), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(G330), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n886), .B(new_n613), .C1(new_n1058), .C2(new_n908), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n837), .B1(new_n696), .B2(new_n792), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n833), .B1(new_n1060), .B2(new_n1043), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT119), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(KEYINPUT119), .B(new_n833), .C1(new_n1060), .C2(new_n1043), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1055), .A2(new_n1066), .A3(new_n832), .A4(new_n1044), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1059), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1057), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1051), .A2(new_n1053), .A3(new_n1068), .A4(new_n1056), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n981), .A3(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1051), .A2(new_n701), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n733), .A2(G128), .B1(G132), .B2(new_n725), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n742), .A2(new_n798), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(KEYINPUT54), .B(G143), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1074), .B(new_n1077), .C1(new_n750), .C2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n736), .A2(G137), .B1(new_n745), .B2(G50), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n343), .B1(new_n738), .B2(G159), .ZN(new_n1081));
  INV_X1    g0881(.A(G125), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1081), .C1(new_n1082), .C2(new_n716), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n733), .A2(G283), .B1(G116), .B2(new_n725), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n554), .B2(new_n750), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n254), .B(new_n743), .C1(new_n753), .C2(G294), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n745), .A2(G68), .B1(new_n738), .B2(G77), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n319), .C2(new_n799), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1079), .A2(new_n1083), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n764), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n704), .B1(new_n407), .B2(new_n816), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n884), .C2(new_n767), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1072), .A2(new_n1073), .A3(new_n1092), .ZN(G378));
  INV_X1    g0893(.A(new_n885), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1058), .B1(new_n904), .B2(new_n900), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n902), .A2(new_n1095), .A3(KEYINPUT122), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT122), .B1(new_n902), .B2(new_n1095), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n294), .A2(new_n642), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n306), .B(new_n1099), .Z(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1097), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1102), .A2(new_n902), .A3(new_n1095), .A4(KEYINPUT122), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1094), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n902), .A2(new_n1095), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1102), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1096), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n885), .A3(new_n1104), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n701), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n704), .B1(new_n207), .B2(new_n816), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n750), .A2(new_n800), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n736), .A2(G132), .B1(G150), .B2(new_n738), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n742), .B2(new_n1078), .C1(new_n734), .C2(new_n1082), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G128), .C2(new_n725), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n753), .A2(G124), .ZN(new_n1122));
  AOI211_X1 g0922(.A(G33), .B(G41), .C1(new_n745), .C2(G159), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n211), .A2(new_n726), .B1(new_n750), .B2(new_n309), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n744), .A2(new_n202), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n995), .B(new_n1126), .C1(G97), .C2(new_n736), .ZN(new_n1127));
  AOI211_X1 g0927(.A(G41), .B(new_n254), .C1(new_n738), .C2(G68), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n808), .C2(new_n716), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1125), .B(new_n1129), .C1(G116), .C2(new_n733), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT58), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(KEYINPUT58), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n207), .B1(new_n341), .B2(G41), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n1124), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1114), .B1(new_n796), .B2(new_n1134), .C1(new_n1110), .C2(new_n767), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT121), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1113), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1059), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1071), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1139), .A2(KEYINPUT57), .A3(new_n1106), .A4(new_n1112), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n981), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1111), .A2(new_n885), .A3(new_n1104), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n885), .B1(new_n1111), .B2(new_n1104), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT57), .B1(new_n1144), .B2(new_n1139), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1137), .B1(new_n1141), .B2(new_n1145), .ZN(G375));
  INV_X1    g0946(.A(new_n932), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1065), .A2(new_n1059), .A3(new_n1067), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1069), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n254), .B(new_n957), .C1(new_n753), .C2(G303), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n759), .A2(G97), .B1(new_n738), .B2(new_n310), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n567), .C2(new_n799), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n733), .A2(G294), .B1(G283), .B2(new_n725), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n319), .B2(new_n750), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n733), .A2(G132), .B1(G137), .B2(new_n725), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n798), .B2(new_n750), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n343), .B(new_n1126), .C1(new_n753), .C2(G128), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n759), .A2(G159), .B1(new_n738), .B2(G50), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n799), .C2(new_n1078), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1152), .A2(new_n1154), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n764), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n704), .B1(new_n203), .B2(new_n816), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1042), .B2(new_n766), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n701), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1149), .A2(new_n1166), .ZN(G381));
  NAND3_X1  g0967(.A1(new_n984), .A2(new_n784), .A3(new_n1015), .ZN(new_n1168));
  OR4_X1    g0968(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1168), .ZN(new_n1169));
  OR4_X1    g0969(.A1(G378), .A2(new_n1169), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g0970(.A1(new_n643), .A2(G213), .ZN(new_n1171));
  OR3_X1    g0971(.A1(G375), .A2(G378), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(G407), .A2(G213), .A3(new_n1172), .ZN(G409));
  INV_X1    g0973(.A(new_n1168), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n784), .B1(new_n984), .B2(new_n1015), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(G390), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1020), .B(new_n1039), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(G387), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n950), .A4(new_n979), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT61), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G378), .B(new_n1137), .C1(new_n1141), .C2(new_n1145), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1073), .A2(new_n1092), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1072), .A2(new_n1185), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1144), .A2(new_n1147), .A3(new_n1139), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1113), .A2(new_n1136), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1148), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1148), .A2(new_n1191), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n981), .A4(new_n1069), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1166), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n819), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1195), .A2(new_n819), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1190), .A2(new_n1171), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1183), .B1(new_n1201), .B2(KEYINPUT63), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1171), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1198), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(G2897), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT125), .Z(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1196), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1207), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1204), .A2(KEYINPUT124), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(KEYINPUT124), .B2(new_n1204), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT63), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1200), .B2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(KEYINPUT123), .B(KEYINPUT63), .C1(new_n1204), .C2(new_n1199), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1202), .B(new_n1212), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1190), .A2(new_n1171), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1210), .A2(new_n1208), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1204), .A2(KEYINPUT62), .A3(new_n1199), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT62), .B1(new_n1204), .B2(new_n1199), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(KEYINPUT126), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1182), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1200), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1204), .A2(KEYINPUT62), .A3(new_n1199), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT126), .B1(new_n1228), .B2(new_n1220), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1217), .B1(new_n1224), .B2(new_n1229), .ZN(G405));
  INV_X1    g1030(.A(KEYINPUT127), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1199), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(new_n1182), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1199), .A2(new_n1231), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1184), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G375), .B2(new_n1186), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1233), .B(new_n1236), .ZN(G402));
endmodule


