//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  AND2_X1   g000(.A1(KEYINPUT74), .A2(G953), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT74), .A2(G953), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT22), .Z(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT67), .B(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT70), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT70), .A2(G119), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G128), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n195), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n199), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT23), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(G110), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT78), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n207), .B(G110), .C1(new_n201), .C2(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n212), .A2(KEYINPUT79), .A3(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT16), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G125), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(G146), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n211), .B2(new_n213), .ZN(new_n221));
  INV_X1    g035(.A(new_n218), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n197), .A2(new_n200), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT24), .B(G110), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n219), .A2(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n209), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n210), .A2(new_n220), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n224), .A2(new_n226), .ZN(new_n231));
  INV_X1    g045(.A(G110), .ZN(new_n232));
  INV_X1    g046(.A(new_n204), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n232), .B(new_n233), .C1(new_n224), .C2(new_n195), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n201), .A2(G110), .A3(new_n204), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT80), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n230), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n194), .B1(new_n228), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  OAI22_X1  g055(.A1(new_n237), .A2(KEYINPUT80), .B1(new_n224), .B2(new_n226), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n234), .A2(new_n235), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n219), .B(new_n229), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n209), .A2(new_n227), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n193), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT81), .B(KEYINPUT25), .Z(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n240), .A2(new_n246), .A3(new_n241), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G217), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(G234), .B2(new_n241), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT77), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n249), .A2(KEYINPUT82), .A3(new_n251), .A4(new_n254), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n253), .A2(G902), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n240), .A2(KEYINPUT83), .A3(new_n246), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT83), .B1(new_n240), .B2(new_n246), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT66), .B1(new_n264), .B2(G137), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n192), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n264), .B2(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n268), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT72), .B1(new_n270), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n220), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n282), .A2(KEYINPUT1), .A3(new_n203), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(G143), .B2(new_n220), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n196), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT68), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n282), .B(new_n288), .C1(new_n196), .C2(new_n285), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n283), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT73), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT64), .B1(new_n282), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(G143), .B(G146), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT0), .A4(G128), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT0), .B(G128), .Z(new_n297));
  AOI22_X1  g111(.A1(new_n293), .A2(new_n296), .B1(new_n282), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n272), .A2(new_n268), .A3(new_n273), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G131), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(G131), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT65), .A3(new_n275), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n270), .A2(new_n275), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n275), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n310));
  INV_X1    g124(.A(new_n283), .ZN(new_n311));
  INV_X1    g125(.A(new_n289), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT1), .B1(new_n280), .B2(G146), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n288), .B1(new_n317), .B2(new_n282), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n311), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n309), .A2(new_n310), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n291), .A2(new_n304), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT30), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n304), .B(new_n323), .C1(new_n305), .C2(new_n290), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT70), .B(G119), .Z(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G116), .ZN(new_n327));
  OR2_X1    g141(.A1(KEYINPUT71), .A2(G116), .ZN(new_n328));
  NAND2_X1  g142(.A1(KEYINPUT71), .A2(G116), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(G119), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT2), .A2(G113), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT2), .A2(G113), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n327), .A2(new_n333), .A3(new_n334), .A4(new_n330), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n303), .A2(new_n301), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n341), .B2(new_n298), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n291), .A2(new_n342), .A3(new_n320), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n189), .A2(G210), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT27), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT26), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(KEYINPUT26), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n348), .A2(G101), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(G101), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT75), .B(KEYINPUT31), .Z(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n339), .A2(new_n343), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n309), .A2(new_n319), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT28), .B1(new_n342), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n304), .B1(new_n305), .B2(new_n290), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n338), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n343), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n360), .B2(KEYINPUT28), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(new_n352), .ZN(new_n362));
  INV_X1    g176(.A(new_n324), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n321), .B2(KEYINPUT30), .ZN(new_n364));
  INV_X1    g178(.A(new_n338), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n343), .B(new_n352), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT75), .A2(KEYINPUT31), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n355), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n343), .B1(new_n364), .B2(new_n365), .ZN(new_n377));
  INV_X1    g191(.A(new_n352), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n377), .A2(KEYINPUT76), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n361), .A2(new_n352), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT76), .B1(new_n377), .B2(new_n378), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n321), .A2(new_n338), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n343), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n357), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT29), .A3(new_n352), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n241), .ZN(new_n390));
  OAI21_X1  g204(.A(G472), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n263), .B1(new_n376), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n196), .A2(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n280), .A2(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G134), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n264), .B1(new_n393), .B2(new_n394), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n328), .A2(new_n329), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G122), .ZN(new_n399));
  INV_X1    g213(.A(G122), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G116), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n396), .A2(new_n397), .B1(new_n402), .B2(G107), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n404), .A3(new_n401), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(KEYINPUT14), .A3(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G107), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT98), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n405), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n403), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n396), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n402), .A2(G107), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n399), .B2(new_n401), .ZN(new_n418));
  INV_X1    g232(.A(new_n395), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G134), .B1(new_n420), .B2(new_n394), .ZN(new_n422));
  OAI221_X1 g236(.A(new_n415), .B1(new_n416), .B2(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT9), .B(G234), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(new_n252), .A3(G953), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n414), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n425), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n415), .B1(new_n421), .B2(new_n422), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n416), .A2(new_n418), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n427), .B1(new_n430), .B2(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n241), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n241), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(KEYINPUT99), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT99), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n432), .B2(new_n241), .ZN(new_n441));
  AOI211_X1 g255(.A(G902), .B(new_n435), .C1(new_n426), .C2(new_n431), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n445));
  XNOR2_X1  g259(.A(G113), .B(G122), .ZN(new_n446));
  INV_X1    g260(.A(G104), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n214), .B2(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n219), .B1(G146), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n189), .A2(G214), .A3(new_n344), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT95), .B1(KEYINPUT94), .B2(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(KEYINPUT95), .B2(G143), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(new_n189), .A3(G214), .A4(new_n344), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G131), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n274), .A3(new_n457), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n452), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(KEYINPUT18), .A2(G131), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n462), .A3(new_n457), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n229), .B1(new_n214), .B2(new_n220), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n462), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n458), .A2(KEYINPUT96), .A3(new_n466), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n449), .B1(new_n461), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT17), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n459), .A2(new_n474), .A3(new_n460), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n458), .A2(KEYINPUT17), .A3(G131), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n223), .A3(new_n219), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n448), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G475), .A2(G902), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n445), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n445), .A3(new_n480), .ZN(new_n483));
  INV_X1    g297(.A(new_n478), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n448), .B1(new_n473), .B2(new_n477), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n241), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n482), .A2(new_n483), .B1(G475), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G952), .ZN(new_n488));
  AOI211_X1 g302(.A(G953), .B(new_n488), .C1(G234), .C2(G237), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n241), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT21), .B(G898), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n444), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G221), .B1(new_n424), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G110), .B(G140), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n189), .A2(G227), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT3), .B1(new_n447), .B2(G107), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT3), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n417), .A3(G104), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n447), .A2(G107), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(G101), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n447), .A2(KEYINPUT87), .A3(G107), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n447), .B2(G107), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n417), .A2(KEYINPUT86), .A3(G104), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n509), .A2(new_n510), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(G101), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n501), .B1(new_n319), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(G101), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n290), .A2(KEYINPUT88), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n294), .B1(G128), .B2(new_n313), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n283), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT12), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n341), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n506), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT85), .A4(new_n505), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(G101), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT4), .A3(new_n517), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT4), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n530), .A2(new_n534), .A3(G101), .A4(new_n531), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n298), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n319), .A2(KEYINPUT10), .A3(new_n515), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n528), .A2(new_n536), .A3(new_n537), .A4(new_n340), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n526), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n523), .A2(new_n341), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n500), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n536), .A3(new_n537), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n341), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(new_n500), .A3(new_n538), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G469), .B1(new_n547), .B2(G902), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n500), .A3(new_n538), .A4(new_n526), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT90), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n539), .A2(new_n551), .A3(new_n500), .A4(new_n542), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n500), .B1(new_n545), .B2(new_n538), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G469), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n241), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n496), .B1(new_n548), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G210), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G110), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT92), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n515), .A2(new_n337), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n327), .A2(KEYINPUT5), .A3(new_n330), .ZN(new_n567));
  INV_X1    g381(.A(G113), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n198), .A2(G116), .A3(new_n199), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT5), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT91), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n567), .A2(KEYINPUT91), .A3(new_n571), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n338), .A2(new_n535), .A3(new_n533), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n515), .A2(new_n337), .ZN(new_n578));
  INV_X1    g392(.A(new_n574), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n572), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n338), .A2(new_n533), .A3(new_n535), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n564), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n582), .A3(KEYINPUT6), .ZN(new_n583));
  OR3_X1    g397(.A1(new_n298), .A2(KEYINPUT93), .A3(new_n212), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n290), .A2(new_n212), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT93), .B1(new_n298), .B2(new_n212), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G224), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n587), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT6), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n591), .B(new_n565), .C1(new_n575), .C2(new_n576), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n583), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT7), .B1(new_n588), .B2(G953), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n582), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n564), .B(KEYINPUT8), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n566), .B1(new_n567), .B2(new_n571), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n337), .B1(new_n579), .B2(new_n572), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n519), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n241), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n562), .B1(new_n593), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n583), .A2(new_n590), .A3(new_n592), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n561), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n560), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n494), .A2(new_n558), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n392), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  NAND2_X1  g428(.A1(new_n548), .A2(new_n557), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n495), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n263), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n370), .A2(new_n241), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n617), .A2(new_n618), .A3(new_n372), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n263), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n558), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n372), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT100), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n611), .A2(new_n493), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n486), .A2(G475), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n479), .A2(new_n445), .A3(new_n480), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n481), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n433), .A2(new_n434), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n432), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n426), .A2(new_n431), .A3(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n241), .A2(G478), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT101), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n629), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n626), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n621), .A2(new_n625), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT102), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G6));
  NOR3_X1   g459(.A1(new_n626), .A2(new_n444), .A3(new_n629), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n621), .A2(new_n625), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n244), .A2(new_n245), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n259), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n257), .A2(new_n258), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n612), .A2(new_n372), .A3(new_n620), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND3_X1  g471(.A1(new_n391), .A2(new_n374), .A3(new_n375), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n607), .A2(new_n610), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n559), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n616), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT103), .B(G900), .Z(new_n663));
  AOI21_X1  g477(.A(new_n489), .B1(new_n490), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n444), .A2(new_n629), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XOR2_X1   g481(.A(new_n664), .B(KEYINPUT39), .Z(new_n668));
  AND2_X1   g482(.A1(new_n558), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT40), .ZN(new_n670));
  INV_X1    g484(.A(new_n377), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n378), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n291), .A2(new_n320), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n673), .A2(new_n342), .B1(new_n321), .B2(new_n338), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n378), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n241), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n376), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n660), .A2(KEYINPUT104), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n607), .A2(new_n610), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT38), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n679), .A2(KEYINPUT38), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n654), .A2(new_n560), .A3(new_n444), .A4(new_n487), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n670), .A2(new_n678), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT105), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  INV_X1    g504(.A(new_n664), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n629), .A2(new_n636), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n659), .A2(new_n662), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  NAND2_X1  g508(.A1(new_n557), .A2(new_n495), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n555), .A2(new_n241), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n556), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n553), .B1(new_n549), .B2(KEYINPUT90), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n699), .B2(new_n552), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT106), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n695), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n641), .A2(new_n658), .A3(new_n622), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n646), .A2(new_n658), .A3(new_n622), .A4(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  AOI21_X1  g521(.A(new_n496), .B1(new_n700), .B2(new_n556), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n700), .B2(KEYINPUT106), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n697), .B(G902), .C1(new_n699), .C2(new_n552), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n611), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n696), .A2(new_n697), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(G469), .A3(new_n701), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n611), .A4(new_n708), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n659), .A3(new_n494), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NAND2_X1  g533(.A1(new_n263), .A2(KEYINPUT109), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n257), .A2(new_n721), .A3(new_n258), .A4(new_n262), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n661), .A2(new_n444), .A3(new_n487), .A4(new_n492), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT108), .B1(new_n387), .B2(new_n357), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  INV_X1    g540(.A(new_n357), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n726), .B(new_n727), .C1(new_n674), .C2(new_n385), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n725), .A2(new_n378), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n355), .A2(new_n369), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n371), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n620), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n723), .A2(new_n724), .A3(new_n732), .A4(new_n702), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND4_X1  g548(.A1(new_n620), .A2(new_n692), .A3(new_n654), .A4(new_n731), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n717), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n717), .A2(new_n739), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n660), .A2(new_n560), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n744), .A2(new_n615), .A3(new_n495), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n658), .A2(new_n745), .A3(new_n622), .A4(new_n692), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n376), .A2(new_n391), .B1(new_n720), .B2(new_n722), .ZN(new_n747));
  AND4_X1   g561(.A1(KEYINPUT42), .A2(new_n558), .A3(new_n692), .A4(new_n744), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n743), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n274), .ZN(G33));
  NAND4_X1  g564(.A1(new_n487), .A2(new_n443), .A3(new_n439), .A4(new_n691), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n392), .A2(new_n745), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n624), .A2(new_n654), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n624), .A2(KEYINPUT114), .A3(new_n654), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT43), .B1(new_n487), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n487), .A2(new_n636), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n758), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g579(.A(G469), .B1(new_n547), .B2(KEYINPUT45), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT112), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(KEYINPUT112), .B1(KEYINPUT45), .B2(new_n547), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(G469), .A2(G902), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT46), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n557), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n770), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n496), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n765), .A2(new_n668), .A3(new_n744), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  AND2_X1   g591(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n778));
  NOR2_X1   g592(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n692), .A2(new_n744), .A3(new_n263), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n658), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n780), .B(new_n782), .C1(new_n775), .C2(new_n779), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  INV_X1    g598(.A(G953), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n488), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n746), .A2(new_n743), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n747), .A2(new_n748), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n745), .A2(new_n654), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n436), .A2(new_n438), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n629), .A2(new_n791), .A3(new_n664), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n658), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n732), .A2(new_n692), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n789), .A2(new_n796), .A3(new_n754), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n703), .A2(new_n733), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n706), .A3(new_n718), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n487), .A2(new_n791), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n637), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT118), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n626), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n621), .A2(new_n805), .A3(new_n625), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n613), .A3(KEYINPUT53), .A4(new_n655), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n797), .A2(new_n799), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n659), .B(new_n662), .C1(new_n665), .C2(new_n692), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n444), .A2(new_n487), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n611), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n654), .A3(new_n664), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n678), .A3(new_n558), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n739), .B1(new_n717), .B2(new_n736), .ZN(new_n814));
  AOI211_X1 g628(.A(KEYINPUT110), .B(new_n735), .C1(new_n713), .C2(new_n716), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n809), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n741), .A2(KEYINPUT52), .A3(new_n809), .A4(new_n813), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n816), .A2(new_n817), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT120), .A3(new_n808), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT119), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n392), .A2(new_n745), .A3(new_n753), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n749), .A2(new_n830), .A3(new_n795), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n798), .A2(new_n718), .A3(new_n832), .A4(new_n706), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n713), .A2(new_n716), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n658), .A2(new_n494), .A3(new_n654), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n703), .A2(new_n706), .A3(new_n733), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n806), .A2(new_n613), .A3(new_n655), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n831), .A2(new_n833), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n829), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT119), .B1(new_n823), .B2(new_n824), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n827), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n827), .A2(new_n843), .A3(KEYINPUT121), .A4(new_n844), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n825), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n840), .A3(new_n829), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n838), .A2(new_n839), .A3(new_n833), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n797), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n851), .A2(KEYINPUT53), .B1(new_n825), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n847), .A2(new_n848), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n763), .A2(new_n858), .A3(new_n489), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n763), .B2(new_n489), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n702), .A2(new_n744), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n861), .A2(new_n654), .A3(new_n732), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n622), .A2(new_n489), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n678), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n629), .A2(new_n636), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n723), .A2(new_n732), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n859), .B2(new_n860), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n684), .A2(new_n702), .A3(new_n560), .A4(new_n685), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT50), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n870), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n864), .B(new_n868), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n861), .A2(new_n869), .A3(new_n744), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n780), .B1(new_n775), .B2(new_n779), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n715), .A2(new_n496), .A3(new_n557), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n857), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n638), .A2(new_n640), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n488), .B(G953), .C1(new_n866), .C2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n834), .B2(new_n870), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n861), .A2(new_n747), .A3(new_n863), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT48), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(KEYINPUT48), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n876), .A2(new_n880), .A3(new_n857), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n786), .B1(new_n856), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n715), .A2(new_n557), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n686), .B(new_n678), .C1(KEYINPUT49), .C2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n762), .A2(new_n496), .A3(new_n560), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n723), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT116), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n894), .B(new_n897), .C1(KEYINPUT49), .C2(new_n893), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n241), .B1(new_n827), .B2(new_n843), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n583), .A2(new_n592), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n590), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n901), .B2(new_n902), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n189), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  AOI22_X1  g723(.A1(new_n851), .A2(new_n828), .B1(new_n822), .B2(new_n826), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n241), .A4(new_n769), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n912));
  INV_X1    g726(.A(new_n769), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n770), .B(KEYINPUT57), .Z(new_n916));
  AND3_X1   g730(.A1(new_n827), .A2(new_n843), .A3(new_n844), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n844), .B1(new_n827), .B2(new_n843), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n555), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n908), .B1(new_n915), .B2(new_n920), .ZN(G54));
  AND2_X1   g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n900), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n479), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(KEYINPUT124), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT124), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n900), .A2(new_n479), .A3(new_n922), .ZN(new_n927));
  INV_X1    g741(.A(new_n908), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  NOR2_X1   g746(.A1(new_n634), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n917), .B2(new_n918), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n928), .ZN(new_n935));
  INV_X1    g749(.A(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n856), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n634), .ZN(G63));
  OAI21_X1  g752(.A(new_n928), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n827), .B2(new_n843), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n942), .B2(new_n652), .ZN(new_n943));
  NAND2_X1  g757(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n260), .A2(new_n261), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n910), .B2(new_n941), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n491), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n785), .B1(new_n950), .B2(G224), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n852), .B2(new_n189), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n903), .B1(G898), .B2(new_n189), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(G69));
  INV_X1    g768(.A(new_n189), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(G227), .A3(G900), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n741), .A2(new_n809), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n688), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n783), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n392), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n802), .A2(new_n804), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n669), .A3(new_n744), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n776), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(new_n955), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n956), .B1(new_n961), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n364), .B(new_n451), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n973));
  INV_X1    g787(.A(G227), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n974), .A3(G900), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n955), .B(new_n975), .C1(new_n973), .C2(G900), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n783), .A2(new_n789), .A3(new_n754), .ZN(new_n977));
  INV_X1    g791(.A(new_n811), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n775), .A2(new_n668), .A3(new_n978), .A4(new_n747), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n977), .A2(new_n776), .A3(new_n957), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n970), .B(new_n976), .C1(new_n980), .C2(new_n955), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n972), .A2(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n980), .B2(new_n852), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n378), .A3(new_n671), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n967), .A2(new_n852), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n984), .B1(new_n961), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n672), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n986), .A2(new_n989), .A3(new_n928), .ZN(new_n990));
  INV_X1    g804(.A(new_n984), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n379), .A2(new_n383), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n366), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n990), .B1(new_n854), .B2(new_n993), .ZN(G57));
endmodule


