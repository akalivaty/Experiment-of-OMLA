

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752;

  OR2_X1 U377 ( .A1(n656), .A2(KEYINPUT85), .ZN(n501) );
  INV_X1 U378 ( .A(G953), .ZN(n730) );
  XNOR2_X1 U379 ( .A(n484), .B(n483), .ZN(n656) );
  XNOR2_X2 U380 ( .A(n513), .B(n368), .ZN(n491) );
  OR2_X2 U381 ( .A1(n662), .A2(G902), .ZN(n513) );
  NOR2_X2 U382 ( .A1(n582), .A2(n581), .ZN(n720) );
  XNOR2_X1 U383 ( .A(n509), .B(KEYINPUT106), .ZN(n557) );
  NOR2_X2 U384 ( .A1(n596), .A2(n723), .ZN(n562) );
  XNOR2_X2 U385 ( .A(n414), .B(n361), .ZN(n634) );
  AND2_X1 U386 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U387 ( .A(KEYINPUT46), .ZN(n563) );
  XNOR2_X1 U388 ( .A(n469), .B(n468), .ZN(n519) );
  BUF_X1 U389 ( .A(n509), .Z(n693) );
  XNOR2_X1 U390 ( .A(n536), .B(n535), .ZN(n731) );
  AND2_X1 U391 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U392 ( .A(n548), .B(n547), .ZN(n551) );
  XNOR2_X1 U393 ( .A(n489), .B(n488), .ZN(n526) );
  AND2_X1 U394 ( .A1(n643), .A2(n504), .ZN(n354) );
  OR2_X1 U395 ( .A1(n541), .A2(n450), .ZN(n355) );
  XOR2_X1 U396 ( .A(n400), .B(n399), .Z(n356) );
  OR2_X1 U397 ( .A1(n680), .A2(n577), .ZN(n578) );
  NAND2_X1 U398 ( .A1(n505), .A2(n354), .ZN(n507) );
  INV_X1 U399 ( .A(KEYINPUT70), .ZN(n590) );
  XNOR2_X1 U400 ( .A(n458), .B(G122), .ZN(n459) );
  XNOR2_X1 U401 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U402 ( .A(n564), .B(n563), .ZN(n593) );
  XNOR2_X1 U403 ( .A(n460), .B(n459), .ZN(n462) );
  NOR2_X1 U404 ( .A1(n598), .A2(n602), .ZN(n573) );
  NAND2_X1 U405 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U406 ( .A(n512), .B(KEYINPUT1), .ZN(n368) );
  XNOR2_X1 U407 ( .A(n453), .B(n452), .ZN(n514) );
  OR2_X1 U408 ( .A1(n526), .A2(n493), .ZN(n495) );
  OR2_X1 U409 ( .A1(n566), .A2(n565), .ZN(n721) );
  INV_X1 U410 ( .A(KEYINPUT60), .ZN(n628) );
  XNOR2_X2 U411 ( .A(KEYINPUT64), .B(G143), .ZN(n358) );
  INV_X1 U412 ( .A(G128), .ZN(n357) );
  XNOR2_X2 U413 ( .A(n358), .B(n357), .ZN(n421) );
  XNOR2_X2 U414 ( .A(n421), .B(G134), .ZN(n479) );
  XNOR2_X1 U415 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n359), .B(G131), .ZN(n465) );
  XNOR2_X2 U417 ( .A(n479), .B(n465), .ZN(n414) );
  INV_X1 U418 ( .A(KEYINPUT69), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n360), .B(G137), .ZN(n372) );
  XNOR2_X1 U420 ( .A(n372), .B(KEYINPUT93), .ZN(n361) );
  XNOR2_X1 U421 ( .A(G110), .B(G107), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n362), .B(G104), .ZN(n739) );
  XNOR2_X1 U423 ( .A(KEYINPUT4), .B(G101), .ZN(n403) );
  XNOR2_X1 U424 ( .A(n739), .B(n403), .ZN(n429) );
  NAND2_X1 U425 ( .A1(n730), .A2(G227), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n363), .B(G140), .ZN(n365) );
  XNOR2_X1 U427 ( .A(G146), .B(KEYINPUT94), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n429), .B(n366), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n634), .B(n367), .ZN(n662) );
  XNOR2_X1 U431 ( .A(KEYINPUT71), .B(G469), .ZN(n512) );
  NAND2_X1 U432 ( .A1(n730), .A2(G234), .ZN(n370) );
  INV_X1 U433 ( .A(KEYINPUT8), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n475) );
  NAND2_X1 U435 ( .A1(G221), .A2(n475), .ZN(n377) );
  INV_X1 U436 ( .A(KEYINPUT24), .ZN(n371) );
  NAND2_X1 U437 ( .A1(n372), .A2(n371), .ZN(n375) );
  INV_X1 U438 ( .A(n372), .ZN(n373) );
  NAND2_X1 U439 ( .A1(n373), .A2(KEYINPUT24), .ZN(n374) );
  NAND2_X1 U440 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n384) );
  XOR2_X1 U442 ( .A(KEYINPUT23), .B(G110), .Z(n379) );
  XNOR2_X1 U443 ( .A(G119), .B(G128), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n382) );
  XNOR2_X1 U445 ( .A(G146), .B(G125), .ZN(n426) );
  INV_X1 U446 ( .A(KEYINPUT10), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n380), .B(G140), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n426), .B(n381), .ZN(n632) );
  XNOR2_X1 U449 ( .A(n382), .B(n632), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n651) );
  INV_X1 U451 ( .A(G902), .ZN(n480) );
  NAND2_X1 U452 ( .A1(n651), .A2(n480), .ZN(n391) );
  XNOR2_X1 U453 ( .A(KEYINPUT15), .B(G902), .ZN(n436) );
  NAND2_X1 U454 ( .A1(n436), .A2(G234), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n385), .B(KEYINPUT20), .ZN(n392) );
  NAND2_X1 U456 ( .A1(G217), .A2(n392), .ZN(n389) );
  XOR2_X1 U457 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n387) );
  XNOR2_X1 U458 ( .A(KEYINPUT78), .B(KEYINPUT96), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U460 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X2 U461 ( .A(n391), .B(n390), .ZN(n490) );
  INV_X1 U462 ( .A(n490), .ZN(n396) );
  NAND2_X1 U463 ( .A1(G221), .A2(n392), .ZN(n394) );
  XOR2_X1 U464 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n393) );
  XNOR2_X1 U465 ( .A(n394), .B(n393), .ZN(n690) );
  INV_X1 U466 ( .A(n690), .ZN(n395) );
  NAND2_X1 U467 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n397), .B(KEYINPUT66), .ZN(n688) );
  OR2_X1 U469 ( .A1(n491), .A2(n688), .ZN(n510) );
  XNOR2_X1 U470 ( .A(n510), .B(KEYINPUT107), .ZN(n418) );
  XNOR2_X1 U471 ( .A(G146), .B(G137), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n398), .B(KEYINPUT99), .ZN(n400) );
  XOR2_X1 U473 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n399) );
  NOR2_X1 U474 ( .A1(G953), .A2(G237), .ZN(n463) );
  NAND2_X1 U475 ( .A1(n463), .A2(G210), .ZN(n402) );
  XOR2_X1 U476 ( .A(KEYINPUT75), .B(KEYINPUT100), .Z(n401) );
  XNOR2_X1 U477 ( .A(n402), .B(n401), .ZN(n404) );
  XNOR2_X1 U478 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U479 ( .A(n356), .B(n405), .ZN(n411) );
  INV_X1 U480 ( .A(n411), .ZN(n410) );
  XNOR2_X1 U481 ( .A(G119), .B(G116), .ZN(n406) );
  XNOR2_X1 U482 ( .A(n406), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U483 ( .A(G113), .B(KEYINPUT72), .ZN(n407) );
  XNOR2_X1 U484 ( .A(n408), .B(n407), .ZN(n434) );
  INV_X1 U485 ( .A(n434), .ZN(n409) );
  NAND2_X1 U486 ( .A1(n410), .A2(n409), .ZN(n413) );
  NAND2_X1 U487 ( .A1(n411), .A2(n434), .ZN(n412) );
  NAND2_X1 U488 ( .A1(n413), .A2(n412), .ZN(n415) );
  XNOR2_X2 U489 ( .A(n415), .B(n414), .ZN(n645) );
  NAND2_X1 U490 ( .A1(n645), .A2(n480), .ZN(n416) );
  XNOR2_X2 U491 ( .A(n416), .B(G472), .ZN(n509) );
  INV_X1 U492 ( .A(KEYINPUT6), .ZN(n417) );
  XNOR2_X1 U493 ( .A(n509), .B(n417), .ZN(n568) );
  NAND2_X1 U494 ( .A1(n418), .A2(n568), .ZN(n420) );
  INV_X1 U495 ( .A(KEYINPUT33), .ZN(n419) );
  XNOR2_X1 U496 ( .A(n420), .B(n419), .ZN(n684) );
  INV_X1 U497 ( .A(n421), .ZN(n424) );
  NAND2_X1 U498 ( .A1(n730), .A2(G224), .ZN(n422) );
  XNOR2_X1 U499 ( .A(n422), .B(KEYINPUT79), .ZN(n423) );
  XNOR2_X1 U500 ( .A(n424), .B(n423), .ZN(n428) );
  XNOR2_X1 U501 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n425) );
  XNOR2_X1 U502 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U503 ( .A(n428), .B(n427), .ZN(n431) );
  INV_X1 U504 ( .A(n429), .ZN(n430) );
  XNOR2_X1 U505 ( .A(n431), .B(n430), .ZN(n435) );
  XNOR2_X1 U506 ( .A(KEYINPUT16), .B(G122), .ZN(n432) );
  XNOR2_X1 U507 ( .A(n432), .B(KEYINPUT74), .ZN(n433) );
  XNOR2_X1 U508 ( .A(n434), .B(n433), .ZN(n742) );
  XNOR2_X1 U509 ( .A(n435), .B(n742), .ZN(n616) );
  INV_X1 U510 ( .A(n436), .ZN(n609) );
  OR2_X2 U511 ( .A1(n616), .A2(n609), .ZN(n441) );
  INV_X1 U512 ( .A(G237), .ZN(n437) );
  NAND2_X1 U513 ( .A1(n480), .A2(n437), .ZN(n442) );
  NAND2_X1 U514 ( .A1(n442), .A2(G210), .ZN(n439) );
  INV_X1 U515 ( .A(KEYINPUT90), .ZN(n438) );
  XNOR2_X1 U516 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X2 U517 ( .A(n441), .B(n440), .ZN(n572) );
  NAND2_X1 U518 ( .A1(n442), .A2(G214), .ZN(n674) );
  NAND2_X1 U519 ( .A1(n572), .A2(n674), .ZN(n444) );
  XNOR2_X1 U520 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n443) );
  XNOR2_X1 U521 ( .A(n444), .B(n443), .ZN(n565) );
  INV_X1 U522 ( .A(n565), .ZN(n451) );
  NAND2_X1 U523 ( .A1(G234), .A2(G237), .ZN(n445) );
  XNOR2_X1 U524 ( .A(n445), .B(KEYINPUT14), .ZN(n447) );
  NAND2_X1 U525 ( .A1(n447), .A2(G952), .ZN(n446) );
  XNOR2_X1 U526 ( .A(n446), .B(KEYINPUT91), .ZN(n703) );
  AND2_X1 U527 ( .A1(n703), .A2(n730), .ZN(n541) );
  NAND2_X1 U528 ( .A1(G902), .A2(n447), .ZN(n542) );
  INV_X1 U529 ( .A(G898), .ZN(n448) );
  NAND2_X1 U530 ( .A1(n448), .A2(G953), .ZN(n449) );
  XNOR2_X1 U531 ( .A(n449), .B(KEYINPUT92), .ZN(n743) );
  NOR2_X1 U532 ( .A1(n542), .A2(n743), .ZN(n450) );
  NAND2_X1 U533 ( .A1(n451), .A2(n355), .ZN(n453) );
  XNOR2_X1 U534 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n452) );
  OR2_X1 U535 ( .A1(n684), .A2(n514), .ZN(n455) );
  INV_X1 U536 ( .A(KEYINPUT34), .ZN(n454) );
  XNOR2_X1 U537 ( .A(n455), .B(n454), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n457) );
  XNOR2_X1 U539 ( .A(G104), .B(KEYINPUT101), .ZN(n456) );
  XNOR2_X1 U540 ( .A(n457), .B(n456), .ZN(n460) );
  XOR2_X1 U541 ( .A(G113), .B(G143), .Z(n458) );
  INV_X1 U542 ( .A(n632), .ZN(n461) );
  XNOR2_X1 U543 ( .A(n462), .B(n461), .ZN(n467) );
  NAND2_X1 U544 ( .A1(G214), .A2(n463), .ZN(n464) );
  XNOR2_X1 U545 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U546 ( .A(n467), .B(n466), .ZN(n624) );
  NAND2_X1 U547 ( .A1(n624), .A2(n480), .ZN(n469) );
  XOR2_X1 U548 ( .A(KEYINPUT13), .B(G475), .Z(n468) );
  XNOR2_X1 U549 ( .A(G116), .B(KEYINPUT104), .ZN(n470) );
  XNOR2_X1 U550 ( .A(n470), .B(KEYINPUT9), .ZN(n474) );
  XOR2_X1 U551 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n472) );
  XNOR2_X1 U552 ( .A(G107), .B(G122), .ZN(n471) );
  XNOR2_X1 U553 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U554 ( .A(n474), .B(n473), .Z(n477) );
  AND2_X1 U555 ( .A1(n475), .A2(G217), .ZN(n476) );
  XNOR2_X1 U556 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U557 ( .A(n479), .B(n478), .ZN(n658) );
  NAND2_X1 U558 ( .A1(n658), .A2(n480), .ZN(n481) );
  XNOR2_X1 U559 ( .A(n481), .B(G478), .ZN(n521) );
  AND2_X1 U560 ( .A1(n519), .A2(n521), .ZN(n580) );
  NAND2_X1 U561 ( .A1(n482), .A2(n580), .ZN(n484) );
  INV_X1 U562 ( .A(KEYINPUT35), .ZN(n483) );
  INV_X1 U563 ( .A(n514), .ZN(n486) );
  OR2_X1 U564 ( .A1(n519), .A2(n521), .ZN(n539) );
  NOR2_X1 U565 ( .A1(n539), .A2(n690), .ZN(n485) );
  NAND2_X1 U566 ( .A1(n486), .A2(n485), .ZN(n489) );
  INV_X1 U567 ( .A(KEYINPUT73), .ZN(n487) );
  XNOR2_X1 U568 ( .A(n487), .B(KEYINPUT22), .ZN(n488) );
  INV_X1 U569 ( .A(n490), .ZN(n496) );
  OR2_X1 U570 ( .A1(n568), .A2(n496), .ZN(n492) );
  OR2_X1 U571 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U572 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n494) );
  XNOR2_X2 U573 ( .A(n495), .B(n494), .ZN(n505) );
  NOR2_X1 U574 ( .A1(n557), .A2(n496), .ZN(n497) );
  NAND2_X1 U575 ( .A1(n497), .A2(n491), .ZN(n498) );
  OR2_X1 U576 ( .A1(n526), .A2(n498), .ZN(n643) );
  AND2_X1 U577 ( .A1(n643), .A2(KEYINPUT44), .ZN(n499) );
  AND2_X1 U578 ( .A1(n505), .A2(n499), .ZN(n500) );
  NAND2_X1 U579 ( .A1(n501), .A2(n500), .ZN(n503) );
  INV_X1 U580 ( .A(KEYINPUT85), .ZN(n506) );
  INV_X1 U581 ( .A(KEYINPUT44), .ZN(n504) );
  NAND2_X1 U582 ( .A1(n506), .A2(n504), .ZN(n502) );
  NAND2_X1 U583 ( .A1(n503), .A2(n502), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U585 ( .A1(n508), .A2(n656), .ZN(n532) );
  INV_X1 U586 ( .A(n693), .ZN(n517) );
  OR2_X1 U587 ( .A1(n510), .A2(n517), .ZN(n696) );
  NOR2_X1 U588 ( .A1(n696), .A2(n514), .ZN(n511) );
  XNOR2_X1 U589 ( .A(n511), .B(KEYINPUT31), .ZN(n725) );
  XNOR2_X1 U590 ( .A(n513), .B(n512), .ZN(n549) );
  OR2_X1 U591 ( .A1(n688), .A2(n549), .ZN(n554) );
  OR2_X1 U592 ( .A1(n514), .A2(n554), .ZN(n516) );
  INV_X1 U593 ( .A(KEYINPUT98), .ZN(n515) );
  XNOR2_X1 U594 ( .A(n516), .B(n515), .ZN(n518) );
  NAND2_X1 U595 ( .A1(n518), .A2(n517), .ZN(n715) );
  NAND2_X1 U596 ( .A1(n725), .A2(n715), .ZN(n525) );
  XNOR2_X1 U597 ( .A(KEYINPUT102), .B(n519), .ZN(n523) );
  INV_X1 U598 ( .A(n523), .ZN(n520) );
  NAND2_X1 U599 ( .A1(n520), .A2(n521), .ZN(n726) );
  INV_X1 U600 ( .A(n521), .ZN(n522) );
  NAND2_X1 U601 ( .A1(n523), .A2(n522), .ZN(n723) );
  AND2_X1 U602 ( .A1(n726), .A2(n723), .ZN(n524) );
  XNOR2_X1 U603 ( .A(n524), .B(KEYINPUT105), .ZN(n680) );
  NAND2_X1 U604 ( .A1(n525), .A2(n680), .ZN(n530) );
  INV_X1 U605 ( .A(n526), .ZN(n529) );
  INV_X1 U606 ( .A(n491), .ZN(n597) );
  OR2_X1 U607 ( .A1(n568), .A2(n490), .ZN(n527) );
  NOR2_X1 U608 ( .A1(n597), .A2(n527), .ZN(n528) );
  NAND2_X1 U609 ( .A1(n529), .A2(n528), .ZN(n631) );
  AND2_X1 U610 ( .A1(n530), .A2(n631), .ZN(n531) );
  XNOR2_X1 U611 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n535) );
  INV_X1 U612 ( .A(KEYINPUT38), .ZN(n537) );
  XNOR2_X1 U613 ( .A(n572), .B(n537), .ZN(n675) );
  NAND2_X1 U614 ( .A1(n675), .A2(n674), .ZN(n538) );
  XNOR2_X1 U615 ( .A(KEYINPUT111), .B(n538), .ZN(n681) );
  INV_X1 U616 ( .A(n539), .ZN(n677) );
  NAND2_X1 U617 ( .A1(n681), .A2(n677), .ZN(n540) );
  XOR2_X1 U618 ( .A(KEYINPUT41), .B(n540), .Z(n705) );
  INV_X1 U619 ( .A(n541), .ZN(n545) );
  NOR2_X1 U620 ( .A1(G900), .A2(n542), .ZN(n543) );
  NAND2_X1 U621 ( .A1(G953), .A2(n543), .ZN(n544) );
  NAND2_X1 U622 ( .A1(n545), .A2(n544), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n490), .A2(n555), .ZN(n546) );
  NOR2_X1 U624 ( .A1(n690), .A2(n546), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n570), .A2(n557), .ZN(n548) );
  XOR2_X1 U626 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n547) );
  INV_X1 U627 ( .A(n549), .ZN(n550) );
  NAND2_X1 U628 ( .A1(n551), .A2(n550), .ZN(n566) );
  NOR2_X1 U629 ( .A1(n705), .A2(n566), .ZN(n553) );
  XNOR2_X1 U630 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n552) );
  XNOR2_X1 U631 ( .A(n553), .B(n552), .ZN(n747) );
  XNOR2_X1 U632 ( .A(n554), .B(KEYINPUT109), .ZN(n556) );
  NAND2_X1 U633 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U634 ( .A1(n557), .A2(n674), .ZN(n558) );
  XNOR2_X1 U635 ( .A(n558), .B(KEYINPUT30), .ZN(n559) );
  NOR2_X1 U636 ( .A1(n560), .A2(n559), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n579), .A2(n675), .ZN(n561) );
  XOR2_X1 U638 ( .A(n561), .B(KEYINPUT39), .Z(n596) );
  XNOR2_X1 U639 ( .A(n562), .B(KEYINPUT40), .ZN(n752) );
  NOR2_X1 U640 ( .A1(n747), .A2(n752), .ZN(n564) );
  NOR2_X1 U641 ( .A1(n721), .A2(KEYINPUT47), .ZN(n567) );
  AND2_X1 U642 ( .A1(n567), .A2(n680), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n568), .A2(n674), .ZN(n569) );
  NOR2_X1 U644 ( .A1(n723), .A2(n569), .ZN(n571) );
  NAND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n598) );
  INV_X1 U646 ( .A(n572), .ZN(n602) );
  XNOR2_X1 U647 ( .A(n573), .B(KEYINPUT36), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n574), .A2(n597), .ZN(n575) );
  XNOR2_X1 U649 ( .A(n575), .B(KEYINPUT113), .ZN(n749) );
  NOR2_X1 U650 ( .A1(n576), .A2(n749), .ZN(n589) );
  INV_X1 U651 ( .A(KEYINPUT47), .ZN(n577) );
  XNOR2_X1 U652 ( .A(n578), .B(KEYINPUT83), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n721), .A2(KEYINPUT47), .ZN(n584) );
  INV_X1 U654 ( .A(n579), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n580), .A2(n572), .ZN(n581) );
  INV_X1 U656 ( .A(n720), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT82), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n595) );
  INV_X1 U661 ( .A(KEYINPUT48), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n595), .B(n594), .ZN(n605) );
  NOR2_X1 U663 ( .A1(n596), .A2(n726), .ZN(n729) );
  NOR2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n601) );
  INV_X1 U665 ( .A(KEYINPUT108), .ZN(n599) );
  XNOR2_X1 U666 ( .A(n599), .B(KEYINPUT43), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n601), .B(n600), .ZN(n603) );
  AND2_X1 U668 ( .A1(n603), .A2(n602), .ZN(n630) );
  OR2_X1 U669 ( .A1(n729), .A2(n630), .ZN(n604) );
  NOR2_X2 U670 ( .A1(n605), .A2(n604), .ZN(n635) );
  NAND2_X1 U671 ( .A1(n731), .A2(n635), .ZN(n670) );
  INV_X1 U672 ( .A(KEYINPUT65), .ZN(n606) );
  NAND2_X1 U673 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  NAND2_X1 U674 ( .A1(n670), .A2(n607), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n608), .A2(n609), .ZN(n612) );
  NAND2_X1 U676 ( .A1(n609), .A2(KEYINPUT2), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n610), .A2(KEYINPUT65), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U679 ( .A(n670), .ZN(n669) );
  NAND2_X1 U680 ( .A1(n669), .A2(KEYINPUT2), .ZN(n613) );
  AND2_X2 U681 ( .A1(n614), .A2(n613), .ZN(n661) );
  NAND2_X1 U682 ( .A1(n661), .A2(G210), .ZN(n618) );
  XNOR2_X1 U683 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n615) );
  XNOR2_X1 U684 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U685 ( .A(n618), .B(n617), .ZN(n620) );
  INV_X1 U686 ( .A(G952), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n619), .A2(G953), .ZN(n659) );
  NAND2_X1 U688 ( .A1(n620), .A2(n659), .ZN(n622) );
  INV_X1 U689 ( .A(KEYINPUT56), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n622), .B(n621), .ZN(G51) );
  NAND2_X1 U691 ( .A1(n661), .A2(G475), .ZN(n626) );
  XOR2_X1 U692 ( .A(KEYINPUT88), .B(KEYINPUT59), .Z(n623) );
  XNOR2_X1 U693 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n627), .A2(n659), .ZN(n629) );
  XNOR2_X1 U696 ( .A(n629), .B(n628), .ZN(G60) );
  XOR2_X1 U697 ( .A(G140), .B(n630), .Z(G42) );
  XNOR2_X1 U698 ( .A(n631), .B(G101), .ZN(G3) );
  XOR2_X1 U699 ( .A(KEYINPUT4), .B(n632), .Z(n633) );
  XNOR2_X1 U700 ( .A(n634), .B(n633), .ZN(n638) );
  XNOR2_X1 U701 ( .A(n638), .B(KEYINPUT126), .ZN(n636) );
  XOR2_X1 U702 ( .A(n636), .B(n635), .Z(n637) );
  NAND2_X1 U703 ( .A1(n637), .A2(n730), .ZN(n642) );
  XNOR2_X1 U704 ( .A(G227), .B(n638), .ZN(n639) );
  NAND2_X1 U705 ( .A1(n639), .A2(G900), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n640), .A2(G953), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n642), .A2(n641), .ZN(G72) );
  XNOR2_X1 U708 ( .A(n643), .B(G110), .ZN(G12) );
  NAND2_X1 U709 ( .A1(n661), .A2(G472), .ZN(n647) );
  XOR2_X1 U710 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n648), .A2(n659), .ZN(n650) );
  XOR2_X1 U714 ( .A(KEYINPUT89), .B(KEYINPUT63), .Z(n649) );
  XNOR2_X1 U715 ( .A(n650), .B(n649), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n661), .A2(G217), .ZN(n653) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT120), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n654), .A2(n659), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n655), .B(KEYINPUT121), .ZN(G66) );
  XNOR2_X1 U721 ( .A(n656), .B(G122), .ZN(G24) );
  XNOR2_X1 U722 ( .A(n505), .B(G119), .ZN(G21) );
  NAND2_X1 U723 ( .A1(n661), .A2(G478), .ZN(n657) );
  XOR2_X1 U724 ( .A(n658), .B(n657), .Z(n660) );
  INV_X1 U725 ( .A(n659), .ZN(n666) );
  NOR2_X1 U726 ( .A1(n660), .A2(n666), .ZN(G63) );
  NAND2_X1 U727 ( .A1(n661), .A2(G469), .ZN(n665) );
  XOR2_X1 U728 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n663) );
  XNOR2_X1 U729 ( .A(n662), .B(n663), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n665), .B(n664), .ZN(n667) );
  NOR2_X1 U731 ( .A1(n667), .A2(n666), .ZN(G54) );
  XOR2_X1 U732 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n668) );
  NOR2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U734 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n670), .A2(n671), .ZN(n672) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n710) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U738 ( .A(KEYINPUT117), .B(n676), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n679), .B(KEYINPUT118), .ZN(n683) );
  NAND2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n686) );
  INV_X1 U743 ( .A(n684), .ZN(n685) );
  NAND2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n687), .B(KEYINPUT119), .ZN(n701) );
  NAND2_X1 U746 ( .A1(n491), .A2(n688), .ZN(n689) );
  XNOR2_X1 U747 ( .A(n689), .B(KEYINPUT50), .ZN(n695) );
  NAND2_X1 U748 ( .A1(n490), .A2(n690), .ZN(n691) );
  XNOR2_X1 U749 ( .A(KEYINPUT49), .B(n691), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U751 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U753 ( .A(KEYINPUT51), .B(n698), .ZN(n699) );
  NOR2_X1 U754 ( .A1(n705), .A2(n699), .ZN(n700) );
  OR2_X1 U755 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n702), .B(KEYINPUT52), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U758 ( .A1(n705), .A2(n684), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n706), .A2(G953), .ZN(n707) );
  NAND2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U761 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n711), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U763 ( .A1(n723), .A2(n715), .ZN(n712) );
  XOR2_X1 U764 ( .A(G104), .B(n712), .Z(G6) );
  XOR2_X1 U765 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n714) );
  XNOR2_X1 U766 ( .A(G107), .B(KEYINPUT27), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n714), .B(n713), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n726), .A2(n715), .ZN(n716) );
  XOR2_X1 U769 ( .A(n717), .B(n716), .Z(G9) );
  NOR2_X1 U770 ( .A1(n721), .A2(n726), .ZN(n719) );
  XNOR2_X1 U771 ( .A(G128), .B(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(G30) );
  XOR2_X1 U773 ( .A(G143), .B(n720), .Z(G45) );
  NOR2_X1 U774 ( .A1(n721), .A2(n723), .ZN(n722) );
  XOR2_X1 U775 ( .A(G146), .B(n722), .Z(G48) );
  NOR2_X1 U776 ( .A1(n723), .A2(n725), .ZN(n724) );
  XOR2_X1 U777 ( .A(G113), .B(n724), .Z(G15) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U779 ( .A(G116), .B(KEYINPUT115), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(G18) );
  XOR2_X1 U781 ( .A(G134), .B(n729), .Z(G36) );
  AND2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n736) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(KEYINPUT122), .ZN(n733) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n733), .ZN(n734) );
  AND2_X1 U786 ( .A1(n734), .A2(G898), .ZN(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U788 ( .A(n737), .B(KEYINPUT125), .Z(n746) );
  XOR2_X1 U789 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n738) );
  XNOR2_X1 U790 ( .A(n738), .B(G101), .ZN(n740) );
  XOR2_X1 U791 ( .A(n740), .B(n739), .Z(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(G69) );
  XNOR2_X1 U795 ( .A(G137), .B(n747), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n748), .B(KEYINPUT127), .ZN(G39) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT116), .ZN(n750) );
  XNOR2_X1 U798 ( .A(n750), .B(KEYINPUT37), .ZN(n751) );
  XNOR2_X1 U799 ( .A(G125), .B(n751), .ZN(G27) );
  XOR2_X1 U800 ( .A(G131), .B(n752), .Z(G33) );
endmodule

