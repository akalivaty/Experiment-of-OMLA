

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765;

  AND2_X1 U374 ( .A1(n387), .A2(n385), .ZN(n384) );
  XOR2_X1 U375 ( .A(n752), .B(n506), .Z(n351) );
  XOR2_X1 U376 ( .A(n598), .B(KEYINPUT109), .Z(n352) );
  XNOR2_X2 U377 ( .A(n628), .B(KEYINPUT64), .ZN(n632) );
  INV_X2 U378 ( .A(KEYINPUT71), .ZN(n398) );
  XNOR2_X2 U379 ( .A(n474), .B(n473), .ZN(n557) );
  XNOR2_X2 U380 ( .A(n592), .B(KEYINPUT39), .ZN(n624) );
  XNOR2_X2 U381 ( .A(n593), .B(KEYINPUT40), .ZN(n764) );
  AND2_X2 U382 ( .A1(n624), .A2(n676), .ZN(n593) );
  AND2_X1 U383 ( .A1(n614), .A2(n613), .ZN(n617) );
  NOR2_X1 U384 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U385 ( .A(n619), .ZN(n700) );
  INV_X2 U386 ( .A(G146), .ZN(n410) );
  NAND2_X1 U387 ( .A1(n372), .A2(n371), .ZN(n628) );
  NAND2_X1 U388 ( .A1(n402), .A2(n401), .ZN(n400) );
  XNOR2_X1 U389 ( .A(n617), .B(n616), .ZN(n406) );
  AND2_X1 U390 ( .A1(n531), .A2(KEYINPUT44), .ZN(n532) );
  OR2_X1 U391 ( .A1(n763), .A2(KEYINPUT89), .ZN(n531) );
  NAND2_X1 U392 ( .A1(n380), .A2(n554), .ZN(n645) );
  XNOR2_X1 U393 ( .A(n437), .B(n360), .ZN(n503) );
  XNOR2_X1 U394 ( .A(n478), .B(G140), .ZN(n501) );
  NOR2_X2 U395 ( .A1(n584), .A2(n522), .ZN(n701) );
  INV_X1 U396 ( .A(n602), .ZN(n353) );
  XNOR2_X1 U397 ( .A(n521), .B(n520), .ZN(n354) );
  XNOR2_X1 U398 ( .A(n391), .B(KEYINPUT19), .ZN(n670) );
  OR2_X2 U399 ( .A1(n377), .A2(n374), .ZN(n581) );
  AND2_X2 U400 ( .A1(n399), .A2(n403), .ZN(n368) );
  XNOR2_X2 U401 ( .A(n369), .B(G134), .ZN(n397) );
  XNOR2_X2 U402 ( .A(n410), .B(G125), .ZN(n437) );
  INV_X1 U403 ( .A(G137), .ZN(n478) );
  INV_X1 U404 ( .A(KEYINPUT10), .ZN(n360) );
  NAND2_X1 U405 ( .A1(n635), .A2(n512), .ZN(n589) );
  XNOR2_X1 U406 ( .A(n471), .B(n470), .ZN(n525) );
  OR2_X1 U407 ( .A1(n550), .A2(n551), .ZN(n691) );
  NAND2_X1 U408 ( .A1(n376), .A2(n512), .ZN(n375) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n487) );
  INV_X1 U410 ( .A(KEYINPUT111), .ZN(n395) );
  NAND2_X1 U411 ( .A1(n581), .A2(n582), .ZN(n583) );
  NAND2_X1 U412 ( .A1(n458), .A2(n627), .ZN(n389) );
  INV_X1 U413 ( .A(KEYINPUT87), .ZN(n401) );
  XNOR2_X1 U414 ( .A(n503), .B(n502), .ZN(n752) );
  XNOR2_X1 U415 ( .A(n361), .B(n423), .ZN(n507) );
  XNOR2_X1 U416 ( .A(n424), .B(n363), .ZN(n361) );
  INV_X1 U417 ( .A(KEYINPUT85), .ZN(n363) );
  NAND2_X1 U418 ( .A1(n754), .A2(n626), .ZN(n371) );
  NAND2_X1 U419 ( .A1(n352), .A2(n355), .ZN(n618) );
  BUF_X1 U420 ( .A(n584), .Z(n554) );
  XNOR2_X1 U421 ( .A(n433), .B(n432), .ZN(n547) );
  XNOR2_X1 U422 ( .A(n431), .B(KEYINPUT105), .ZN(n432) );
  XNOR2_X1 U423 ( .A(n575), .B(n500), .ZN(n597) );
  NOR2_X1 U424 ( .A1(n669), .A2(n713), .ZN(n580) );
  NOR2_X1 U425 ( .A1(n669), .A2(n602), .ZN(n675) );
  NAND2_X1 U426 ( .A1(n603), .A2(n675), .ZN(n365) );
  INV_X1 U427 ( .A(G237), .ZN(n457) );
  XOR2_X1 U428 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n489) );
  XOR2_X1 U429 ( .A(KEYINPUT78), .B(G113), .Z(n494) );
  XNOR2_X1 U430 ( .A(G137), .B(G116), .ZN(n493) );
  NOR2_X1 U431 ( .A1(n405), .A2(n404), .ZN(n403) );
  INV_X1 U432 ( .A(n686), .ZN(n404) );
  NOR2_X1 U433 ( .A1(n644), .A2(KEYINPUT87), .ZN(n405) );
  XNOR2_X1 U434 ( .A(n501), .B(n479), .ZN(n481) );
  INV_X1 U435 ( .A(KEYINPUT68), .ZN(n443) );
  XNOR2_X1 U436 ( .A(KEYINPUT95), .B(KEYINPUT17), .ZN(n442) );
  XNOR2_X1 U437 ( .A(KEYINPUT18), .B(KEYINPUT94), .ZN(n441) );
  NAND2_X1 U438 ( .A1(G234), .A2(G237), .ZN(n461) );
  BUF_X1 U439 ( .A(n525), .Z(n540) );
  NAND2_X1 U440 ( .A1(G469), .A2(G902), .ZN(n378) );
  INV_X1 U441 ( .A(G953), .ZN(n463) );
  INV_X1 U442 ( .A(KEYINPUT3), .ZN(n450) );
  XNOR2_X1 U443 ( .A(KEYINPUT77), .B(KEYINPUT16), .ZN(n447) );
  XNOR2_X1 U444 ( .A(G113), .B(G104), .ZN(n452) );
  XNOR2_X1 U445 ( .A(n412), .B(n411), .ZN(n413) );
  INV_X1 U446 ( .A(G122), .ZN(n411) );
  NOR2_X1 U447 ( .A1(n692), .A2(n691), .ZN(n579) );
  XNOR2_X1 U448 ( .A(n591), .B(n394), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n590), .B(n395), .ZN(n394) );
  NAND2_X1 U450 ( .A1(n383), .A2(n390), .ZN(n622) );
  XNOR2_X1 U451 ( .A(n351), .B(n511), .ZN(n651) );
  AND2_X1 U452 ( .A1(n373), .A2(n627), .ZN(n372) );
  NOR2_X1 U453 ( .A1(n600), .A2(n599), .ZN(n684) );
  XNOR2_X1 U454 ( .A(n367), .B(n366), .ZN(n599) );
  INV_X1 U455 ( .A(KEYINPUT36), .ZN(n366) );
  NOR2_X1 U456 ( .A1(n618), .A2(n622), .ZN(n367) );
  XNOR2_X1 U457 ( .A(n382), .B(n519), .ZN(n642) );
  NOR2_X1 U458 ( .A1(n575), .A2(n596), .ZN(n576) );
  NOR2_X1 U459 ( .A1(n386), .A2(n460), .ZN(n385) );
  XNOR2_X1 U460 ( .A(n381), .B(KEYINPUT67), .ZN(n380) );
  XNOR2_X1 U461 ( .A(n549), .B(n548), .ZN(n678) );
  NOR2_X1 U462 ( .A1(n727), .A2(G953), .ZN(n364) );
  NOR2_X1 U463 ( .A1(n678), .A2(n460), .ZN(n355) );
  XNOR2_X1 U464 ( .A(n589), .B(n588), .ZN(n699) );
  NOR2_X1 U465 ( .A1(n600), .A2(n518), .ZN(n356) );
  XOR2_X1 U466 ( .A(KEYINPUT86), .B(n726), .Z(n357) );
  AND2_X1 U467 ( .A1(n619), .A2(n575), .ZN(n358) );
  AND2_X1 U468 ( .A1(n644), .A2(KEYINPUT87), .ZN(n359) );
  BUF_X1 U469 ( .A(n463), .Z(n755) );
  NAND2_X1 U470 ( .A1(n730), .A2(G469), .ZN(n379) );
  NAND2_X1 U471 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X2 U472 ( .A(n622), .B(KEYINPUT38), .ZN(n689) );
  NOR2_X2 U473 ( .A1(n541), .A2(n597), .ZN(n362) );
  NAND2_X1 U474 ( .A1(n384), .A2(n390), .ZN(n391) );
  BUF_X2 U475 ( .A(n630), .Z(n741) );
  XNOR2_X2 U476 ( .A(n362), .B(n524), .ZN(n697) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n646) );
  NAND2_X1 U478 ( .A1(n357), .A2(n364), .ZN(n728) );
  XNOR2_X1 U479 ( .A(n503), .B(n413), .ZN(n415) );
  INV_X1 U480 ( .A(n365), .ZN(n610) );
  NAND2_X1 U481 ( .A1(n365), .A2(KEYINPUT47), .ZN(n608) );
  NAND2_X2 U482 ( .A1(n368), .A2(n400), .ZN(n754) );
  NOR2_X1 U483 ( .A1(n596), .A2(n597), .ZN(n598) );
  XNOR2_X2 U484 ( .A(n589), .B(n587), .ZN(n575) );
  INV_X1 U485 ( .A(n754), .ZN(n629) );
  XNOR2_X1 U486 ( .A(n369), .B(G143), .ZN(n414) );
  XNOR2_X2 U487 ( .A(n398), .B(G131), .ZN(n369) );
  NAND2_X1 U488 ( .A1(n370), .A2(n626), .ZN(n392) );
  OR2_X1 U489 ( .A1(n754), .A2(n741), .ZN(n370) );
  NAND2_X1 U490 ( .A1(n630), .A2(n626), .ZN(n373) );
  NOR2_X1 U491 ( .A1(n730), .A2(n375), .ZN(n374) );
  INV_X1 U492 ( .A(G469), .ZN(n376) );
  XNOR2_X2 U493 ( .A(n498), .B(n484), .ZN(n730) );
  XNOR2_X2 U494 ( .A(n581), .B(n485), .ZN(n619) );
  NAND2_X1 U495 ( .A1(n642), .A2(n645), .ZN(n521) );
  NAND2_X1 U496 ( .A1(n557), .A2(n358), .ZN(n381) );
  NAND2_X1 U497 ( .A1(n557), .A2(n356), .ZN(n382) );
  AND2_X1 U498 ( .A1(n387), .A2(n389), .ZN(n383) );
  INV_X1 U499 ( .A(n389), .ZN(n386) );
  OR2_X2 U500 ( .A1(n656), .A2(n388), .ZN(n387) );
  OR2_X1 U501 ( .A1(n627), .A2(n458), .ZN(n388) );
  NAND2_X1 U502 ( .A1(n656), .A2(n458), .ZN(n390) );
  XNOR2_X1 U503 ( .A(n392), .B(KEYINPUT83), .ZN(n725) );
  NAND2_X1 U504 ( .A1(n607), .A2(n689), .ZN(n592) );
  AND2_X2 U505 ( .A1(n396), .A2(n393), .ZN(n607) );
  XNOR2_X1 U506 ( .A(n585), .B(n586), .ZN(n396) );
  XNOR2_X2 U507 ( .A(n753), .B(n477), .ZN(n498) );
  XNOR2_X2 U508 ( .A(n397), .B(n476), .ZN(n753) );
  XNOR2_X2 U509 ( .A(n439), .B(KEYINPUT4), .ZN(n476) );
  XNOR2_X2 U510 ( .A(G143), .B(G128), .ZN(n439) );
  NAND2_X1 U511 ( .A1(n406), .A2(n359), .ZN(n399) );
  INV_X1 U512 ( .A(n406), .ZN(n402) );
  XNOR2_X2 U513 ( .A(n530), .B(n529), .ZN(n763) );
  AND2_X1 U514 ( .A1(n611), .A2(n610), .ZN(n407) );
  XOR2_X1 U515 ( .A(n417), .B(n416), .Z(n408) );
  XOR2_X1 U516 ( .A(G128), .B(G119), .Z(n409) );
  XNOR2_X1 U517 ( .A(n615), .B(KEYINPUT48), .ZN(n616) );
  INV_X1 U518 ( .A(G104), .ZN(n479) );
  XNOR2_X1 U519 ( .A(n490), .B(KEYINPUT5), .ZN(n491) );
  INV_X1 U520 ( .A(n587), .ZN(n588) );
  XNOR2_X1 U521 ( .A(n492), .B(n491), .ZN(n496) );
  INV_X1 U522 ( .A(G478), .ZN(n431) );
  XNOR2_X1 U523 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U524 ( .A(n418), .B(n408), .ZN(n419) );
  INV_X1 U525 ( .A(KEYINPUT63), .ZN(n640) );
  NAND2_X1 U526 ( .A1(G214), .A2(n487), .ZN(n412) );
  XNOR2_X1 U527 ( .A(n415), .B(n414), .ZN(n420) );
  XNOR2_X1 U528 ( .A(n452), .B(KEYINPUT104), .ZN(n418) );
  XOR2_X1 U529 ( .A(KEYINPUT103), .B(KEYINPUT12), .Z(n417) );
  XNOR2_X1 U530 ( .A(G140), .B(KEYINPUT11), .ZN(n416) );
  INV_X1 U531 ( .A(G902), .ZN(n512) );
  NAND2_X1 U532 ( .A1(n646), .A2(n512), .ZN(n422) );
  XOR2_X1 U533 ( .A(KEYINPUT13), .B(G475), .Z(n421) );
  XNOR2_X1 U534 ( .A(n422), .B(n421), .ZN(n550) );
  XOR2_X1 U535 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n424) );
  NAND2_X1 U536 ( .A1(G234), .A2(n755), .ZN(n423) );
  NAND2_X1 U537 ( .A1(G217), .A2(n507), .ZN(n430) );
  XNOR2_X1 U538 ( .A(G134), .B(KEYINPUT9), .ZN(n428) );
  XNOR2_X1 U539 ( .A(G122), .B(G116), .ZN(n425) );
  XNOR2_X1 U540 ( .A(n425), .B(G107), .ZN(n449) );
  XNOR2_X1 U541 ( .A(n439), .B(KEYINPUT7), .ZN(n426) );
  XNOR2_X1 U542 ( .A(n449), .B(n426), .ZN(n427) );
  XNOR2_X1 U543 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U544 ( .A(n430), .B(n429), .ZN(n737) );
  NOR2_X1 U545 ( .A1(G902), .A2(n737), .ZN(n433) );
  INV_X1 U546 ( .A(n547), .ZN(n551) );
  XNOR2_X1 U547 ( .A(G902), .B(KEYINPUT15), .ZN(n456) );
  NAND2_X1 U548 ( .A1(G234), .A2(n456), .ZN(n434) );
  XNOR2_X1 U549 ( .A(KEYINPUT20), .B(n434), .ZN(n513) );
  AND2_X1 U550 ( .A1(n513), .A2(G221), .ZN(n435) );
  XNOR2_X1 U551 ( .A(n435), .B(KEYINPUT21), .ZN(n704) );
  INV_X1 U552 ( .A(n704), .ZN(n522) );
  NOR2_X1 U553 ( .A1(n691), .A2(n522), .ZN(n472) );
  NAND2_X1 U554 ( .A1(n463), .A2(G224), .ZN(n436) );
  XNOR2_X1 U555 ( .A(n436), .B(KEYINPUT82), .ZN(n438) );
  XNOR2_X1 U556 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U557 ( .A(n440), .B(n476), .ZN(n446) );
  XNOR2_X1 U558 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U559 ( .A(n443), .B(G101), .ZN(n475) );
  XNOR2_X1 U560 ( .A(n444), .B(n475), .ZN(n445) );
  XNOR2_X1 U561 ( .A(n446), .B(n445), .ZN(n455) );
  XNOR2_X1 U562 ( .A(n447), .B(G110), .ZN(n448) );
  XNOR2_X1 U563 ( .A(n449), .B(n448), .ZN(n454) );
  XNOR2_X1 U564 ( .A(n450), .B(G119), .ZN(n490) );
  INV_X1 U565 ( .A(n490), .ZN(n451) );
  XNOR2_X1 U566 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U567 ( .A(n454), .B(n453), .ZN(n747) );
  XNOR2_X1 U568 ( .A(n455), .B(n747), .ZN(n656) );
  INV_X1 U569 ( .A(n456), .ZN(n627) );
  NAND2_X1 U570 ( .A1(n512), .A2(n457), .ZN(n459) );
  NAND2_X1 U571 ( .A1(n459), .A2(G210), .ZN(n458) );
  NAND2_X1 U572 ( .A1(n459), .A2(G214), .ZN(n688) );
  INV_X1 U573 ( .A(n688), .ZN(n460) );
  XNOR2_X1 U574 ( .A(n461), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U575 ( .A1(n465), .A2(G902), .ZN(n462) );
  XOR2_X1 U576 ( .A(KEYINPUT97), .B(n462), .Z(n569) );
  INV_X1 U577 ( .A(n569), .ZN(n464) );
  NOR2_X1 U578 ( .A1(G898), .A2(n755), .ZN(n748) );
  NAND2_X1 U579 ( .A1(n464), .A2(n748), .ZN(n468) );
  NAND2_X1 U580 ( .A1(G952), .A2(n465), .ZN(n719) );
  NOR2_X1 U581 ( .A1(G953), .A2(n719), .ZN(n467) );
  INV_X1 U582 ( .A(KEYINPUT96), .ZN(n466) );
  XNOR2_X1 U583 ( .A(n467), .B(n466), .ZN(n571) );
  NAND2_X1 U584 ( .A1(n468), .A2(n571), .ZN(n469) );
  NAND2_X1 U585 ( .A1(n670), .A2(n469), .ZN(n471) );
  INV_X1 U586 ( .A(KEYINPUT0), .ZN(n470) );
  NAND2_X1 U587 ( .A1(n472), .A2(n525), .ZN(n474) );
  INV_X1 U588 ( .A(KEYINPUT22), .ZN(n473) );
  XNOR2_X1 U589 ( .A(G146), .B(n475), .ZN(n477) );
  XNOR2_X1 U590 ( .A(G107), .B(G110), .ZN(n483) );
  NAND2_X1 U591 ( .A1(G227), .A2(n755), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U593 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U594 ( .A(KEYINPUT1), .ZN(n485) );
  INV_X1 U595 ( .A(KEYINPUT93), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n619), .B(n486), .ZN(n600) );
  NAND2_X1 U597 ( .A1(n487), .A2(G210), .ZN(n488) );
  XNOR2_X1 U598 ( .A(n489), .B(n488), .ZN(n492) );
  XNOR2_X1 U599 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U600 ( .A(n498), .B(n497), .ZN(n635) );
  XNOR2_X1 U601 ( .A(KEYINPUT101), .B(G472), .ZN(n587) );
  INV_X1 U602 ( .A(KEYINPUT108), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n499), .B(KEYINPUT6), .ZN(n500) );
  INV_X1 U604 ( .A(n501), .ZN(n502) );
  XOR2_X1 U605 ( .A(KEYINPUT23), .B(KEYINPUT74), .Z(n505) );
  XNOR2_X1 U606 ( .A(KEYINPUT98), .B(KEYINPUT81), .ZN(n504) );
  XNOR2_X1 U607 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U608 ( .A1(G221), .A2(n507), .ZN(n510) );
  XOR2_X1 U609 ( .A(KEYINPUT24), .B(G110), .Z(n508) );
  XNOR2_X1 U610 ( .A(n508), .B(n409), .ZN(n509) );
  XNOR2_X1 U611 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U612 ( .A1(n651), .A2(n512), .ZN(n517) );
  XOR2_X1 U613 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n515) );
  AND2_X1 U614 ( .A1(n513), .A2(G217), .ZN(n514) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X2 U616 ( .A(n517), .B(n516), .ZN(n584) );
  NAND2_X1 U617 ( .A1(n597), .A2(n554), .ZN(n518) );
  XNOR2_X1 U618 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n519) );
  INV_X1 U619 ( .A(KEYINPUT90), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n521), .B(n520), .ZN(n562) );
  OR2_X2 U621 ( .A1(n562), .A2(KEYINPUT65), .ZN(n533) );
  NAND2_X1 U622 ( .A1(n701), .A2(n700), .ZN(n541) );
  XOR2_X1 U623 ( .A(KEYINPUT91), .B(KEYINPUT33), .Z(n523) );
  XNOR2_X1 U624 ( .A(KEYINPUT75), .B(n523), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n697), .A2(n540), .ZN(n527) );
  XOR2_X1 U626 ( .A(KEYINPUT76), .B(KEYINPUT34), .Z(n526) );
  XNOR2_X1 U627 ( .A(n527), .B(n526), .ZN(n528) );
  AND2_X1 U628 ( .A1(n550), .A2(n551), .ZN(n604) );
  NAND2_X1 U629 ( .A1(n528), .A2(n604), .ZN(n530) );
  INV_X1 U630 ( .A(KEYINPUT35), .ZN(n529) );
  NAND2_X1 U631 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U632 ( .A1(n763), .A2(n354), .ZN(n537) );
  NOR2_X1 U633 ( .A1(KEYINPUT65), .A2(KEYINPUT89), .ZN(n535) );
  INV_X1 U634 ( .A(KEYINPUT44), .ZN(n534) );
  AND2_X1 U635 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U636 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U637 ( .A1(n539), .A2(n538), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n763), .A2(KEYINPUT89), .ZN(n561) );
  INV_X1 U639 ( .A(n540), .ZN(n545) );
  OR2_X1 U640 ( .A1(n575), .A2(n541), .ZN(n710) );
  NOR2_X1 U641 ( .A1(n545), .A2(n710), .ZN(n543) );
  XNOR2_X1 U642 ( .A(KEYINPUT31), .B(KEYINPUT102), .ZN(n542) );
  XNOR2_X1 U643 ( .A(n543), .B(n542), .ZN(n682) );
  NAND2_X1 U644 ( .A1(n575), .A2(n701), .ZN(n544) );
  NOR2_X1 U645 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U646 ( .A1(n581), .A2(n546), .ZN(n665) );
  NAND2_X1 U647 ( .A1(n682), .A2(n665), .ZN(n553) );
  AND2_X1 U648 ( .A1(n547), .A2(n550), .ZN(n549) );
  INV_X1 U649 ( .A(KEYINPUT106), .ZN(n548) );
  INV_X1 U650 ( .A(n678), .ZN(n676) );
  INV_X1 U651 ( .A(n550), .ZN(n552) );
  NAND2_X1 U652 ( .A1(n552), .A2(n551), .ZN(n681) );
  XNOR2_X1 U653 ( .A(KEYINPUT107), .B(n681), .ZN(n625) );
  NOR2_X1 U654 ( .A1(n676), .A2(n625), .ZN(n693) );
  INV_X1 U655 ( .A(n693), .ZN(n603) );
  NAND2_X1 U656 ( .A1(n553), .A2(n603), .ZN(n559) );
  INV_X1 U657 ( .A(n554), .ZN(n705) );
  AND2_X1 U658 ( .A1(n619), .A2(n705), .ZN(n555) );
  AND2_X1 U659 ( .A1(n597), .A2(n555), .ZN(n556) );
  AND2_X1 U660 ( .A1(n557), .A2(n556), .ZN(n662) );
  INV_X1 U661 ( .A(n662), .ZN(n558) );
  AND2_X1 U662 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U663 ( .A1(n561), .A2(n560), .ZN(n564) );
  AND2_X1 U664 ( .A1(n354), .A2(KEYINPUT65), .ZN(n563) );
  NOR2_X1 U665 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U666 ( .A1(n566), .A2(n565), .ZN(n568) );
  INV_X1 U667 ( .A(KEYINPUT45), .ZN(n567) );
  XNOR2_X1 U668 ( .A(n568), .B(n567), .ZN(n630) );
  NOR2_X1 U669 ( .A1(G900), .A2(n569), .ZN(n570) );
  NAND2_X1 U670 ( .A1(n570), .A2(G953), .ZN(n572) );
  NAND2_X1 U671 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U672 ( .A1(n573), .A2(n704), .ZN(n582) );
  XOR2_X1 U673 ( .A(KEYINPUT73), .B(n582), .Z(n574) );
  NAND2_X1 U674 ( .A1(n574), .A2(n584), .ZN(n596) );
  XNOR2_X1 U675 ( .A(KEYINPUT28), .B(n576), .ZN(n577) );
  NAND2_X1 U676 ( .A1(n577), .A2(n581), .ZN(n669) );
  NAND2_X1 U677 ( .A1(n689), .A2(n688), .ZN(n692) );
  XOR2_X1 U678 ( .A(KEYINPUT41), .B(KEYINPUT113), .Z(n578) );
  XNOR2_X1 U679 ( .A(n579), .B(n578), .ZN(n713) );
  XNOR2_X1 U680 ( .A(n580), .B(KEYINPUT42), .ZN(n765) );
  INV_X1 U681 ( .A(KEYINPUT79), .ZN(n586) );
  NAND2_X1 U682 ( .A1(n699), .A2(n688), .ZN(n591) );
  XOR2_X1 U683 ( .A(KEYINPUT112), .B(KEYINPUT30), .Z(n590) );
  NOR2_X1 U684 ( .A1(n764), .A2(n765), .ZN(n595) );
  INV_X1 U685 ( .A(KEYINPUT46), .ZN(n594) );
  XNOR2_X1 U686 ( .A(n595), .B(n594), .ZN(n601) );
  NOR2_X1 U687 ( .A1(n601), .A2(n684), .ZN(n614) );
  INV_X1 U688 ( .A(n670), .ZN(n602) );
  INV_X1 U689 ( .A(n604), .ZN(n605) );
  NOR2_X1 U690 ( .A1(n605), .A2(n622), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n674) );
  NAND2_X1 U692 ( .A1(n608), .A2(n674), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(KEYINPUT84), .ZN(n612) );
  XNOR2_X1 U694 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n611) );
  NOR2_X1 U695 ( .A1(n612), .A2(n407), .ZN(n613) );
  XNOR2_X1 U696 ( .A(KEYINPUT72), .B(KEYINPUT88), .ZN(n615) );
  XOR2_X1 U697 ( .A(n618), .B(KEYINPUT110), .Z(n620) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n621), .B(KEYINPUT43), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n644) );
  NAND2_X1 U701 ( .A1(n624), .A2(n625), .ZN(n686) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n629), .A2(KEYINPUT2), .ZN(n631) );
  NOR2_X2 U704 ( .A1(n631), .A2(n741), .ZN(n724) );
  NOR2_X4 U705 ( .A1(n632), .A2(n724), .ZN(n733) );
  NAND2_X1 U706 ( .A1(n733), .A2(G472), .ZN(n637) );
  XOR2_X1 U707 ( .A(KEYINPUT92), .B(KEYINPUT114), .Z(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U711 ( .A(G952), .ZN(n638) );
  AND2_X1 U712 ( .A1(n638), .A2(G953), .ZN(n740) );
  NOR2_X2 U713 ( .A1(n639), .A2(n740), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G57) );
  XNOR2_X1 U715 ( .A(n642), .B(G119), .ZN(G21) );
  XOR2_X1 U716 ( .A(G140), .B(KEYINPUT117), .Z(n643) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(G42) );
  XNOR2_X1 U718 ( .A(n645), .B(G110), .ZN(G12) );
  NAND2_X1 U719 ( .A1(n733), .A2(G475), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT59), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X2 U722 ( .A1(n649), .A2(n740), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U724 ( .A1(n733), .A2(G217), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT125), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n654), .A2(n740), .ZN(G66) );
  NAND2_X1 U728 ( .A1(n733), .A2(G210), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X2 U732 ( .A1(n659), .A2(n740), .ZN(n661) );
  XOR2_X1 U733 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(G51) );
  XOR2_X1 U735 ( .A(G101), .B(n662), .Z(G3) );
  NOR2_X1 U736 ( .A1(n678), .A2(n665), .ZN(n664) );
  XNOR2_X1 U737 ( .A(G104), .B(KEYINPUT115), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n664), .B(n663), .ZN(G6) );
  NOR2_X1 U739 ( .A1(n681), .A2(n665), .ZN(n667) );
  XNOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U742 ( .A(G107), .B(n668), .ZN(G9) );
  XOR2_X1 U743 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NOR2_X1 U744 ( .A1(n669), .A2(n681), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n671), .A2(n353), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G30) );
  XNOR2_X1 U747 ( .A(G143), .B(n674), .ZN(G45) );
  NAND2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U749 ( .A(G146), .B(n677), .ZN(G48) );
  NOR2_X1 U750 ( .A1(n678), .A2(n682), .ZN(n679) );
  XOR2_X1 U751 ( .A(KEYINPUT116), .B(n679), .Z(n680) );
  XNOR2_X1 U752 ( .A(G113), .B(n680), .ZN(G15) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U754 ( .A(G116), .B(n683), .Z(G18) );
  XNOR2_X1 U755 ( .A(G125), .B(n684), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n685), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U757 ( .A(G134), .B(n686), .ZN(G36) );
  XOR2_X1 U758 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n729) );
  INV_X1 U759 ( .A(n697), .ZN(n687) );
  NOR2_X1 U760 ( .A1(n713), .A2(n687), .ZN(n722) );
  NOR2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U765 ( .A(KEYINPUT119), .B(n696), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n702), .B(KEYINPUT50), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n699), .A2(n703), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U771 ( .A(n706), .B(KEYINPUT49), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U774 ( .A(KEYINPUT51), .B(n711), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(n714), .Z(n715) );
  NAND2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U778 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n717) );
  XNOR2_X1 U779 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U781 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U782 ( .A(KEYINPUT121), .B(n723), .ZN(n727) );
  NOR2_X1 U783 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(G75) );
  XNOR2_X1 U785 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n730), .B(KEYINPUT57), .ZN(n731) );
  XNOR2_X1 U787 ( .A(n732), .B(n731), .ZN(n735) );
  NAND2_X1 U788 ( .A1(n733), .A2(G469), .ZN(n734) );
  XOR2_X1 U789 ( .A(n735), .B(n734), .Z(n736) );
  NOR2_X1 U790 ( .A1(n740), .A2(n736), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n733), .A2(G478), .ZN(n738) );
  XNOR2_X1 U792 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(G63) );
  NOR2_X1 U794 ( .A1(n741), .A2(G953), .ZN(n746) );
  NAND2_X1 U795 ( .A1(G224), .A2(G953), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(KEYINPUT126), .ZN(n743) );
  XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  AND2_X1 U798 ( .A1(n744), .A2(G898), .ZN(n745) );
  NOR2_X1 U799 ( .A1(n746), .A2(n745), .ZN(n751) );
  XOR2_X1 U800 ( .A(G101), .B(n747), .Z(n749) );
  NOR2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U802 ( .A(n751), .B(n750), .Z(G69) );
  XOR2_X1 U803 ( .A(n753), .B(n752), .Z(n757) );
  XNOR2_X1 U804 ( .A(n754), .B(n757), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n761) );
  XNOR2_X1 U806 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U810 ( .A(KEYINPUT127), .B(n762), .Z(G72) );
  XNOR2_X1 U811 ( .A(n763), .B(G122), .ZN(G24) );
  XOR2_X1 U812 ( .A(n764), .B(G131), .Z(G33) );
  XOR2_X1 U813 ( .A(n765), .B(G137), .Z(G39) );
endmodule

