//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT66), .B1(new_n203), .B2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(new_n206), .A3(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(G113gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT67), .A4(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G127gat), .B(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n206), .A2(G120gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n208), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n214), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  INV_X1    g023(.A(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227));
  NOR3_X1   g026(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(KEYINPUT73), .A3(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT73), .B1(new_n226), .B2(new_n227), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT71), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(G155gat), .B2(G162gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n230), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  OAI22_X1  g040(.A1(new_n234), .A2(new_n235), .B1(new_n241), .B2(KEYINPUT72), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(KEYINPUT72), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n223), .B(new_n231), .C1(new_n242), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n239), .A2(G155gat), .A3(G162gat), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT71), .B1(new_n236), .B2(new_n237), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n229), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT73), .ZN(new_n252));
  INV_X1    g051(.A(new_n227), .ZN(new_n253));
  NOR2_X1   g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n232), .A3(new_n233), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n243), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n223), .B1(new_n257), .B2(new_n231), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n246), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n231), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(KEYINPUT74), .A3(new_n222), .A4(new_n245), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n222), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n220), .B1(new_n213), .B2(new_n216), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n231), .A4(new_n257), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n263), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n222), .A2(new_n260), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n231), .A3(new_n257), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n266), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277));
  OR3_X1    g076(.A1(new_n276), .A2(new_n277), .A3(new_n270), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n276), .B2(new_n270), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n272), .B1(new_n263), .B2(new_n269), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n271), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G1gat), .B(G29gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT0), .ZN(new_n284));
  XNOR2_X1  g083(.A(G57gat), .B(G85gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT77), .B1(new_n282), .B2(new_n287), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n286), .B(new_n271), .C1(new_n280), .C2(new_n281), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n289), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n282), .A2(KEYINPUT77), .A3(new_n287), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n290), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n298));
  XOR2_X1   g097(.A(G8gat), .B(G36gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT70), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(G211gat), .ZN(new_n304));
  INV_X1    g103(.A(G218gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(KEYINPUT22), .B2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G211gat), .B(G218gat), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT25), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(KEYINPUT24), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(G169gat), .ZN(new_n320));
  INV_X1    g119(.A(G176gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G183gat), .ZN(new_n325));
  INV_X1    g124(.A(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT24), .A3(new_n316), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n318), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n318), .A2(new_n324), .A3(new_n328), .A4(new_n330), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n314), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT27), .B(G183gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n326), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n325), .A2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G183gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n340), .A3(new_n326), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT65), .A3(KEYINPUT28), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n337), .A2(new_n342), .A3(new_n316), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n311), .B1(new_n334), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n314), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n317), .B1(new_n323), .B2(new_n322), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n330), .B1(new_n352), .B2(new_n328), .ZN(new_n353));
  AND4_X1   g152(.A1(new_n330), .A2(new_n318), .A3(new_n324), .A4(new_n328), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n355), .B2(new_n348), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n309), .B(new_n350), .C1(new_n356), .C2(new_n311), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n310), .B1(new_n355), .B2(new_n348), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT68), .B(KEYINPUT29), .Z(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n334), .B2(new_n349), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n310), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n302), .B(new_n357), .C1(new_n361), .C2(new_n309), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n359), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n355), .B2(new_n348), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n350), .B1(new_n366), .B2(new_n311), .ZN(new_n367));
  INV_X1    g166(.A(new_n309), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n302), .A4(new_n357), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n357), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(new_n310), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n309), .B1(new_n373), .B2(new_n350), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT69), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n357), .C1(new_n361), .C2(new_n309), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n302), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n298), .B1(new_n297), .B2(new_n380), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n295), .A2(new_n291), .A3(new_n293), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT78), .B(new_n379), .C1(new_n382), .C2(new_n290), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n222), .A2(new_n355), .A3(new_n348), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n267), .B1(new_n334), .B2(new_n349), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G227gat), .ZN(new_n387));
  INV_X1    g186(.A(G233gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n391));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n387), .A2(new_n388), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n384), .A2(new_n385), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n390), .A2(new_n391), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n390), .B2(new_n391), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(KEYINPUT32), .A3(new_n396), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n245), .A2(new_n359), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n368), .ZN(new_n408));
  INV_X1    g207(.A(new_n260), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n309), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(G228gat), .A3(G233gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n309), .B2(new_n359), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n408), .B(new_n414), .C1(new_n409), .C2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT31), .B(G50gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n413), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n413), .B2(new_n416), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G22gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OR3_X1    g222(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n406), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n381), .A2(new_n383), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n429));
  AND4_X1   g228(.A1(KEYINPUT82), .A2(new_n282), .A3(KEYINPUT6), .A4(new_n287), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n263), .A2(new_n269), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT75), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n432), .A2(new_n273), .A3(new_n279), .A4(new_n278), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n286), .B1(new_n433), .B2(new_n271), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT82), .B1(new_n434), .B2(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n302), .ZN(new_n438));
  INV_X1    g237(.A(new_n377), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n376), .B1(new_n369), .B2(new_n357), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(KEYINPUT79), .A3(new_n364), .A4(new_n370), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n371), .B2(new_n378), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n406), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n426), .A2(KEYINPUT35), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n381), .A2(new_n383), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n426), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n265), .A2(new_n268), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n266), .B1(new_n263), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n274), .A2(new_n266), .A3(new_n275), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(KEYINPUT39), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n452), .B1(new_n259), .B2(new_n262), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n266), .ZN(new_n460));
  AND4_X1   g259(.A1(KEYINPUT40), .A2(new_n456), .A3(new_n460), .A4(new_n286), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n287), .B1(new_n454), .B2(new_n455), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT40), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n434), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n426), .B1(new_n464), .B2(new_n445), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n369), .A2(new_n466), .A3(new_n357), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n369), .A2(KEYINPUT80), .A3(new_n466), .A4(new_n357), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n302), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT37), .B1(new_n439), .B2(new_n440), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT38), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n466), .B1(new_n367), .B2(new_n309), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n368), .B(new_n350), .C1(new_n356), .C2(new_n311), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT38), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n471), .A2(KEYINPUT81), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT81), .B1(new_n471), .B2(new_n477), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n474), .B(new_n362), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n465), .B1(new_n437), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n406), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n451), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n449), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G29gat), .A2(G36gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT84), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n492), .A2(new_n497), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n491), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n486), .A2(new_n487), .ZN(new_n501));
  NOR4_X1   g300(.A1(new_n500), .A2(new_n501), .A3(new_n488), .A4(new_n494), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT16), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(G1gat), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  OAI221_X1 g306(.A(new_n506), .B1(KEYINPUT86), .B2(new_n507), .C1(G1gat), .C2(new_n504), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n503), .A2(new_n510), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT87), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT13), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G197gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT11), .B(G169gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n522), .B(new_n523), .Z(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT12), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT18), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n512), .B(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n510), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n518), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n529), .A2(KEYINPUT18), .A3(new_n518), .A4(new_n532), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n520), .A2(new_n526), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n519), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n513), .B(KEYINPUT88), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(new_n511), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n536), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n525), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT89), .B1(new_n485), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n448), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n545), .B1(new_n428), .B2(KEYINPUT35), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n481), .A2(new_n483), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n450), .B2(new_n426), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT89), .B(new_n543), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  INV_X1    g354(.A(G85gat), .ZN(new_n556));
  INV_X1    g355(.A(G92gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(KEYINPUT8), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G99gat), .B(G106gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n552), .B1(new_n503), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n530), .A2(new_n531), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G134gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(new_n237), .ZN(new_n572));
  INV_X1    g371(.A(new_n568), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n565), .B2(new_n566), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n581), .A2(new_n585), .B1(new_n586), .B2(KEYINPUT90), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(KEYINPUT90), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G127gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n510), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT91), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n594), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n598), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n589), .B(new_n561), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(KEYINPUT10), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n561), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT94), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n609), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(KEYINPUT95), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(KEYINPUT95), .ZN(new_n623));
  NOR4_X1   g422(.A1(new_n615), .A2(new_n619), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n621), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n619), .B1(new_n611), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n580), .A2(new_n604), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n551), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n297), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g433(.A(new_n445), .B1(new_n631), .B2(new_n632), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT16), .B(G8gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n635), .B2(G8gat), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n639), .A2(new_n641), .B1(new_n636), .B2(new_n645), .ZN(G1325gat));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n632), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n647), .A2(G15gat), .A3(new_n406), .ZN(new_n648));
  OAI21_X1  g447(.A(G15gat), .B1(new_n647), .B2(new_n483), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(G1326gat));
  OAI21_X1  g449(.A(new_n426), .B1(new_n631), .B2(new_n632), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT43), .B(G22gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  NOR2_X1   g452(.A1(new_n544), .A2(new_n550), .ZN(new_n654));
  INV_X1    g453(.A(new_n297), .ZN(new_n655));
  INV_X1    g454(.A(new_n628), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n604), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n579), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n654), .A2(G29gat), .A3(new_n655), .A4(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT45), .Z(new_n661));
  NAND3_X1  g460(.A1(new_n484), .A2(new_n449), .A3(KEYINPUT101), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n546), .B2(new_n548), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n579), .A2(KEYINPUT44), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n580), .B1(new_n546), .B2(new_n548), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT44), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n667), .B2(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n543), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n537), .A2(new_n542), .A3(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n657), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n655), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n679), .ZN(G1328gat));
  INV_X1    g479(.A(new_n445), .ZN(new_n681));
  NOR4_X1   g480(.A1(new_n654), .A2(G36gat), .A3(new_n681), .A4(new_n659), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT46), .ZN(new_n683));
  OAI21_X1  g482(.A(G36gat), .B1(new_n678), .B2(new_n681), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(new_n483), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n686), .A3(new_n677), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G43gat), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n687), .A2(KEYINPUT102), .A3(G43gat), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n406), .A2(G43gat), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n551), .A2(KEYINPUT103), .A3(new_n658), .A4(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n658), .B(new_n692), .C1(new_n544), .C2(new_n550), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT47), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n690), .A2(new_n691), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n688), .A2(new_n694), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT47), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n698), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(G1330gat));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n654), .A2(new_n659), .ZN(new_n706));
  INV_X1    g505(.A(new_n426), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(G50gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT105), .Z(new_n710));
  NAND3_X1  g509(.A1(new_n671), .A2(new_n426), .A3(new_n677), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n705), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT48), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT106), .B1(new_n706), .B2(new_n708), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n715), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n717), .ZN(G1331gat));
  AND2_X1   g517(.A1(new_n662), .A2(new_n664), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n675), .A2(new_n580), .A3(new_n604), .A4(new_n656), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n655), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT107), .B(G57gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n681), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n721), .B2(new_n483), .ZN(new_n730));
  INV_X1    g529(.A(new_n406), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n583), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n721), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n721), .A2(new_n707), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n584), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n675), .A2(new_n603), .A3(new_n656), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n671), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n671), .A2(KEYINPUT109), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743), .B2(new_n655), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n485), .A2(new_n580), .A3(new_n604), .A4(new_n676), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(KEYINPUT110), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n746), .A2(KEYINPUT110), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n656), .B1(new_n745), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n556), .A3(new_n297), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n744), .A2(new_n753), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n557), .A3(new_n445), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g555(.A(G92gat), .B1(new_n739), .B2(new_n681), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n445), .A3(new_n742), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n755), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(new_n756), .ZN(G1337gat));
  AOI21_X1  g561(.A(G99gat), .B1(new_n752), .B2(new_n731), .ZN(new_n763));
  INV_X1    g562(.A(new_n743), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n686), .A2(G99gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(G1338gat));
  OR3_X1    g565(.A1(new_n751), .A2(G106gat), .A3(new_n707), .ZN(new_n767));
  OAI21_X1  g566(.A(G106gat), .B1(new_n739), .B2(new_n707), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n741), .A2(new_n426), .A3(new_n742), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n767), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(G1339gat));
  NAND3_X1  g574(.A1(new_n297), .A2(new_n446), .A3(new_n707), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n777));
  AOI21_X1  g576(.A(new_n618), .B1(new_n611), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT54), .B1(new_n608), .B2(new_n609), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n615), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n780), .A2(KEYINPUT114), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT114), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n624), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n781), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT115), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n537), .A2(new_n542), .A3(KEYINPUT99), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT99), .B1(new_n537), .B2(new_n542), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n784), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n533), .A2(new_n534), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n517), .B2(new_n519), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n524), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n628), .A2(new_n792), .A3(new_n537), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n580), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n784), .A2(new_n786), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n792), .A2(new_n537), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n795), .A2(new_n580), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n795), .A2(new_n537), .A3(new_n580), .A4(new_n792), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  INV_X1    g599(.A(new_n793), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n675), .B2(new_n795), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n580), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n803), .A3(new_n604), .ZN(new_n804));
  INV_X1    g603(.A(new_n629), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT112), .B1(new_n805), .B2(new_n675), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n676), .A2(new_n807), .A3(new_n629), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n776), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n675), .ZN(new_n812));
  INV_X1    g611(.A(new_n543), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n206), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n811), .B2(new_n814), .ZN(G1340gat));
  NOR2_X1   g614(.A1(KEYINPUT117), .A2(G120gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n811), .B2(new_n628), .ZN(new_n817));
  NAND2_X1  g616(.A1(KEYINPUT117), .A2(G120gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT118), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n817), .B(new_n819), .ZN(G1341gat));
  AND3_X1   g619(.A1(new_n811), .A2(G127gat), .A3(new_n603), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(KEYINPUT119), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(KEYINPUT119), .ZN(new_n823));
  AOI21_X1  g622(.A(G127gat), .B1(new_n811), .B2(new_n603), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n826), .A3(new_n580), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT120), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n811), .B2(new_n580), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(KEYINPUT56), .B2(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1343gat));
  NOR2_X1   g631(.A1(new_n655), .A2(new_n445), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n686), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n804), .A2(new_n810), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(new_n837), .B2(new_n426), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n707), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n784), .A2(new_n543), .A3(new_n785), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n580), .B1(new_n842), .B2(new_n793), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n603), .B1(new_n844), .B2(new_n799), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n809), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT121), .B(new_n841), .C1(new_n809), .C2(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n836), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n224), .B1(new_n852), .B2(new_n543), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n707), .B(new_n836), .C1(new_n804), .C2(new_n810), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n813), .A2(G141gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n675), .B(new_n835), .C1(new_n838), .C2(new_n850), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n859), .A2(G141gat), .B1(new_n854), .B2(new_n855), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n853), .A2(new_n858), .B1(new_n860), .B2(new_n857), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n854), .A2(new_n225), .A3(new_n628), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G148gat), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n852), .B2(new_n628), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n834), .A2(new_n656), .ZN(new_n866));
  INV_X1    g665(.A(new_n841), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n804), .B2(new_n810), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n604), .B1(new_n797), .B2(new_n843), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n543), .B2(new_n805), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n426), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n483), .B(new_n866), .C1(new_n868), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n863), .B1(new_n872), .B2(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n862), .B1(new_n865), .B2(new_n873), .ZN(G1345gat));
  NAND3_X1  g673(.A1(new_n854), .A2(new_n236), .A3(new_n603), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n852), .A2(new_n603), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n236), .ZN(G1346gat));
  NAND3_X1  g676(.A1(new_n854), .A2(new_n237), .A3(new_n580), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n852), .A2(new_n580), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n237), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n297), .A2(new_n681), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n837), .A2(new_n427), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n675), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n813), .A2(new_n320), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(G1348gat));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n628), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(G176gat), .ZN(G1349gat));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n336), .B1(new_n888), .B2(G183gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n882), .A2(new_n603), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n882), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n604), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n888), .A2(new_n325), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT60), .B(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895));
  INV_X1    g694(.A(new_n890), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n882), .B2(new_n603), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n894), .A2(new_n898), .ZN(G1350gat));
  OAI22_X1  g698(.A1(new_n891), .A2(new_n579), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(G1351gat));
  NOR2_X1   g701(.A1(new_n686), .A2(new_n707), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n837), .A2(new_n881), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n837), .A2(KEYINPUT123), .A3(new_n881), .A4(new_n903), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n676), .A2(G197gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n483), .B(new_n881), .C1(new_n868), .C2(new_n871), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n913), .B2(new_n813), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G197gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n913), .A2(KEYINPUT125), .A3(new_n813), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n911), .A2(new_n912), .B1(new_n915), .B2(new_n916), .ZN(G1352gat));
  OAI21_X1  g716(.A(G204gat), .B1(new_n913), .B2(new_n656), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n656), .A2(G204gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n837), .A2(new_n881), .A3(new_n903), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT126), .B1(new_n920), .B2(KEYINPUT62), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n920), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n922));
  OAI221_X1 g721(.A(new_n918), .B1(KEYINPUT62), .B2(new_n920), .C1(new_n921), .C2(new_n922), .ZN(G1353gat));
  NAND4_X1  g722(.A1(new_n906), .A2(new_n304), .A3(new_n603), .A4(new_n907), .ZN(new_n924));
  OAI21_X1  g723(.A(G211gat), .B1(new_n913), .B2(new_n604), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g726(.A(KEYINPUT63), .B(G211gat), .C1(new_n913), .C2(new_n604), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n927), .B2(new_n929), .ZN(G1354gat));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n580), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n913), .A2(new_n931), .ZN(new_n934));
  OAI21_X1  g733(.A(G218gat), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n906), .A2(new_n305), .A3(new_n580), .A4(new_n907), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1355gat));
endmodule


