

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794;

  XNOR2_X1 U371 ( .A(n733), .B(KEYINPUT62), .ZN(n734) );
  XNOR2_X1 U372 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U373 ( .A(n718), .B(KEYINPUT59), .ZN(n719) );
  BUF_X1 U374 ( .A(n654), .Z(n739) );
  INV_X1 U375 ( .A(n614), .ZN(n348) );
  XNOR2_X1 U376 ( .A(n607), .B(KEYINPUT108), .ZN(n436) );
  BUF_X1 U377 ( .A(n623), .Z(n624) );
  XNOR2_X1 U378 ( .A(G113), .B(G143), .ZN(n473) );
  XOR2_X1 U379 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n531) );
  XNOR2_X1 U380 ( .A(KEYINPUT16), .B(G122), .ZN(n492) );
  XNOR2_X1 U381 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n543) );
  XNOR2_X1 U382 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n495) );
  INV_X2 U383 ( .A(G128), .ZN(n460) );
  AND2_X4 U384 ( .A1(G902), .A2(G469), .ZN(n399) );
  NAND2_X2 U385 ( .A1(n624), .A2(n669), .ZN(n591) );
  XNOR2_X2 U386 ( .A(n349), .B(n348), .ZN(n630) );
  NAND2_X2 U387 ( .A1(n360), .A2(n612), .ZN(n349) );
  XNOR2_X2 U388 ( .A(n550), .B(n549), .ZN(n659) );
  NAND2_X1 U389 ( .A1(G234), .A2(G237), .ZN(n506) );
  XNOR2_X1 U390 ( .A(G146), .B(G137), .ZN(n533) );
  XOR2_X1 U391 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n530) );
  XOR2_X1 U392 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n476) );
  XNOR2_X1 U393 ( .A(G101), .B(G146), .ZN(n523) );
  INV_X1 U394 ( .A(G237), .ZN(n502) );
  XNOR2_X1 U395 ( .A(KEYINPUT3), .B(G119), .ZN(n490) );
  XNOR2_X1 U396 ( .A(KEYINPUT74), .B(KEYINPUT8), .ZN(n435) );
  INV_X1 U397 ( .A(G902), .ZN(n427) );
  XOR2_X1 U398 ( .A(n611), .B(KEYINPUT67), .Z(n350) );
  AND2_X1 U399 ( .A1(n638), .A2(n673), .ZN(n351) );
  AND2_X2 U400 ( .A1(n752), .A2(G469), .ZN(n405) );
  XNOR2_X2 U401 ( .A(n782), .B(n527), .ZN(n752) );
  AND2_X2 U402 ( .A1(n364), .A2(n379), .ZN(n363) );
  NAND2_X1 U403 ( .A1(n571), .A2(n570), .ZN(n601) );
  AND2_X1 U404 ( .A1(n370), .A2(n368), .ZN(n379) );
  INV_X1 U405 ( .A(n603), .ZN(n414) );
  NAND2_X1 U406 ( .A1(n374), .A2(n371), .ZN(n794) );
  INV_X1 U407 ( .A(n780), .ZN(n384) );
  NOR2_X1 U408 ( .A1(n649), .A2(KEYINPUT79), .ZN(n385) );
  AND2_X1 U409 ( .A1(n351), .A2(n377), .ZN(n372) );
  INV_X1 U410 ( .A(n570), .ZN(n578) );
  NOR2_X1 U411 ( .A1(n633), .A2(n563), .ZN(n404) );
  XNOR2_X1 U412 ( .A(n504), .B(n503), .ZN(n633) );
  XNOR2_X1 U413 ( .A(n747), .B(n390), .ZN(n726) );
  XNOR2_X1 U414 ( .A(n537), .B(n391), .ZN(n747) );
  XNOR2_X1 U415 ( .A(n392), .B(n490), .ZN(n537) );
  XNOR2_X1 U416 ( .A(n491), .B(G104), .ZN(n525) );
  XNOR2_X1 U417 ( .A(G146), .B(G125), .ZN(n498) );
  XNOR2_X1 U418 ( .A(G110), .B(G107), .ZN(n491) );
  INV_X1 U419 ( .A(KEYINPUT32), .ZN(n377) );
  INV_X8 U420 ( .A(G953), .ZN(n786) );
  INV_X1 U421 ( .A(KEYINPUT79), .ZN(n381) );
  INV_X1 U422 ( .A(KEYINPUT4), .ZN(n493) );
  NAND2_X1 U423 ( .A1(n362), .A2(n395), .ZN(n361) );
  NAND2_X1 U424 ( .A1(n382), .A2(n381), .ZN(n358) );
  AND2_X1 U425 ( .A1(n413), .A2(n416), .ZN(n395) );
  NAND2_X1 U426 ( .A1(n414), .A2(KEYINPUT44), .ZN(n413) );
  AND2_X1 U427 ( .A1(n415), .A2(KEYINPUT82), .ZN(n394) );
  OR2_X1 U428 ( .A1(n599), .A2(KEYINPUT83), .ZN(n409) );
  NOR2_X1 U429 ( .A1(n604), .A2(KEYINPUT44), .ZN(n369) );
  AND2_X1 U430 ( .A1(n440), .A2(KEYINPUT48), .ZN(n439) );
  XNOR2_X1 U431 ( .A(n393), .B(KEYINPUT85), .ZN(n603) );
  NAND2_X1 U432 ( .A1(n794), .A2(n602), .ZN(n393) );
  NOR2_X1 U433 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U434 ( .A1(n629), .A2(n451), .ZN(n449) );
  AND2_X1 U435 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U436 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U437 ( .A1(n649), .A2(KEYINPUT79), .ZN(n387) );
  XNOR2_X1 U438 ( .A(n356), .B(KEYINPUT109), .ZN(n355) );
  AND2_X1 U439 ( .A1(n610), .A2(n688), .ZN(n354) );
  AND2_X1 U440 ( .A1(n610), .A2(n631), .ZN(n357) );
  NOR2_X1 U441 ( .A1(n690), .A2(n693), .ZN(n615) );
  XNOR2_X1 U442 ( .A(n431), .B(n430), .ZN(n669) );
  BUF_X1 U443 ( .A(n576), .Z(n673) );
  INV_X1 U444 ( .A(n776), .ZN(n352) );
  OR2_X1 U445 ( .A1(n552), .A2(n551), .ZN(n553) );
  AND2_X1 U446 ( .A1(KEYINPUT82), .A2(KEYINPUT44), .ZN(n367) );
  XNOR2_X1 U447 ( .A(n525), .B(n492), .ZN(n391) );
  NOR2_X1 U448 ( .A1(n434), .A2(G953), .ZN(n433) );
  XNOR2_X1 U449 ( .A(n498), .B(KEYINPUT10), .ZN(n784) );
  INV_X1 U450 ( .A(G234), .ZN(n434) );
  XNOR2_X1 U451 ( .A(G116), .B(G134), .ZN(n463) );
  XNOR2_X2 U452 ( .A(G902), .B(KEYINPUT15), .ZN(n651) );
  XNOR2_X1 U453 ( .A(G107), .B(KEYINPUT104), .ZN(n464) );
  XNOR2_X1 U454 ( .A(G116), .B(G113), .ZN(n489) );
  XNOR2_X1 U455 ( .A(G134), .B(G131), .ZN(n519) );
  NOR2_X2 U456 ( .A1(G953), .A2(G237), .ZN(n532) );
  XOR2_X2 U457 ( .A(G104), .B(G122), .Z(n474) );
  XNOR2_X1 U458 ( .A(KEYINPUT101), .B(KEYINPUT12), .ZN(n475) );
  XNOR2_X2 U459 ( .A(G128), .B(KEYINPUT24), .ZN(n545) );
  XOR2_X1 U460 ( .A(G140), .B(G131), .Z(n480) );
  XNOR2_X2 U461 ( .A(G119), .B(G110), .ZN(n546) );
  XNOR2_X2 U462 ( .A(G140), .B(G137), .ZN(n544) );
  XOR2_X1 U463 ( .A(KEYINPUT91), .B(KEYINPUT89), .Z(n496) );
  XNOR2_X2 U464 ( .A(n353), .B(n350), .ZN(n360) );
  NAND2_X1 U465 ( .A1(n436), .A2(n354), .ZN(n353) );
  NAND2_X1 U466 ( .A1(n355), .A2(n632), .ZN(n769) );
  NAND2_X1 U467 ( .A1(n436), .A2(n357), .ZN(n356) );
  XNOR2_X1 U468 ( .A(n785), .B(KEYINPUT71), .ZN(n650) );
  XNOR2_X2 U469 ( .A(n655), .B(KEYINPUT78), .ZN(n785) );
  NAND2_X2 U470 ( .A1(n359), .A2(n358), .ZN(n655) );
  AND2_X2 U471 ( .A1(n386), .A2(n383), .ZN(n359) );
  NAND2_X1 U472 ( .A1(n360), .A2(n352), .ZN(n780) );
  NAND2_X1 U473 ( .A1(n363), .A2(n361), .ZN(n378) );
  NAND2_X1 U474 ( .A1(n365), .A2(n415), .ZN(n362) );
  NAND2_X1 U475 ( .A1(n365), .A2(n394), .ZN(n364) );
  NAND2_X1 U476 ( .A1(n412), .A2(n411), .ZN(n365) );
  NAND2_X1 U477 ( .A1(n515), .A2(n366), .ZN(n518) );
  NAND2_X1 U478 ( .A1(n680), .A2(n366), .ZN(n590) );
  NAND2_X1 U479 ( .A1(n593), .A2(n366), .ZN(n761) );
  NAND2_X1 U480 ( .A1(n685), .A2(n366), .ZN(n582) );
  XNOR2_X2 U481 ( .A(n389), .B(n514), .ZN(n366) );
  NAND2_X1 U482 ( .A1(n414), .A2(n367), .ZN(n370) );
  NAND2_X1 U483 ( .A1(n369), .A2(n603), .ZN(n368) );
  INV_X1 U484 ( .A(n601), .ZN(n373) );
  OR2_X1 U485 ( .A1(n351), .A2(n377), .ZN(n375) );
  NAND2_X1 U486 ( .A1(n601), .A2(KEYINPUT32), .ZN(n376) );
  XNOR2_X2 U487 ( .A(n378), .B(n605), .ZN(n654) );
  INV_X1 U488 ( .A(n388), .ZN(n382) );
  NAND2_X1 U489 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U490 ( .A1(n438), .A2(n398), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n639), .A2(n513), .ZN(n389) );
  XNOR2_X1 U492 ( .A(n404), .B(n403), .ZN(n639) );
  XNOR2_X1 U493 ( .A(n520), .B(n501), .ZN(n390) );
  XNOR2_X2 U494 ( .A(n494), .B(n493), .ZN(n520) );
  XNOR2_X1 U495 ( .A(n489), .B(n488), .ZN(n392) );
  XNOR2_X2 U496 ( .A(n623), .B(KEYINPUT1), .ZN(n577) );
  XNOR2_X2 U497 ( .A(n528), .B(n521), .ZN(n782) );
  XNOR2_X2 U498 ( .A(n520), .B(n519), .ZN(n528) );
  NAND2_X1 U499 ( .A1(n428), .A2(n427), .ZN(n426) );
  INV_X1 U500 ( .A(KEYINPUT84), .ZN(n585) );
  INV_X1 U501 ( .A(G221), .ZN(n458) );
  INV_X1 U502 ( .A(KEYINPUT34), .ZN(n454) );
  NAND2_X1 U503 ( .A1(n726), .A2(n651), .ZN(n504) );
  XNOR2_X1 U504 ( .A(n432), .B(n554), .ZN(n576) );
  XNOR2_X1 U505 ( .A(n435), .B(n433), .ZN(n541) );
  AND2_X1 U506 ( .A1(n446), .A2(n396), .ZN(n445) );
  NAND2_X1 U507 ( .A1(n793), .A2(KEYINPUT46), .ZN(n446) );
  INV_X1 U508 ( .A(KEYINPUT82), .ZN(n416) );
  INV_X1 U509 ( .A(G469), .ZN(n428) );
  INV_X1 U510 ( .A(KEYINPUT96), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n465) );
  NAND2_X1 U512 ( .A1(n423), .A2(KEYINPUT77), .ZN(n422) );
  NAND2_X1 U513 ( .A1(n651), .A2(n606), .ZN(n420) );
  AND2_X1 U514 ( .A1(n620), .A2(n687), .ZN(n608) );
  INV_X1 U515 ( .A(KEYINPUT65), .ZN(n430) );
  NOR2_X1 U516 ( .A1(n576), .A2(n672), .ZN(n431) );
  INV_X1 U517 ( .A(KEYINPUT75), .ZN(n406) );
  XNOR2_X1 U518 ( .A(n452), .B(n400), .ZN(n584) );
  NAND2_X1 U519 ( .A1(n453), .A2(n632), .ZN(n452) );
  INV_X1 U520 ( .A(KEYINPUT19), .ZN(n403) );
  OR2_X1 U521 ( .A1(n786), .A2(G952), .ZN(n736) );
  INV_X1 U522 ( .A(KEYINPUT81), .ZN(n572) );
  INV_X1 U523 ( .A(n629), .ZN(n447) );
  AND2_X1 U524 ( .A1(n769), .A2(n648), .ZN(n396) );
  OR2_X1 U525 ( .A1(n739), .A2(n785), .ZN(n397) );
  AND2_X1 U526 ( .A1(n437), .A2(n442), .ZN(n398) );
  XOR2_X1 U527 ( .A(KEYINPUT73), .B(KEYINPUT35), .Z(n400) );
  AND2_X1 U528 ( .A1(KEYINPUT46), .A2(n450), .ZN(n401) );
  INV_X1 U529 ( .A(KEYINPUT77), .ZN(n606) );
  INV_X1 U530 ( .A(KEYINPUT83), .ZN(n417) );
  INV_X1 U531 ( .A(KEYINPUT48), .ZN(n450) );
  BUF_X1 U532 ( .A(n633), .Z(n402) );
  NOR2_X1 U533 ( .A1(n405), .A2(n399), .ZN(n429) );
  NAND2_X1 U534 ( .A1(n407), .A2(n406), .ZN(n666) );
  NAND2_X1 U535 ( .A1(n397), .A2(n662), .ZN(n407) );
  NAND2_X1 U536 ( .A1(n439), .A2(n441), .ZN(n438) );
  XNOR2_X2 U537 ( .A(n591), .B(KEYINPUT97), .ZN(n607) );
  NAND2_X1 U538 ( .A1(n408), .A2(n650), .ZN(n424) );
  NOR2_X1 U539 ( .A1(n419), .A2(n421), .ZN(n408) );
  XNOR2_X1 U540 ( .A(n586), .B(n585), .ZN(n600) );
  NAND2_X2 U541 ( .A1(n429), .A2(n425), .ZN(n623) );
  XNOR2_X1 U542 ( .A(n582), .B(n454), .ZN(n453) );
  NAND2_X1 U543 ( .A1(n410), .A2(n409), .ZN(n412) );
  INV_X1 U544 ( .A(n600), .ZN(n410) );
  NAND2_X1 U545 ( .A1(n600), .A2(n417), .ZN(n411) );
  NAND2_X1 U546 ( .A1(n599), .A2(KEYINPUT83), .ZN(n415) );
  NAND2_X1 U547 ( .A1(n418), .A2(n420), .ZN(n419) );
  NAND2_X1 U548 ( .A1(n654), .A2(n606), .ZN(n418) );
  NOR2_X1 U549 ( .A1(n654), .A2(n422), .ZN(n421) );
  INV_X1 U550 ( .A(n651), .ZN(n423) );
  XNOR2_X1 U551 ( .A(n424), .B(KEYINPUT76), .ZN(n653) );
  OR2_X1 U552 ( .A1(n752), .A2(n426), .ZN(n425) );
  NAND2_X1 U553 ( .A1(n577), .A2(n669), .ZN(n587) );
  XNOR2_X2 U554 ( .A(n518), .B(n517), .ZN(n571) );
  NAND2_X1 U555 ( .A1(n659), .A2(n427), .ZN(n432) );
  NAND2_X1 U556 ( .A1(n444), .A2(n450), .ZN(n437) );
  NAND2_X1 U557 ( .A1(n448), .A2(n445), .ZN(n444) );
  NAND2_X1 U558 ( .A1(n443), .A2(KEYINPUT46), .ZN(n440) );
  INV_X1 U559 ( .A(n444), .ZN(n441) );
  NAND2_X1 U560 ( .A1(n443), .A2(n401), .ZN(n442) );
  INV_X1 U561 ( .A(n630), .ZN(n443) );
  NAND2_X1 U562 ( .A1(n630), .A2(n449), .ZN(n448) );
  INV_X1 U563 ( .A(KEYINPUT46), .ZN(n451) );
  NAND2_X1 U564 ( .A1(n584), .A2(KEYINPUT44), .ZN(n586) );
  BUF_X1 U565 ( .A(n732), .Z(n751) );
  INV_X1 U566 ( .A(n544), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n484), .B(G475), .ZN(n485) );
  XNOR2_X1 U568 ( .A(n486), .B(n485), .ZN(n595) );
  BUF_X1 U569 ( .A(n584), .Z(n604) );
  NAND2_X1 U570 ( .A1(n651), .A2(G234), .ZN(n457) );
  XNOR2_X1 U571 ( .A(n455), .B(KEYINPUT20), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n457), .B(n456), .ZN(n552) );
  OR2_X1 U573 ( .A1(n552), .A2(n458), .ZN(n459) );
  XNOR2_X1 U574 ( .A(n459), .B(KEYINPUT21), .ZN(n672) );
  XNOR2_X2 U575 ( .A(G143), .B(KEYINPUT64), .ZN(n461) );
  XNOR2_X2 U576 ( .A(n461), .B(n460), .ZN(n494) );
  BUF_X1 U577 ( .A(n494), .Z(n462) );
  XNOR2_X1 U578 ( .A(n463), .B(G122), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U580 ( .A(n467), .B(n466), .Z(n468) );
  XNOR2_X1 U581 ( .A(n462), .B(n468), .ZN(n470) );
  NAND2_X1 U582 ( .A1(n541), .A2(G217), .ZN(n469) );
  XNOR2_X1 U583 ( .A(n470), .B(n469), .ZN(n716) );
  NAND2_X1 U584 ( .A1(n716), .A2(n427), .ZN(n472) );
  XNOR2_X1 U585 ( .A(KEYINPUT105), .B(G478), .ZN(n471) );
  XNOR2_X1 U586 ( .A(n472), .B(n471), .ZN(n583) );
  XNOR2_X1 U587 ( .A(n474), .B(n473), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U589 ( .A(n478), .B(n477), .Z(n483) );
  NAND2_X1 U590 ( .A1(G214), .A2(n532), .ZN(n479) );
  XNOR2_X1 U591 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U592 ( .A(n481), .B(n784), .ZN(n482) );
  XNOR2_X1 U593 ( .A(n483), .B(n482), .ZN(n718) );
  NOR2_X1 U594 ( .A1(G902), .A2(n718), .ZN(n486) );
  XNOR2_X1 U595 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n484) );
  NAND2_X1 U596 ( .A1(n583), .A2(n595), .ZN(n690) );
  NOR2_X1 U597 ( .A1(n672), .A2(n690), .ZN(n487) );
  XNOR2_X1 U598 ( .A(n487), .B(KEYINPUT106), .ZN(n515) );
  XNOR2_X1 U599 ( .A(G101), .B(KEYINPUT66), .ZN(n488) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n500) );
  NAND2_X1 U601 ( .A1(n786), .A2(G224), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U604 ( .A1(n427), .A2(n502), .ZN(n505) );
  NAND2_X1 U605 ( .A1(n505), .A2(G210), .ZN(n503) );
  AND2_X1 U606 ( .A1(n505), .A2(G214), .ZN(n563) );
  XNOR2_X1 U607 ( .A(n506), .B(KEYINPUT14), .ZN(n509) );
  NAND2_X1 U608 ( .A1(n509), .A2(G902), .ZN(n507) );
  XNOR2_X1 U609 ( .A(KEYINPUT94), .B(n507), .ZN(n559) );
  INV_X1 U610 ( .A(n559), .ZN(n508) );
  NOR2_X1 U611 ( .A1(G898), .A2(n786), .ZN(n746) );
  NAND2_X1 U612 ( .A1(n508), .A2(n746), .ZN(n512) );
  NAND2_X1 U613 ( .A1(n509), .A2(G952), .ZN(n510) );
  XNOR2_X1 U614 ( .A(n510), .B(KEYINPUT92), .ZN(n704) );
  NOR2_X1 U615 ( .A1(n704), .A2(G953), .ZN(n511) );
  XNOR2_X1 U616 ( .A(n511), .B(KEYINPUT93), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n512), .A2(n562), .ZN(n513) );
  INV_X1 U618 ( .A(KEYINPUT0), .ZN(n514) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n516), .B(KEYINPUT22), .ZN(n517) );
  NAND2_X1 U621 ( .A1(n786), .A2(G227), .ZN(n522) );
  XNOR2_X1 U622 ( .A(n522), .B(KEYINPUT72), .ZN(n524) );
  XNOR2_X1 U623 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U624 ( .A(n526), .B(n525), .ZN(n527) );
  BUF_X1 U625 ( .A(n577), .Z(n670) );
  INV_X1 U626 ( .A(n670), .ZN(n556) );
  BUF_X1 U627 ( .A(n528), .Z(n529) );
  XNOR2_X1 U628 ( .A(n531), .B(n530), .ZN(n536) );
  NAND2_X1 U629 ( .A1(n532), .A2(G210), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U631 ( .A(n536), .B(n535), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U633 ( .A(n529), .B(n539), .ZN(n733) );
  NAND2_X1 U634 ( .A1(n733), .A2(n427), .ZN(n540) );
  XNOR2_X2 U635 ( .A(n540), .B(G472), .ZN(n620) );
  INV_X1 U636 ( .A(n620), .ZN(n676) );
  NAND2_X1 U637 ( .A1(n541), .A2(G221), .ZN(n542) );
  XNOR2_X1 U638 ( .A(n542), .B(n784), .ZN(n550) );
  XNOR2_X1 U639 ( .A(n544), .B(n543), .ZN(n548) );
  XNOR2_X1 U640 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U642 ( .A(G217), .ZN(n551) );
  XNOR2_X1 U643 ( .A(n553), .B(KEYINPUT25), .ZN(n554) );
  AND2_X1 U644 ( .A1(n676), .A2(n673), .ZN(n555) );
  AND2_X1 U645 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U646 ( .A1(n571), .A2(n557), .ZN(n602) );
  XOR2_X1 U647 ( .A(G110), .B(KEYINPUT115), .Z(n558) );
  XNOR2_X1 U648 ( .A(n602), .B(n558), .ZN(G12) );
  XNOR2_X1 U649 ( .A(n620), .B(KEYINPUT6), .ZN(n570) );
  INV_X1 U650 ( .A(n583), .ZN(n594) );
  OR2_X1 U651 ( .A1(n595), .A2(n594), .ZN(n773) );
  NOR2_X1 U652 ( .A1(n559), .A2(G900), .ZN(n560) );
  NAND2_X1 U653 ( .A1(G953), .A2(n560), .ZN(n561) );
  NAND2_X1 U654 ( .A1(n562), .A2(n561), .ZN(n617) );
  INV_X1 U655 ( .A(n563), .ZN(n687) );
  NAND2_X1 U656 ( .A1(n617), .A2(n687), .ZN(n564) );
  NOR2_X1 U657 ( .A1(n564), .A2(n672), .ZN(n565) );
  NAND2_X1 U658 ( .A1(n673), .A2(n565), .ZN(n566) );
  NOR2_X1 U659 ( .A1(n773), .A2(n566), .ZN(n567) );
  NAND2_X1 U660 ( .A1(n578), .A2(n567), .ZN(n634) );
  OR2_X1 U661 ( .A1(n634), .A2(n670), .ZN(n568) );
  XNOR2_X1 U662 ( .A(n568), .B(KEYINPUT43), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n569), .A2(n402), .ZN(n649) );
  XNOR2_X1 U664 ( .A(n649), .B(G140), .ZN(G42) );
  NOR2_X1 U665 ( .A1(n601), .A2(n670), .ZN(n573) );
  XNOR2_X1 U666 ( .A(n573), .B(n572), .ZN(n575) );
  INV_X1 U667 ( .A(n673), .ZN(n574) );
  NAND2_X1 U668 ( .A1(n575), .A2(n574), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(G101), .ZN(G3) );
  XNOR2_X1 U670 ( .A(n587), .B(KEYINPUT107), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U672 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n581), .B(n580), .ZN(n685) );
  NOR2_X1 U674 ( .A1(n595), .A2(n583), .ZN(n632) );
  XOR2_X1 U675 ( .A(G122), .B(n604), .Z(G24) );
  BUF_X1 U676 ( .A(n587), .Z(n588) );
  INV_X1 U677 ( .A(n588), .ZN(n589) );
  AND2_X1 U678 ( .A1(n589), .A2(n620), .ZN(n680) );
  XOR2_X1 U679 ( .A(KEYINPUT31), .B(n590), .Z(n775) );
  INV_X1 U680 ( .A(n607), .ZN(n592) );
  NOR2_X1 U681 ( .A1(n592), .A2(n620), .ZN(n593) );
  NAND2_X1 U682 ( .A1(n775), .A2(n761), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n776) );
  NAND2_X1 U684 ( .A1(n773), .A2(n776), .ZN(n692) );
  NAND2_X1 U685 ( .A1(n596), .A2(n692), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U687 ( .A(n670), .B(KEYINPUT90), .ZN(n638) );
  INV_X1 U688 ( .A(KEYINPUT45), .ZN(n605) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT30), .ZN(n609) );
  AND2_X1 U690 ( .A1(n609), .A2(n617), .ZN(n610) );
  XNOR2_X1 U691 ( .A(n633), .B(KEYINPUT38), .ZN(n688) );
  XNOR2_X1 U692 ( .A(KEYINPUT80), .B(KEYINPUT39), .ZN(n611) );
  INV_X1 U693 ( .A(n773), .ZN(n612) );
  INV_X1 U694 ( .A(KEYINPUT110), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT40), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n688), .A2(n687), .ZN(n693) );
  XNOR2_X1 U697 ( .A(KEYINPUT41), .B(n615), .ZN(n706) );
  INV_X1 U698 ( .A(n672), .ZN(n616) );
  AND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  AND2_X1 U700 ( .A1(n673), .A2(n618), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U702 ( .A(KEYINPUT28), .ZN(n621) );
  XNOR2_X1 U703 ( .A(n622), .B(n621), .ZN(n640) );
  NAND2_X1 U704 ( .A1(n640), .A2(n624), .ZN(n625) );
  NOR2_X1 U705 ( .A1(n706), .A2(n625), .ZN(n628) );
  INV_X1 U706 ( .A(KEYINPUT111), .ZN(n626) );
  XNOR2_X1 U707 ( .A(n626), .B(KEYINPUT42), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n628), .B(n627), .ZN(n793) );
  INV_X1 U709 ( .A(n793), .ZN(n629) );
  INV_X1 U710 ( .A(n402), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n634), .A2(n402), .ZN(n636) );
  XNOR2_X1 U712 ( .A(KEYINPUT36), .B(KEYINPUT86), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n779) );
  AND2_X1 U715 ( .A1(n639), .A2(n624), .ZN(n641) );
  AND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n770) );
  NAND2_X1 U717 ( .A1(n770), .A2(n692), .ZN(n643) );
  INV_X1 U718 ( .A(KEYINPUT70), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n644), .A2(KEYINPUT47), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n644), .A2(KEYINPUT47), .ZN(n645) );
  AND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  AND2_X1 U723 ( .A1(n779), .A2(n647), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n423), .A2(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n658) );
  INV_X1 U726 ( .A(n739), .ZN(n657) );
  INV_X1 U727 ( .A(KEYINPUT2), .ZN(n662) );
  NOR2_X1 U728 ( .A1(n655), .A2(n662), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n667) );
  AND2_X2 U730 ( .A1(n658), .A2(n667), .ZN(n732) );
  AND2_X2 U731 ( .A1(n751), .A2(G217), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  INV_X1 U733 ( .A(n736), .ZN(n757) );
  NOR2_X1 U734 ( .A1(n661), .A2(n757), .ZN(G66) );
  NAND2_X1 U735 ( .A1(n662), .A2(KEYINPUT75), .ZN(n663) );
  NOR2_X1 U736 ( .A1(n785), .A2(n663), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n739), .A2(n664), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n711) );
  NOR2_X1 U740 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(KEYINPUT50), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n675) );
  XOR2_X1 U743 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n681) );
  OR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(n682), .Z(n684) );
  INV_X1 U749 ( .A(n706), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n700) );
  BUF_X1 U751 ( .A(n685), .Z(n686) );
  INV_X1 U752 ( .A(n686), .ZN(n705) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U755 ( .A(KEYINPUT119), .B(n691), .Z(n696) );
  INV_X1 U756 ( .A(n692), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n705), .A2(n697), .ZN(n698) );
  XOR2_X1 U760 ( .A(KEYINPUT120), .B(n698), .Z(n699) );
  NAND2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U762 ( .A(n701), .B(KEYINPUT121), .ZN(n702) );
  XNOR2_X1 U763 ( .A(n702), .B(KEYINPUT52), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n709), .B(KEYINPUT122), .ZN(n710) );
  NAND2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U769 ( .A(n712), .B(KEYINPUT123), .ZN(n713) );
  NAND2_X1 U770 ( .A1(n713), .A2(n786), .ZN(n714) );
  XOR2_X1 U771 ( .A(KEYINPUT53), .B(n714), .Z(G75) );
  NAND2_X1 U772 ( .A1(n732), .A2(G478), .ZN(n715) );
  XOR2_X1 U773 ( .A(n716), .B(n715), .Z(n717) );
  NOR2_X1 U774 ( .A1(n717), .A2(n757), .ZN(G63) );
  XOR2_X1 U775 ( .A(n443), .B(G131), .Z(G33) );
  NAND2_X1 U776 ( .A1(n732), .A2(G475), .ZN(n720) );
  XNOR2_X1 U777 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U778 ( .A1(n721), .A2(n736), .ZN(n723) );
  INV_X1 U779 ( .A(KEYINPUT60), .ZN(n722) );
  XNOR2_X1 U780 ( .A(n723), .B(n722), .ZN(G60) );
  NAND2_X1 U781 ( .A1(n732), .A2(G210), .ZN(n728) );
  XNOR2_X1 U782 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n724) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT55), .ZN(n725) );
  XNOR2_X1 U784 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U785 ( .A1(n729), .A2(n736), .ZN(n731) );
  INV_X1 U786 ( .A(KEYINPUT56), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n731), .B(n730), .ZN(G51) );
  NAND2_X1 U788 ( .A1(n732), .A2(G472), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U791 ( .A(n738), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U792 ( .A1(n739), .A2(G953), .ZN(n745) );
  XOR2_X1 U793 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n741) );
  NAND2_X1 U794 ( .A1(G224), .A2(G953), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U796 ( .A1(G898), .A2(n742), .ZN(n743) );
  XOR2_X1 U797 ( .A(KEYINPUT126), .B(n743), .Z(n744) );
  NOR2_X1 U798 ( .A1(n745), .A2(n744), .ZN(n750) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n748), .B(KEYINPUT127), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(G69) );
  NAND2_X1 U802 ( .A1(n751), .A2(G469), .ZN(n756) );
  XOR2_X1 U803 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n753) );
  XNOR2_X1 U804 ( .A(n753), .B(KEYINPUT58), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n752), .B(n754), .ZN(n755) );
  XNOR2_X1 U806 ( .A(n756), .B(n755), .ZN(n758) );
  NOR2_X1 U807 ( .A1(n758), .A2(n757), .ZN(G54) );
  NOR2_X1 U808 ( .A1(n761), .A2(n773), .ZN(n759) );
  XOR2_X1 U809 ( .A(KEYINPUT112), .B(n759), .Z(n760) );
  XNOR2_X1 U810 ( .A(G104), .B(n760), .ZN(G6) );
  NOR2_X1 U811 ( .A1(n761), .A2(n776), .ZN(n766) );
  XOR2_X1 U812 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n763) );
  XNOR2_X1 U813 ( .A(G107), .B(KEYINPUT113), .ZN(n762) );
  XNOR2_X1 U814 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U815 ( .A(KEYINPUT26), .B(n764), .ZN(n765) );
  XNOR2_X1 U816 ( .A(n766), .B(n765), .ZN(G9) );
  XOR2_X1 U817 ( .A(G128), .B(KEYINPUT29), .Z(n768) );
  NAND2_X1 U818 ( .A1(n770), .A2(n352), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(G30) );
  XNOR2_X1 U820 ( .A(G143), .B(n769), .ZN(G45) );
  NAND2_X1 U821 ( .A1(n770), .A2(n612), .ZN(n771) );
  XNOR2_X1 U822 ( .A(n771), .B(KEYINPUT116), .ZN(n772) );
  XNOR2_X1 U823 ( .A(G146), .B(n772), .ZN(G48) );
  NOR2_X1 U824 ( .A1(n773), .A2(n775), .ZN(n774) );
  XOR2_X1 U825 ( .A(G113), .B(n774), .Z(G15) );
  NOR2_X1 U826 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U827 ( .A(G116), .B(n777), .Z(G18) );
  XOR2_X1 U828 ( .A(G125), .B(KEYINPUT37), .Z(n778) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(G27) );
  XOR2_X1 U830 ( .A(G134), .B(n780), .Z(n781) );
  XNOR2_X1 U831 ( .A(n781), .B(KEYINPUT117), .ZN(G36) );
  BUF_X1 U832 ( .A(n782), .Z(n783) );
  XNOR2_X1 U833 ( .A(n783), .B(n784), .ZN(n788) );
  XNOR2_X1 U834 ( .A(n785), .B(n788), .ZN(n787) );
  NAND2_X1 U835 ( .A1(n787), .A2(n786), .ZN(n792) );
  XNOR2_X1 U836 ( .A(n788), .B(G227), .ZN(n789) );
  NAND2_X1 U837 ( .A1(n789), .A2(G900), .ZN(n790) );
  NAND2_X1 U838 ( .A1(n790), .A2(G953), .ZN(n791) );
  NAND2_X1 U839 ( .A1(n792), .A2(n791), .ZN(G72) );
  XOR2_X1 U840 ( .A(G137), .B(n447), .Z(G39) );
  XNOR2_X1 U841 ( .A(n794), .B(G119), .ZN(G21) );
endmodule

