//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G567), .B1(G2106), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n465), .A2(new_n472), .A3(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n471), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(new_n468), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(G138), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n461), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT3), .B1(new_n469), .B2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(KEYINPUT71), .B(new_n487), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n468), .B2(new_n470), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n488), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n498));
  OAI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n479), .A2(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n495), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XOR2_X1   g083(.A(KEYINPUT5), .B(G543), .Z(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT72), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .A3(G651), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n515), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n515), .B2(new_n517), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n512), .A2(KEYINPUT73), .A3(new_n521), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n520), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(new_n519), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n536), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n532), .A2(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n520), .A2(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n523), .A2(G52), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n514), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n523), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n520), .A2(G81), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n520), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n532), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n523), .A2(new_n562), .A3(G53), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n565));
  OAI221_X1 g140(.A(new_n560), .B1(new_n514), .B2(new_n561), .C1(new_n564), .C2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  AND2_X1   g143(.A1(new_n527), .A2(new_n528), .ZN(G303));
  NAND2_X1  g144(.A1(new_n520), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n523), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(G86), .A2(new_n520), .B1(new_n523), .B2(G48), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n518), .B2(new_n519), .ZN(new_n576));
  AND2_X1   g151(.A1(G73), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n514), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  AOI22_X1  g160(.A1(G85), .A2(new_n520), .B1(new_n523), .B2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  INV_X1    g170(.A(new_n520), .ZN(new_n596));
  OR3_X1    g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n509), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n591), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n591), .B1(new_n603), .B2(G868), .ZN(G321));
  NOR2_X1   g180(.A1(G299), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G868), .B2(G168), .ZN(G280));
  XOR2_X1   g182(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g183(.A(new_n603), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G559), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G860), .B2(new_n603), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT81), .ZN(G148));
  OAI21_X1  g187(.A(KEYINPUT82), .B1(new_n554), .B2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n613), .B(KEYINPUT82), .S(new_n615), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n474), .A2(new_n461), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(G2100), .ZN(new_n622));
  AOI22_X1  g197(.A1(G135), .A2(new_n471), .B1(new_n479), .B2(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n625), .B2(new_n624), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n621), .A2(new_n622), .A3(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n630), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(new_n675), .B(new_n674), .S(new_n667), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G1981), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G1986), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G1986), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  AND3_X1   g261(.A1(new_n680), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n686), .B1(new_n680), .B2(new_n684), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n665), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n680), .A2(new_n684), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(new_n685), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n680), .A2(new_n684), .A3(new_n686), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n664), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(new_n693), .ZN(G229));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT33), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1976), .ZN(new_n701));
  NOR2_X1   g276(.A1(G6), .A2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G305), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n696), .A2(G24), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n589), .B2(new_n696), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n471), .A2(G131), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n479), .A2(G119), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  NOR3_X1   g304(.A1(new_n715), .A2(new_n718), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n695), .B1(new_n714), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n714), .A2(new_n695), .A3(new_n730), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n732), .A2(KEYINPUT36), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT36), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(G162), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G29), .B2(G35), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT29), .B(G2090), .Z(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n740), .B2(KEYINPUT24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(KEYINPUT24), .B2(new_n740), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n465), .A2(new_n472), .A3(new_n475), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n719), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2072), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n719), .A2(G33), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT25), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n471), .A2(G139), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n749), .B(new_n750), .C1(new_n478), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT92), .B(G2067), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n719), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n471), .A2(G140), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT91), .B1(G104), .B2(G2105), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(KEYINPUT91), .A2(G104), .A3(G2105), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(G116), .B2(new_n478), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n479), .A2(G128), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n757), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(new_n719), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n745), .B1(new_n746), .B2(new_n753), .C1(new_n754), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n554), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G16), .B2(G19), .ZN(new_n768));
  INV_X1    g343(.A(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n737), .B2(new_n738), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n768), .A2(new_n769), .B1(new_n739), .B2(new_n744), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n766), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n474), .A2(G105), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n471), .A2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n479), .A2(G129), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND4_X1  g353(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G32), .B(new_n779), .S(G29), .Z(new_n780));
  XOR2_X1   g355(.A(KEYINPUT27), .B(G1996), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n609), .A2(G16), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n696), .A2(G4), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n782), .B1(new_n786), .B2(G1348), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G21), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G168), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1966), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n765), .A2(new_n754), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT30), .B(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  NAND2_X1  g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n793), .A2(new_n719), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n796), .C1(new_n719), .C2(new_n629), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n785), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n773), .A2(new_n787), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n696), .A2(G5), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G171), .B2(new_n696), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n802), .A2(G1961), .B1(new_n753), .B2(new_n746), .ZN(new_n803));
  NOR2_X1   g378(.A1(G27), .A2(G29), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G164), .B2(G29), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n803), .B1(G1961), .B2(new_n802), .C1(G2078), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n805), .A2(G2078), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n696), .A2(G20), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT23), .Z(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G299), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1956), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n800), .A2(new_n806), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT93), .Z(new_n814));
  NOR3_X1   g389(.A1(new_n734), .A2(new_n735), .A3(new_n814), .ZN(G311));
  OR3_X1    g390(.A1(new_n734), .A2(new_n735), .A3(new_n814), .ZN(G150));
  XNOR2_X1  g391(.A(KEYINPUT97), .B(G860), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n603), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(G80), .A2(G543), .ZN(new_n821));
  INV_X1    g396(.A(G67), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n509), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G651), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT94), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT95), .B(G93), .Z(new_n826));
  AOI22_X1  g401(.A1(new_n520), .A2(new_n826), .B1(new_n523), .B2(G55), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n824), .B2(KEYINPUT94), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT96), .ZN(new_n830));
  OR3_X1    g405(.A1(new_n825), .A2(new_n828), .A3(KEYINPUT96), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n553), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n554), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n820), .B(new_n834), .Z(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n818), .B1(new_n836), .B2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(KEYINPUT39), .B2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n830), .A2(new_n831), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n818), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(G145));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT100), .B(G37), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n506), .B(new_n764), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n779), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n752), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n725), .B(KEYINPUT99), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n619), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n479), .A2(G130), .ZN(new_n851));
  OR2_X1    g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(G2104), .C1(G118), .C2(new_n478), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G142), .B2(new_n471), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n850), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n848), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n743), .B(KEYINPUT98), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n629), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n845), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n860), .B(KEYINPUT102), .Z(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  OR3_X1    g438(.A1(new_n848), .A2(new_n863), .A3(new_n856), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n848), .A2(new_n863), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n848), .A2(new_n856), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n862), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n843), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n861), .A2(new_n867), .A3(new_n843), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(G395));
  INV_X1    g449(.A(KEYINPUT110), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n839), .B2(new_n614), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n603), .B(G299), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT106), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n603), .B2(G299), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n877), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n834), .B(new_n610), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n890));
  NAND2_X1  g465(.A1(G303), .A2(G305), .ZN(new_n891));
  NAND2_X1  g466(.A1(G166), .A2(new_n703), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n589), .B(new_n698), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT108), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT107), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n887), .A2(new_n888), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n890), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G868), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n890), .B2(new_n902), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n876), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n907), .A2(new_n875), .A3(G868), .A4(new_n903), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(G295));
  AND2_X1   g484(.A1(new_n906), .A2(new_n908), .ZN(G331));
  NAND3_X1  g485(.A1(new_n832), .A2(G168), .A3(new_n833), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G168), .B1(new_n832), .B2(new_n833), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n912), .A2(G301), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(G301), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n884), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n879), .B(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n915), .B(new_n916), .C1(new_n917), .C2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n883), .ZN(new_n921));
  INV_X1    g496(.A(new_n916), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n899), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n920), .A2(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n899), .A2(KEYINPUT111), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n896), .A2(new_n929), .A3(new_n898), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT43), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n916), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n883), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n877), .A4(new_n916), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n934), .A2(new_n928), .A3(new_n930), .A4(new_n935), .ZN(new_n936));
  AND4_X1   g511(.A1(KEYINPUT43), .A2(new_n936), .A3(new_n844), .A4(new_n924), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n926), .B2(new_n931), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n940), .A2(new_n936), .A3(new_n844), .A4(new_n924), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n943), .ZN(G397));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n779), .B(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n763), .B(G2067), .Z(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n725), .B(new_n728), .Z(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  INV_X1    g526(.A(new_n488), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n485), .B1(new_n493), .B2(KEYINPUT71), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT71), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n952), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n951), .B1(new_n957), .B2(new_n504), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(G160), .A2(G40), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n683), .A3(new_n589), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n950), .A2(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n965), .B2(new_n964), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT46), .B1(new_n962), .B2(new_n945), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT127), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n779), .B1(KEYINPUT46), .B2(new_n945), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n947), .A2(new_n972), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n970), .A2(new_n971), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT47), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n726), .A2(new_n728), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n948), .A2(new_n976), .B1(G2067), .B2(new_n763), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n967), .B(new_n975), .C1(new_n962), .C2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n527), .A2(new_n528), .A3(G8), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT55), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n958), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n506), .A2(KEYINPUT112), .A3(new_n951), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n961), .B1(KEYINPUT50), .B2(new_n958), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n743), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n958), .B2(new_n959), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n495), .B2(new_n505), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n989), .A2(G2090), .B1(new_n995), .B2(G1971), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n980), .A2(new_n981), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n982), .A2(G8), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT115), .B(G1981), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n574), .B(new_n999), .C1(new_n580), .C2(new_n581), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n523), .A2(G48), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT116), .B(G86), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n578), .B(new_n1001), .C1(new_n596), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G1981), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n984), .A2(new_n985), .A3(new_n991), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(KEYINPUT49), .A3(new_n1004), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1006), .A2(G8), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G288), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1012), .A3(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1007), .A2(new_n1012), .A3(G8), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G288), .A2(G1976), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1009), .A2(new_n1018), .B1(new_n703), .B2(new_n999), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1007), .A2(G8), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT117), .Z(new_n1021));
  OAI22_X1  g596(.A1(new_n998), .A2(new_n1017), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1017), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n998), .A2(new_n1023), .A3(KEYINPUT63), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n984), .A2(new_n985), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n992), .B1(new_n1026), .B2(new_n959), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT118), .B1(new_n1027), .B2(G1966), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n984), .B2(new_n985), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1029), .B(new_n790), .C1(new_n1030), .C2(new_n992), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n989), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT119), .B(G2084), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1025), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n996), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n996), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n980), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1024), .A2(G168), .A3(new_n1036), .A4(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(G168), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n986), .B1(new_n984), .B2(new_n985), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n991), .B1(new_n958), .B2(KEYINPUT50), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n961), .B1(KEYINPUT45), .B2(new_n993), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n960), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1047), .A2(new_n1048), .B1(new_n709), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n980), .B1(new_n1051), .B2(new_n1025), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n998), .A2(new_n1052), .A3(new_n1023), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1043), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1022), .B1(new_n1042), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n993), .A2(KEYINPUT112), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n983), .B(G1384), .C1(new_n495), .C2(new_n505), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n959), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1049), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1029), .B1(new_n1059), .B2(new_n790), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1031), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1035), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OR3_X1    g638(.A1(G168), .A2(KEYINPUT123), .A3(new_n1025), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT123), .B1(G168), .B2(new_n1025), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1036), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1066), .B(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1036), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(KEYINPUT125), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(KEYINPUT51), .C1(new_n1036), .C2(new_n1073), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1068), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(G299), .B(KEYINPUT57), .Z(new_n1079));
  OAI21_X1  g654(.A(new_n811), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n995), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n987), .B2(new_n988), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1007), .A2(G2067), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n609), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1080), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1084), .A2(new_n1086), .A3(new_n603), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1089), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1083), .ZN(new_n1095));
  OR4_X1    g670(.A1(KEYINPUT60), .A2(new_n1084), .A3(new_n1086), .A4(new_n609), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1079), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1089), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1050), .B2(G1996), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n995), .A2(KEYINPUT122), .A3(new_n945), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1007), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n554), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1107), .B2(new_n554), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1090), .B1(new_n1101), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1050), .B2(G2078), .ZN(new_n1114));
  INV_X1    g689(.A(G1961), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n989), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G2078), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n995), .A2(KEYINPUT53), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1058), .A2(KEYINPUT53), .A3(new_n1117), .A4(new_n1049), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1114), .A2(new_n1121), .A3(new_n1116), .A4(G301), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1120), .A2(KEYINPUT54), .A3(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT126), .B(KEYINPUT54), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1114), .A2(new_n1121), .A3(new_n1116), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G171), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1114), .A2(new_n1116), .A3(G301), .A4(new_n1118), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1123), .A2(new_n1128), .A3(new_n1053), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1112), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1055), .B1(new_n1078), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1078), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1053), .A2(new_n1126), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1073), .B1(new_n1062), .B2(G8), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT125), .B1(new_n1135), .B2(new_n1069), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1071), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1077), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1068), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1134), .B1(new_n1140), .B2(KEYINPUT62), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1131), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n589), .B(G1986), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n963), .B1(new_n950), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n978), .B1(new_n1142), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g720(.A(G319), .ZN(new_n1147));
  NOR3_X1   g721(.A1(G401), .A2(new_n1147), .A3(G227), .ZN(new_n1148));
  AND3_X1   g722(.A1(new_n689), .A2(new_n693), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g723(.A(new_n870), .ZN(new_n1150));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1150), .B2(new_n868), .ZN(new_n1151));
  NOR2_X1   g725(.A1(new_n941), .A2(new_n942), .ZN(new_n1152));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n1152), .ZN(G308));
  OAI221_X1 g727(.A(new_n1149), .B1(new_n1150), .B2(new_n868), .C1(new_n941), .C2(new_n942), .ZN(G225));
endmodule


