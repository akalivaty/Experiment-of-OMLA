

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761;

  BUF_X1 U372 ( .A(n672), .Z(n623) );
  NOR2_X1 U373 ( .A1(G237), .A2(G953), .ZN(n438) );
  NOR2_X1 U374 ( .A1(n753), .A2(n583), .ZN(n624) );
  OR2_X1 U375 ( .A1(n685), .A2(n675), .ZN(n510) );
  INV_X1 U376 ( .A(G953), .ZN(n745) );
  NAND2_X1 U377 ( .A1(n413), .A2(n649), .ZN(n613) );
  NOR2_X2 U378 ( .A1(n607), .A2(n601), .ZN(n619) );
  XNOR2_X2 U379 ( .A(n379), .B(G131), .ZN(n479) );
  XNOR2_X2 U380 ( .A(G146), .B(KEYINPUT69), .ZN(n379) );
  XNOR2_X2 U381 ( .A(n443), .B(G101), .ZN(n495) );
  XNOR2_X2 U382 ( .A(KEYINPUT3), .B(G119), .ZN(n443) );
  XNOR2_X2 U383 ( .A(n613), .B(KEYINPUT31), .ZN(n731) );
  AND2_X1 U384 ( .A1(n620), .A2(n373), .ZN(n372) );
  XNOR2_X1 U385 ( .A(n371), .B(n370), .ZN(n369) );
  NOR2_X1 U386 ( .A1(n557), .A2(n435), .ZN(n388) );
  NOR2_X1 U387 ( .A1(n733), .A2(n722), .ZN(n387) );
  AND2_X1 U388 ( .A1(n567), .A2(n590), .ZN(n733) );
  XNOR2_X1 U389 ( .A(n594), .B(n593), .ZN(n376) );
  XNOR2_X1 U390 ( .A(n366), .B(n365), .ZN(n435) );
  XNOR2_X1 U391 ( .A(n600), .B(n599), .ZN(n669) );
  AND2_X1 U392 ( .A1(n398), .A2(n396), .ZN(n395) );
  XNOR2_X1 U393 ( .A(n385), .B(KEYINPUT1), .ZN(n610) );
  OR2_X1 U394 ( .A1(n708), .A2(G902), .ZN(n523) );
  XNOR2_X1 U395 ( .A(n368), .B(KEYINPUT65), .ZN(n349) );
  XNOR2_X1 U396 ( .A(n368), .B(KEYINPUT65), .ZN(n350) );
  XNOR2_X1 U397 ( .A(n368), .B(KEYINPUT65), .ZN(n705) );
  NAND2_X2 U398 ( .A1(n419), .A2(n416), .ZN(n368) );
  XOR2_X1 U399 ( .A(n459), .B(G140), .Z(n478) );
  XNOR2_X1 U400 ( .A(G125), .B(KEYINPUT10), .ZN(n459) );
  NAND2_X1 U401 ( .A1(n618), .A2(n667), .ZN(n371) );
  AND2_X1 U402 ( .A1(n431), .A2(n430), .ZN(n429) );
  AND2_X1 U403 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U404 ( .A(G237), .ZN(n448) );
  XNOR2_X1 U405 ( .A(n456), .B(n412), .ZN(n471) );
  INV_X1 U406 ( .A(KEYINPUT8), .ZN(n412) );
  XOR2_X1 U407 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n485) );
  XNOR2_X1 U408 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U409 ( .A(KEYINPUT85), .ZN(n403) );
  NOR2_X1 U410 ( .A1(n672), .A2(KEYINPUT2), .ZN(n407) );
  XNOR2_X1 U411 ( .A(n382), .B(n356), .ZN(n414) );
  NAND2_X1 U412 ( .A1(n383), .A2(n616), .ZN(n382) );
  INV_X1 U413 ( .A(KEYINPUT19), .ZN(n397) );
  OR2_X1 U414 ( .A1(n628), .A2(n397), .ZN(n396) );
  XNOR2_X1 U415 ( .A(n495), .B(n494), .ZN(n360) );
  XNOR2_X1 U416 ( .A(G119), .B(G137), .ZN(n453) );
  XNOR2_X1 U417 ( .A(G128), .B(G110), .ZN(n454) );
  XNOR2_X1 U418 ( .A(n457), .B(n410), .ZN(n409) );
  XNOR2_X1 U419 ( .A(G146), .B(KEYINPUT24), .ZN(n457) );
  XNOR2_X1 U420 ( .A(KEYINPUT95), .B(KEYINPUT83), .ZN(n410) );
  INV_X1 U421 ( .A(KEYINPUT70), .ZN(n460) );
  XNOR2_X1 U422 ( .A(G116), .B(G107), .ZN(n496) );
  OR2_X1 U423 ( .A1(n676), .A2(KEYINPUT66), .ZN(n421) );
  INV_X1 U424 ( .A(KEYINPUT66), .ZN(n417) );
  NOR2_X1 U425 ( .A1(n596), .A2(n541), .ZN(n543) );
  BUF_X1 U426 ( .A(n610), .Z(n639) );
  AND2_X1 U427 ( .A1(n615), .A2(n434), .ZN(n432) );
  INV_X1 U428 ( .A(KEYINPUT104), .ZN(n434) );
  INV_X1 U429 ( .A(KEYINPUT47), .ZN(n365) );
  INV_X1 U430 ( .A(KEYINPUT106), .ZN(n370) );
  XNOR2_X1 U431 ( .A(G116), .B(G113), .ZN(n439) );
  XOR2_X1 U432 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n440) );
  XNOR2_X1 U433 ( .A(n574), .B(KEYINPUT88), .ZN(n575) );
  NAND2_X1 U434 ( .A1(G237), .A2(G234), .ZN(n524) );
  XNOR2_X1 U435 ( .A(n490), .B(n489), .ZN(n692) );
  XNOR2_X1 U436 ( .A(n479), .B(n437), .ZN(n378) );
  XNOR2_X1 U437 ( .A(KEYINPUT4), .B(G137), .ZN(n437) );
  XNOR2_X1 U438 ( .A(G104), .B(G140), .ZN(n511) );
  XOR2_X1 U439 ( .A(KEYINPUT76), .B(KEYINPUT70), .Z(n512) );
  XNOR2_X1 U440 ( .A(KEYINPUT73), .B(G110), .ZN(n517) );
  XNOR2_X1 U441 ( .A(G107), .B(G101), .ZN(n516) );
  XNOR2_X1 U442 ( .A(n401), .B(n622), .ZN(n625) );
  NAND2_X1 U443 ( .A1(n405), .A2(n402), .ZN(n401) );
  AND2_X1 U444 ( .A1(n552), .A2(n551), .ZN(n554) );
  NOR2_X1 U445 ( .A1(n550), .A2(n640), .ZN(n551) );
  AND2_X1 U446 ( .A1(n564), .A2(n628), .ZN(n576) );
  INV_X1 U447 ( .A(KEYINPUT79), .ZN(n362) );
  OR2_X1 U448 ( .A1(n385), .A2(n538), .ZN(n547) );
  NAND2_X1 U449 ( .A1(n395), .A2(n392), .ZN(n587) );
  NAND2_X1 U450 ( .A1(n394), .A2(n393), .ZN(n392) );
  AND2_X1 U451 ( .A1(n628), .A2(n397), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n458), .B(n408), .ZN(n461) );
  XNOR2_X1 U453 ( .A(n411), .B(n409), .ZN(n408) );
  XNOR2_X1 U454 ( .A(n470), .B(n476), .ZN(n700) );
  NAND2_X1 U455 ( .A1(n418), .A2(n417), .ZN(n416) );
  XOR2_X1 U456 ( .A(n692), .B(KEYINPUT59), .Z(n693) );
  XNOR2_X1 U457 ( .A(n686), .B(n687), .ZN(n688) );
  BUF_X1 U458 ( .A(n745), .Z(n367) );
  XNOR2_X1 U459 ( .A(n545), .B(KEYINPUT42), .ZN(n761) );
  NAND2_X1 U460 ( .A1(n436), .A2(n544), .ZN(n545) );
  INV_X1 U461 ( .A(KEYINPUT35), .ZN(n377) );
  AND2_X1 U462 ( .A1(n639), .A2(n598), .ZN(n400) );
  NOR2_X1 U463 ( .A1(n573), .A2(n572), .ZN(n727) );
  AND2_X1 U464 ( .A1(n617), .A2(n639), .ZN(n375) );
  AND2_X1 U465 ( .A1(n413), .A2(n355), .ZN(n351) );
  XNOR2_X1 U466 ( .A(n467), .B(n466), .ZN(n537) );
  OR2_X2 U467 ( .A1(n537), .A2(n642), .ZN(n640) );
  AND2_X1 U468 ( .A1(G217), .A2(n468), .ZN(n352) );
  XOR2_X1 U469 ( .A(n363), .B(n362), .Z(n353) );
  NOR2_X1 U470 ( .A1(n631), .A2(n642), .ZN(n354) );
  AND2_X1 U471 ( .A1(n549), .A2(n614), .ZN(n355) );
  XNOR2_X1 U472 ( .A(KEYINPUT92), .B(KEYINPUT33), .ZN(n356) );
  XOR2_X1 U473 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n357) );
  XNOR2_X1 U474 ( .A(n360), .B(n497), .ZN(n744) );
  XNOR2_X1 U475 ( .A(n358), .B(n691), .ZN(G51) );
  NAND2_X1 U476 ( .A1(n690), .A2(n702), .ZN(n358) );
  XNOR2_X1 U477 ( .A(n359), .B(n696), .ZN(G60) );
  NAND2_X1 U478 ( .A1(n695), .A2(n702), .ZN(n359) );
  NAND2_X1 U479 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U480 ( .A(n386), .B(n575), .ZN(n364) );
  AND2_X1 U481 ( .A1(n422), .A2(n420), .ZN(n419) );
  NOR2_X1 U482 ( .A1(n610), .A2(n640), .ZN(n383) );
  XNOR2_X2 U483 ( .A(n361), .B(n588), .ZN(n595) );
  NAND2_X1 U484 ( .A1(n354), .A2(n413), .ZN(n361) );
  NAND2_X1 U485 ( .A1(n590), .A2(n589), .ZN(n363) );
  NAND2_X1 U486 ( .A1(n376), .A2(n669), .ZN(n391) );
  NAND2_X1 U487 ( .A1(n364), .A2(n582), .ZN(n671) );
  NOR2_X1 U488 ( .A1(n724), .A2(n633), .ZN(n366) );
  NAND2_X1 U489 ( .A1(n471), .A2(G221), .ZN(n411) );
  NAND2_X1 U490 ( .A1(n372), .A2(n369), .ZN(n621) );
  NAND2_X1 U491 ( .A1(n374), .A2(n389), .ZN(n373) );
  NAND2_X1 U492 ( .A1(n390), .A2(n608), .ZN(n374) );
  XNOR2_X2 U493 ( .A(n399), .B(n357), .ZN(n413) );
  NAND2_X1 U494 ( .A1(n595), .A2(n375), .ZN(n667) );
  XNOR2_X1 U495 ( .A(n376), .B(G119), .ZN(G21) );
  XNOR2_X1 U496 ( .A(n607), .B(G122), .ZN(G24) );
  XNOR2_X2 U497 ( .A(n606), .B(n377), .ZN(n607) );
  XNOR2_X2 U498 ( .A(n470), .B(n378), .ZN(n751) );
  XNOR2_X2 U499 ( .A(n501), .B(G134), .ZN(n470) );
  XNOR2_X2 U500 ( .A(n381), .B(n380), .ZN(n501) );
  XNOR2_X2 U501 ( .A(KEYINPUT64), .B(KEYINPUT81), .ZN(n380) );
  XNOR2_X2 U502 ( .A(G143), .B(G128), .ZN(n381) );
  INV_X1 U503 ( .A(n414), .ZN(n415) );
  XNOR2_X2 U504 ( .A(n597), .B(n560), .ZN(n616) );
  NAND2_X1 U505 ( .A1(n384), .A2(n761), .ZN(n556) );
  XNOR2_X1 U506 ( .A(n384), .B(G131), .ZN(G33) );
  XNOR2_X2 U507 ( .A(n555), .B(KEYINPUT40), .ZN(n384) );
  XNOR2_X2 U508 ( .A(n523), .B(n522), .ZN(n385) );
  NOR2_X1 U509 ( .A1(n597), .A2(n385), .ZN(n614) );
  NOR2_X1 U510 ( .A1(n568), .A2(n385), .ZN(n436) );
  INV_X1 U511 ( .A(n391), .ZN(n390) );
  NAND2_X1 U512 ( .A1(n391), .A2(n601), .ZN(n389) );
  INV_X1 U513 ( .A(n570), .ZN(n394) );
  NAND2_X1 U514 ( .A1(n570), .A2(KEYINPUT19), .ZN(n398) );
  NAND2_X1 U515 ( .A1(n587), .A2(n586), .ZN(n399) );
  NAND2_X1 U516 ( .A1(n595), .A2(n400), .ZN(n600) );
  NAND2_X1 U517 ( .A1(n753), .A2(n583), .ZN(n404) );
  XNOR2_X1 U518 ( .A(n407), .B(n406), .ZN(n405) );
  INV_X1 U519 ( .A(KEYINPUT84), .ZN(n406) );
  NAND2_X1 U520 ( .A1(n414), .A2(n413), .ZN(n603) );
  NOR2_X1 U521 ( .A1(n415), .A2(n658), .ZN(n659) );
  NOR2_X1 U522 ( .A1(n638), .A2(n415), .ZN(n653) );
  NAND2_X1 U523 ( .A1(n424), .A2(n423), .ZN(n422) );
  XNOR2_X2 U524 ( .A(n674), .B(KEYINPUT86), .ZN(n424) );
  INV_X1 U525 ( .A(n424), .ZN(n418) );
  AND2_X1 U526 ( .A1(n677), .A2(n421), .ZN(n420) );
  AND2_X1 U527 ( .A1(n676), .A2(KEYINPUT66), .ZN(n423) );
  NAND2_X1 U528 ( .A1(n425), .A2(n429), .ZN(n618) );
  NAND2_X1 U529 ( .A1(n731), .A2(n432), .ZN(n426) );
  NAND2_X1 U530 ( .A1(n433), .A2(n428), .ZN(n427) );
  INV_X1 U531 ( .A(n731), .ZN(n428) );
  OR2_X1 U532 ( .A1(n615), .A2(n434), .ZN(n430) );
  NAND2_X1 U533 ( .A1(n351), .A2(n432), .ZN(n431) );
  NOR2_X1 U534 ( .A1(n351), .A2(n434), .ZN(n433) );
  XNOR2_X2 U535 ( .A(n483), .B(G104), .ZN(n494) );
  INV_X1 U536 ( .A(KEYINPUT48), .ZN(n574) );
  INV_X1 U537 ( .A(KEYINPUT82), .ZN(n622) );
  XNOR2_X1 U538 ( .A(n451), .B(KEYINPUT23), .ZN(n452) );
  XNOR2_X1 U539 ( .A(n453), .B(n452), .ZN(n455) );
  INV_X1 U540 ( .A(KEYINPUT87), .ZN(n626) );
  INV_X1 U541 ( .A(KEYINPUT53), .ZN(n665) );
  XOR2_X1 U542 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n450) );
  XNOR2_X1 U543 ( .A(n438), .B(KEYINPUT74), .ZN(n480) );
  NAND2_X1 U544 ( .A1(n480), .A2(G210), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U546 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U547 ( .A(n444), .B(n495), .ZN(n445) );
  XNOR2_X1 U548 ( .A(n751), .B(n445), .ZN(n678) );
  OR2_X2 U549 ( .A1(n678), .A2(G902), .ZN(n447) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(G472), .ZN(n446) );
  XNOR2_X2 U551 ( .A(n447), .B(n446), .ZN(n597) );
  INV_X1 U552 ( .A(G902), .ZN(n491) );
  NAND2_X1 U553 ( .A1(n448), .A2(n491), .ZN(n508) );
  NAND2_X1 U554 ( .A1(n508), .A2(G214), .ZN(n628) );
  NAND2_X1 U555 ( .A1(n597), .A2(n628), .ZN(n449) );
  XNOR2_X1 U556 ( .A(n450), .B(n449), .ZN(n552) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n451) );
  XNOR2_X1 U558 ( .A(n455), .B(n454), .ZN(n458) );
  NAND2_X1 U559 ( .A1(G234), .A2(n745), .ZN(n456) );
  XNOR2_X1 U560 ( .A(n478), .B(n460), .ZN(n750) );
  XNOR2_X1 U561 ( .A(n461), .B(n750), .ZN(n698) );
  NAND2_X1 U562 ( .A1(n698), .A2(n491), .ZN(n467) );
  XNOR2_X1 U563 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n463) );
  XNOR2_X1 U564 ( .A(G902), .B(KEYINPUT15), .ZN(n670) );
  NAND2_X1 U565 ( .A1(n670), .A2(G234), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n462), .B(KEYINPUT20), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n463), .B(n352), .ZN(n465) );
  XOR2_X1 U568 ( .A(KEYINPUT75), .B(KEYINPUT98), .Z(n464) );
  XNOR2_X1 U569 ( .A(n465), .B(n464), .ZN(n466) );
  AND2_X1 U570 ( .A1(n468), .A2(G221), .ZN(n469) );
  XNOR2_X1 U571 ( .A(n469), .B(KEYINPUT21), .ZN(n540) );
  INV_X1 U572 ( .A(n540), .ZN(n642) );
  AND2_X1 U573 ( .A1(n552), .A2(n549), .ZN(n530) );
  NAND2_X1 U574 ( .A1(n471), .A2(G217), .ZN(n473) );
  XNOR2_X1 U575 ( .A(G122), .B(KEYINPUT7), .ZN(n472) );
  XNOR2_X1 U576 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n496), .B(KEYINPUT9), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U579 ( .A1(n700), .A2(n491), .ZN(n477) );
  XNOR2_X1 U580 ( .A(n477), .B(G478), .ZN(n572) );
  INV_X1 U581 ( .A(n572), .ZN(n532) );
  XNOR2_X1 U582 ( .A(n479), .B(n478), .ZN(n482) );
  NAND2_X1 U583 ( .A1(G214), .A2(n480), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n482), .B(n481), .ZN(n490) );
  XNOR2_X2 U585 ( .A(G122), .B(G113), .ZN(n483) );
  XNOR2_X1 U586 ( .A(G143), .B(KEYINPUT11), .ZN(n484) );
  XNOR2_X1 U587 ( .A(n485), .B(n484), .ZN(n487) );
  XOR2_X1 U588 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n486) );
  XNOR2_X1 U589 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U590 ( .A(n494), .B(n488), .ZN(n489) );
  NAND2_X1 U591 ( .A1(n692), .A2(n491), .ZN(n493) );
  XNOR2_X1 U592 ( .A(KEYINPUT13), .B(G475), .ZN(n492) );
  XNOR2_X1 U593 ( .A(n493), .B(n492), .ZN(n573) );
  NOR2_X1 U594 ( .A1(n532), .A2(n573), .ZN(n604) );
  XNOR2_X1 U595 ( .A(n496), .B(KEYINPUT16), .ZN(n497) );
  XNOR2_X1 U596 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n499) );
  XNOR2_X1 U597 ( .A(G146), .B(KEYINPUT17), .ZN(n498) );
  XNOR2_X1 U598 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n501), .B(n500), .ZN(n506) );
  XNOR2_X1 U600 ( .A(G125), .B(KEYINPUT94), .ZN(n503) );
  NAND2_X1 U601 ( .A1(n745), .A2(G224), .ZN(n502) );
  XNOR2_X1 U602 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n504), .B(n517), .ZN(n505) );
  XNOR2_X1 U604 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U605 ( .A(n744), .B(n507), .ZN(n685) );
  INV_X1 U606 ( .A(n670), .ZN(n675) );
  NAND2_X1 U607 ( .A1(n508), .A2(G210), .ZN(n509) );
  XNOR2_X2 U608 ( .A(n510), .B(n509), .ZN(n570) );
  BUF_X1 U609 ( .A(n570), .Z(n579) );
  NAND2_X1 U610 ( .A1(n604), .A2(n394), .ZN(n528) );
  XNOR2_X1 U611 ( .A(n512), .B(n511), .ZN(n515) );
  NAND2_X1 U612 ( .A1(n745), .A2(G227), .ZN(n513) );
  XNOR2_X1 U613 ( .A(n513), .B(KEYINPUT77), .ZN(n514) );
  XNOR2_X1 U614 ( .A(n515), .B(n514), .ZN(n519) );
  XNOR2_X1 U615 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U616 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U617 ( .A(n751), .B(n520), .ZN(n708) );
  XNOR2_X1 U618 ( .A(KEYINPUT72), .B(G469), .ZN(n521) );
  XNOR2_X1 U619 ( .A(n521), .B(KEYINPUT71), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n524), .B(KEYINPUT14), .ZN(n655) );
  INV_X1 U621 ( .A(G952), .ZN(n681) );
  NAND2_X1 U622 ( .A1(n367), .A2(n681), .ZN(n526) );
  OR2_X1 U623 ( .A1(n367), .A2(G902), .ZN(n525) );
  AND2_X1 U624 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U625 ( .A1(n655), .A2(n527), .ZN(n585) );
  NAND2_X1 U626 ( .A1(G953), .A2(G900), .ZN(n757) );
  NAND2_X1 U627 ( .A1(n585), .A2(n757), .ZN(n538) );
  NOR2_X1 U628 ( .A1(n528), .A2(n547), .ZN(n529) );
  AND2_X1 U629 ( .A1(n530), .A2(n529), .ZN(n722) );
  INV_X1 U630 ( .A(KEYINPUT38), .ZN(n531) );
  XNOR2_X1 U631 ( .A(n570), .B(n531), .ZN(n546) );
  INV_X1 U632 ( .A(n628), .ZN(n569) );
  OR2_X2 U633 ( .A1(n546), .A2(n569), .ZN(n632) );
  INV_X1 U634 ( .A(n632), .ZN(n534) );
  NAND2_X1 U635 ( .A1(n532), .A2(n573), .ZN(n631) );
  INV_X1 U636 ( .A(n631), .ZN(n533) );
  NAND2_X1 U637 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U638 ( .A(KEYINPUT41), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n536), .B(n535), .ZN(n658) );
  INV_X1 U640 ( .A(n658), .ZN(n544) );
  INV_X1 U641 ( .A(n537), .ZN(n596) );
  INV_X1 U642 ( .A(n538), .ZN(n539) );
  AND2_X1 U643 ( .A1(n540), .A2(n539), .ZN(n558) );
  NAND2_X1 U644 ( .A1(n597), .A2(n558), .ZN(n541) );
  XNOR2_X1 U645 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n542) );
  XNOR2_X1 U646 ( .A(n543), .B(n542), .ZN(n568) );
  INV_X1 U647 ( .A(n546), .ZN(n629) );
  INV_X1 U648 ( .A(n547), .ZN(n548) );
  NAND2_X1 U649 ( .A1(n629), .A2(n548), .ZN(n550) );
  INV_X1 U650 ( .A(n640), .ZN(n549) );
  INV_X1 U651 ( .A(KEYINPUT39), .ZN(n553) );
  XNOR2_X1 U652 ( .A(n554), .B(n553), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n581), .A2(n727), .ZN(n555) );
  XNOR2_X1 U654 ( .A(n556), .B(KEYINPUT46), .ZN(n557) );
  INV_X1 U655 ( .A(n727), .ZN(n723) );
  INV_X1 U656 ( .A(n558), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n596), .A2(n559), .ZN(n561) );
  XNOR2_X1 U658 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n561), .A2(n616), .ZN(n562) );
  NOR2_X1 U660 ( .A1(n723), .A2(n562), .ZN(n563) );
  XNOR2_X1 U661 ( .A(n563), .B(KEYINPUT108), .ZN(n564) );
  NAND2_X1 U662 ( .A1(n576), .A2(n394), .ZN(n566) );
  XOR2_X1 U663 ( .A(KEYINPUT36), .B(KEYINPUT90), .Z(n565) );
  XNOR2_X1 U664 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U665 ( .A(n610), .B(KEYINPUT93), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n436), .A2(n587), .ZN(n571) );
  XNOR2_X1 U667 ( .A(n571), .B(KEYINPUT80), .ZN(n724) );
  AND2_X1 U668 ( .A1(n573), .A2(n572), .ZN(n730) );
  NOR2_X1 U669 ( .A1(n727), .A2(n730), .ZN(n633) );
  NAND2_X1 U670 ( .A1(n576), .A2(n639), .ZN(n578) );
  XOR2_X1 U671 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n577) );
  XNOR2_X1 U672 ( .A(n578), .B(n577), .ZN(n580) );
  NAND2_X1 U673 ( .A1(n580), .A2(n579), .ZN(n668) );
  NAND2_X1 U674 ( .A1(n581), .A2(n730), .ZN(n737) );
  AND2_X1 U675 ( .A1(n668), .A2(n737), .ZN(n582) );
  BUF_X2 U676 ( .A(n671), .Z(n753) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n583) );
  NAND2_X1 U678 ( .A1(G953), .A2(G898), .ZN(n584) );
  AND2_X1 U679 ( .A1(n585), .A2(n584), .ZN(n586) );
  INV_X1 U680 ( .A(KEYINPUT22), .ZN(n588) );
  NOR2_X1 U681 ( .A1(n616), .A2(n596), .ZN(n589) );
  NAND2_X1 U682 ( .A1(n595), .A2(n353), .ZN(n594) );
  XNOR2_X1 U683 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n592) );
  INV_X1 U684 ( .A(KEYINPUT67), .ZN(n591) );
  XNOR2_X1 U685 ( .A(n592), .B(n591), .ZN(n593) );
  INV_X1 U686 ( .A(n597), .ZN(n609) );
  AND2_X1 U687 ( .A1(n537), .A2(n609), .ZN(n598) );
  INV_X1 U688 ( .A(KEYINPUT107), .ZN(n599) );
  INV_X1 U689 ( .A(KEYINPUT44), .ZN(n601) );
  INV_X1 U690 ( .A(KEYINPUT34), .ZN(n602) );
  XNOR2_X1 U691 ( .A(n603), .B(n602), .ZN(n605) );
  NAND2_X1 U692 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U693 ( .A1(n607), .A2(n601), .ZN(n608) );
  NOR2_X1 U694 ( .A1(n640), .A2(n609), .ZN(n612) );
  INV_X1 U695 ( .A(n639), .ZN(n611) );
  AND2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n649) );
  INV_X1 U697 ( .A(n633), .ZN(n615) );
  NOR2_X1 U698 ( .A1(n616), .A2(n537), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n619), .B(KEYINPUT89), .ZN(n620) );
  XNOR2_X2 U700 ( .A(n621), .B(KEYINPUT45), .ZN(n672) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n677) );
  NAND2_X1 U702 ( .A1(n625), .A2(n677), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(n626), .ZN(n662) );
  NOR2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n636) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U707 ( .A(KEYINPUT119), .B(n634), .Z(n635) );
  NOR2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n637), .B(KEYINPUT120), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT50), .ZN(n646) );
  XOR2_X1 U712 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n644) );
  NAND2_X1 U713 ( .A1(n642), .A2(n537), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U716 ( .A1(n597), .A2(n647), .ZN(n648) );
  NOR2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U718 ( .A(KEYINPUT51), .B(n650), .Z(n651) );
  NOR2_X1 U719 ( .A1(n658), .A2(n651), .ZN(n652) );
  NOR2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n654), .B(KEYINPUT52), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n655), .A2(G952), .ZN(n656) );
  NOR2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n660) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n663), .B(KEYINPUT121), .ZN(n664) );
  NAND2_X1 U727 ( .A1(n664), .A2(n367), .ZN(n666) );
  XNOR2_X1 U728 ( .A(n666), .B(n665), .ZN(G75) );
  XNOR2_X1 U729 ( .A(n667), .B(G101), .ZN(G3) );
  XNOR2_X1 U730 ( .A(n668), .B(G140), .ZN(G42) );
  XNOR2_X1 U731 ( .A(n669), .B(G110), .ZN(G12) );
  NOR2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n675), .A2(KEYINPUT2), .ZN(n676) );
  NAND2_X1 U735 ( .A1(n705), .A2(G472), .ZN(n680) );
  XOR2_X1 U736 ( .A(KEYINPUT62), .B(n678), .Z(n679) );
  XNOR2_X1 U737 ( .A(n680), .B(n679), .ZN(n682) );
  NAND2_X1 U738 ( .A1(n681), .A2(G953), .ZN(n702) );
  NAND2_X1 U739 ( .A1(n682), .A2(n702), .ZN(n684) );
  XOR2_X1 U740 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n683) );
  XNOR2_X1 U741 ( .A(n684), .B(n683), .ZN(G57) );
  INV_X1 U742 ( .A(KEYINPUT56), .ZN(n691) );
  NAND2_X1 U743 ( .A1(n349), .A2(G210), .ZN(n689) );
  BUF_X1 U744 ( .A(n685), .Z(n686) );
  XNOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n690) );
  INV_X1 U747 ( .A(KEYINPUT60), .ZN(n696) );
  NAND2_X1 U748 ( .A1(n350), .A2(G475), .ZN(n694) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n350), .A2(G217), .ZN(n697) );
  XOR2_X1 U751 ( .A(n698), .B(n697), .Z(n699) );
  INV_X1 U752 ( .A(n702), .ZN(n711) );
  NOR2_X1 U753 ( .A1(n699), .A2(n711), .ZN(G66) );
  NAND2_X1 U754 ( .A1(n705), .A2(G478), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U756 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U757 ( .A(n704), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n349), .A2(G469), .ZN(n710) );
  XOR2_X1 U759 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(KEYINPUT58), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(G54) );
  NAND2_X1 U764 ( .A1(n351), .A2(n727), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(KEYINPUT112), .ZN(n714) );
  XNOR2_X1 U766 ( .A(G104), .B(n714), .ZN(G6) );
  XOR2_X1 U767 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n716) );
  NAND2_X1 U768 ( .A1(n351), .A2(n730), .ZN(n715) );
  XNOR2_X1 U769 ( .A(n716), .B(n715), .ZN(n718) );
  XOR2_X1 U770 ( .A(G107), .B(KEYINPUT26), .Z(n717) );
  XNOR2_X1 U771 ( .A(n718), .B(n717), .ZN(G9) );
  INV_X1 U772 ( .A(n730), .ZN(n719) );
  NOR2_X1 U773 ( .A1(n724), .A2(n719), .ZN(n721) );
  XNOR2_X1 U774 ( .A(G128), .B(KEYINPUT29), .ZN(n720) );
  XNOR2_X1 U775 ( .A(n721), .B(n720), .ZN(G30) );
  XOR2_X1 U776 ( .A(G143), .B(n722), .Z(G45) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U778 ( .A(KEYINPUT114), .B(n725), .Z(n726) );
  XNOR2_X1 U779 ( .A(G146), .B(n726), .ZN(G48) );
  XOR2_X1 U780 ( .A(G113), .B(KEYINPUT115), .Z(n729) );
  NAND2_X1 U781 ( .A1(n731), .A2(n727), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(G15) );
  NAND2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(G116), .ZN(G18) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT116), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n734), .B(KEYINPUT37), .ZN(n735) );
  XNOR2_X1 U787 ( .A(G125), .B(n735), .ZN(G27) );
  XOR2_X1 U788 ( .A(G134), .B(KEYINPUT117), .Z(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(G36) );
  NAND2_X1 U790 ( .A1(n623), .A2(n367), .ZN(n738) );
  XOR2_X1 U791 ( .A(KEYINPUT125), .B(n738), .Z(n743) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n739) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U794 ( .A1(n740), .A2(G898), .ZN(n741) );
  XNOR2_X1 U795 ( .A(KEYINPUT124), .B(n741), .ZN(n742) );
  NAND2_X1 U796 ( .A1(n743), .A2(n742), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n744), .B(G110), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n367), .A2(G898), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n749), .B(n748), .ZN(G69) );
  XNOR2_X1 U801 ( .A(n750), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U802 ( .A(n751), .B(n752), .ZN(n755) );
  XOR2_X1 U803 ( .A(n755), .B(n753), .Z(n754) );
  NOR2_X1 U804 ( .A1(G953), .A2(n754), .ZN(n759) );
  XNOR2_X1 U805 ( .A(n755), .B(G227), .ZN(n756) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U808 ( .A(KEYINPUT127), .B(n760), .Z(G72) );
  XNOR2_X1 U809 ( .A(G137), .B(n761), .ZN(G39) );
endmodule

