

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729;

  INV_X2 U373 ( .A(G953), .ZN(n721) );
  NOR2_X1 U374 ( .A1(G953), .A2(G237), .ZN(n475) );
  XNOR2_X1 U375 ( .A(n523), .B(n522), .ZN(n698) );
  XNOR2_X2 U376 ( .A(n415), .B(KEYINPUT19), .ZN(n550) );
  NAND2_X2 U377 ( .A1(n586), .A2(n585), .ZN(n588) );
  AND2_X1 U378 ( .A1(n521), .A2(n520), .ZN(n523) );
  NOR2_X1 U379 ( .A1(n609), .A2(n608), .ZN(n536) );
  XNOR2_X1 U380 ( .A(n474), .B(n473), .ZN(n595) );
  NOR2_X1 U381 ( .A1(n694), .A2(G902), .ZN(n474) );
  XNOR2_X1 U382 ( .A(n409), .B(G134), .ZN(n431) );
  INV_X2 U383 ( .A(G131), .ZN(n365) );
  XOR2_X1 U384 ( .A(G146), .B(G125), .Z(n438) );
  XNOR2_X1 U385 ( .A(n376), .B(KEYINPUT39), .ZN(n350) );
  BUF_X1 U386 ( .A(n647), .Z(n351) );
  NAND2_X2 U387 ( .A1(n562), .A2(n606), .ZN(n376) );
  XNOR2_X1 U388 ( .A(n535), .B(n534), .ZN(n647) );
  XNOR2_X1 U389 ( .A(n352), .B(KEYINPUT111), .ZN(n609) );
  NOR2_X1 U390 ( .A1(n532), .A2(n527), .ZN(n352) );
  XNOR2_X2 U391 ( .A(n530), .B(KEYINPUT77), .ZN(n562) );
  XNOR2_X2 U392 ( .A(n588), .B(n587), .ZN(n628) );
  XNOR2_X1 U393 ( .A(n676), .B(KEYINPUT91), .ZN(n569) );
  NOR2_X1 U394 ( .A1(n654), .A2(n505), .ZN(n521) );
  XOR2_X1 U395 ( .A(G116), .B(G122), .Z(n432) );
  AND2_X1 U396 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U397 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U398 ( .A(n463), .B(n462), .ZN(n466) );
  XOR2_X1 U399 ( .A(KEYINPUT24), .B(G110), .Z(n459) );
  XNOR2_X1 U400 ( .A(n500), .B(n499), .ZN(n359) );
  AND2_X1 U401 ( .A1(n545), .A2(n544), .ZN(n551) );
  AND2_X1 U402 ( .A1(n638), .A2(KEYINPUT2), .ZN(n378) );
  XNOR2_X1 U403 ( .A(n364), .B(n399), .ZN(n680) );
  XNOR2_X1 U404 ( .A(n712), .B(n398), .ZN(n364) );
  AND2_X1 U405 ( .A1(n564), .A2(n563), .ZN(n570) );
  XNOR2_X1 U406 ( .A(KEYINPUT5), .B(G116), .ZN(n477) );
  XNOR2_X1 U407 ( .A(G119), .B(KEYINPUT78), .ZN(n460) );
  XNOR2_X1 U408 ( .A(n395), .B(n431), .ZN(n481) );
  XNOR2_X1 U409 ( .A(KEYINPUT70), .B(G137), .ZN(n394) );
  XNOR2_X1 U410 ( .A(n711), .B(n384), .ZN(n405) );
  XNOR2_X1 U411 ( .A(n391), .B(KEYINPUT67), .ZN(n384) );
  OR2_X1 U412 ( .A1(n537), .A2(n527), .ZN(n529) );
  INV_X1 U413 ( .A(G237), .ZN(n402) );
  XNOR2_X1 U414 ( .A(n393), .B(n392), .ZN(n704) );
  XOR2_X1 U415 ( .A(G104), .B(G107), .Z(n393) );
  XNOR2_X1 U416 ( .A(G143), .B(G113), .ZN(n440) );
  XOR2_X1 U417 ( .A(G122), .B(G104), .Z(n441) );
  XNOR2_X1 U418 ( .A(n405), .B(G146), .ZN(n483) );
  XNOR2_X1 U419 ( .A(n481), .B(KEYINPUT94), .ZN(n712) );
  XNOR2_X1 U420 ( .A(n405), .B(KEYINPUT80), .ZN(n373) );
  XNOR2_X1 U421 ( .A(n407), .B(n479), .ZN(n703) );
  XNOR2_X1 U422 ( .A(n704), .B(KEYINPUT72), .ZN(n404) );
  XNOR2_X1 U423 ( .A(n631), .B(KEYINPUT87), .ZN(n715) );
  XNOR2_X1 U424 ( .A(n376), .B(KEYINPUT39), .ZN(n533) );
  XNOR2_X1 U425 ( .A(n518), .B(n517), .ZN(n655) );
  AND2_X1 U426 ( .A1(n511), .A2(n510), .ZN(n526) );
  XNOR2_X1 U427 ( .A(n423), .B(KEYINPUT0), .ZN(n424) );
  XNOR2_X1 U428 ( .A(G128), .B(G137), .ZN(n458) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n691) );
  XNOR2_X1 U430 ( .A(n436), .B(n435), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n374), .B(n372), .ZN(n649) );
  XNOR2_X1 U432 ( .A(n375), .B(n703), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n373), .B(n404), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n411), .B(n386), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n547), .B(KEYINPUT42), .ZN(n727) );
  AND2_X1 U436 ( .A1(n368), .A2(n362), .ZN(n676) );
  XNOR2_X1 U437 ( .A(n358), .B(n357), .ZN(n502) );
  INV_X1 U438 ( .A(KEYINPUT35), .ZN(n357) );
  NAND2_X1 U439 ( .A1(n359), .A2(n501), .ZN(n358) );
  NAND2_X1 U440 ( .A1(n551), .A2(n550), .ZN(n667) );
  XNOR2_X1 U441 ( .A(n683), .B(n682), .ZN(n684) );
  INV_X1 U442 ( .A(n566), .ZN(n361) );
  NOR2_X1 U443 ( .A1(n691), .A2(G902), .ZN(n353) );
  NOR2_X1 U444 ( .A1(n362), .A2(n510), .ZN(n354) );
  XOR2_X1 U445 ( .A(n640), .B(KEYINPUT62), .Z(n355) );
  XOR2_X1 U446 ( .A(n548), .B(KEYINPUT46), .Z(n356) );
  XNOR2_X1 U447 ( .A(n434), .B(n433), .ZN(n367) );
  XNOR2_X1 U448 ( .A(n369), .B(KEYINPUT36), .ZN(n368) );
  INV_X1 U449 ( .A(n502), .ZN(n728) );
  NOR2_X1 U450 ( .A1(n592), .A2(n591), .ZN(n363) );
  NAND2_X1 U451 ( .A1(n362), .A2(n360), .ZN(n497) );
  NOR2_X1 U452 ( .A1(n591), .A2(n361), .ZN(n360) );
  INV_X1 U453 ( .A(n592), .ZN(n362) );
  NAND2_X1 U454 ( .A1(n363), .A2(n541), .ZN(n506) );
  XNOR2_X2 U455 ( .A(n365), .B(KEYINPUT69), .ZN(n443) );
  AND2_X1 U456 ( .A1(n576), .A2(n580), .ZN(n369) );
  NOR2_X2 U457 ( .A1(n727), .A2(n647), .ZN(n549) );
  XNOR2_X1 U458 ( .A(n370), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U459 ( .A1(n371), .A2(n643), .ZN(n370) );
  XNOR2_X1 U460 ( .A(n641), .B(n355), .ZN(n371) );
  INV_X1 U461 ( .A(n532), .ZN(n606) );
  AND2_X1 U462 ( .A1(n383), .A2(KEYINPUT2), .ZN(n639) );
  NOR2_X1 U463 ( .A1(n382), .A2(n715), .ZN(n636) );
  NAND2_X2 U464 ( .A1(n379), .A2(n377), .ZN(n685) );
  NAND2_X1 U465 ( .A1(n383), .A2(n378), .ZN(n377) );
  NAND2_X1 U466 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X1 U467 ( .A1(n715), .A2(n637), .ZN(n380) );
  INV_X1 U468 ( .A(n382), .ZN(n381) );
  NAND2_X1 U469 ( .A1(n628), .A2(n698), .ZN(n382) );
  NAND2_X1 U470 ( .A1(n589), .A2(n698), .ZN(n383) );
  XNOR2_X2 U471 ( .A(n390), .B(KEYINPUT68), .ZN(n711) );
  AND2_X2 U472 ( .A1(n526), .A2(n540), .ZN(n388) );
  XNOR2_X1 U473 ( .A(n400), .B(G469), .ZN(n509) );
  XNOR2_X2 U474 ( .A(n414), .B(n413), .ZN(n580) );
  AND2_X1 U475 ( .A1(G227), .A2(n721), .ZN(n385) );
  XOR2_X1 U476 ( .A(n438), .B(n403), .Z(n386) );
  XOR2_X1 U477 ( .A(n529), .B(n528), .Z(n387) );
  NOR2_X1 U478 ( .A1(KEYINPUT84), .A2(n667), .ZN(n389) );
  OR2_X1 U479 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U480 ( .A(KEYINPUT92), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n504), .B(KEYINPUT44), .ZN(n505) );
  XNOR2_X1 U482 ( .A(n397), .B(n385), .ZN(n398) );
  XNOR2_X1 U483 ( .A(n432), .B(KEYINPUT16), .ZN(n407) );
  NAND2_X1 U484 ( .A1(n541), .A2(n565), .ZN(n543) );
  XNOR2_X1 U485 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U486 ( .A(KEYINPUT34), .ZN(n499) );
  INV_X1 U487 ( .A(n697), .ZN(n643) );
  XNOR2_X1 U488 ( .A(n680), .B(n681), .ZN(n682) );
  XNOR2_X1 U489 ( .A(n635), .B(n634), .ZN(G75) );
  XNOR2_X2 U490 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n390) );
  INV_X1 U491 ( .A(G101), .ZN(n391) );
  XNOR2_X1 U492 ( .A(KEYINPUT93), .B(G110), .ZN(n392) );
  XNOR2_X1 U493 ( .A(n483), .B(n404), .ZN(n399) );
  XNOR2_X2 U494 ( .A(G143), .B(G128), .ZN(n409) );
  XNOR2_X1 U495 ( .A(n443), .B(n394), .ZN(n395) );
  XNOR2_X1 U496 ( .A(G140), .B(KEYINPUT95), .ZN(n396) );
  XNOR2_X1 U497 ( .A(n396), .B(KEYINPUT79), .ZN(n397) );
  NOR2_X1 U498 ( .A1(n680), .A2(G902), .ZN(n400) );
  INV_X1 U499 ( .A(n509), .ZN(n545) );
  INV_X1 U500 ( .A(KEYINPUT1), .ZN(n401) );
  XNOR2_X2 U501 ( .A(n545), .B(n401), .ZN(n592) );
  INV_X1 U502 ( .A(G902), .ZN(n417) );
  NAND2_X1 U503 ( .A1(n417), .A2(n402), .ZN(n412) );
  NAND2_X1 U504 ( .A1(n412), .A2(G214), .ZN(n605) );
  XOR2_X1 U505 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n403) );
  XNOR2_X1 U506 ( .A(KEYINPUT3), .B(G119), .ZN(n406) );
  XNOR2_X1 U507 ( .A(n406), .B(G113), .ZN(n479) );
  NAND2_X1 U508 ( .A1(G224), .A2(n721), .ZN(n408) );
  XNOR2_X1 U509 ( .A(n408), .B(KEYINPUT81), .ZN(n410) );
  XNOR2_X1 U510 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U511 ( .A(KEYINPUT15), .B(G902), .ZN(n637) );
  NAND2_X1 U512 ( .A1(n649), .A2(n637), .ZN(n414) );
  AND2_X1 U513 ( .A1(n412), .A2(G210), .ZN(n413) );
  NAND2_X1 U514 ( .A1(n605), .A2(n580), .ZN(n415) );
  NAND2_X1 U515 ( .A1(G234), .A2(G237), .ZN(n416) );
  XNOR2_X1 U516 ( .A(n416), .B(KEYINPUT14), .ZN(n620) );
  NAND2_X1 U517 ( .A1(G953), .A2(n417), .ZN(n418) );
  NAND2_X1 U518 ( .A1(n620), .A2(n418), .ZN(n420) );
  NOR2_X1 U519 ( .A1(G953), .A2(G952), .ZN(n419) );
  NOR2_X1 U520 ( .A1(n420), .A2(n419), .ZN(n525) );
  NAND2_X1 U521 ( .A1(G898), .A2(G953), .ZN(n421) );
  AND2_X1 U522 ( .A1(n525), .A2(n421), .ZN(n422) );
  NAND2_X1 U523 ( .A1(n550), .A2(n422), .ZN(n425) );
  XNOR2_X2 U524 ( .A(n425), .B(n424), .ZN(n512) );
  XOR2_X1 U525 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n428) );
  NAND2_X1 U526 ( .A1(n637), .A2(G234), .ZN(n426) );
  XNOR2_X1 U527 ( .A(n426), .B(KEYINPUT20), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(G221), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n428), .B(n427), .ZN(n538) );
  INV_X1 U530 ( .A(n538), .ZN(n594) );
  XNOR2_X1 U531 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n430) );
  NAND2_X1 U532 ( .A1(G234), .A2(n721), .ZN(n429) );
  XNOR2_X1 U533 ( .A(n430), .B(n429), .ZN(n464) );
  NAND2_X1 U534 ( .A1(n464), .A2(G217), .ZN(n436) );
  XNOR2_X1 U535 ( .A(n431), .B(G107), .ZN(n434) );
  XOR2_X1 U536 ( .A(KEYINPUT7), .B(n432), .Z(n433) );
  XOR2_X1 U537 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n435) );
  XNOR2_X1 U538 ( .A(KEYINPUT104), .B(G478), .ZN(n437) );
  XNOR2_X1 U539 ( .A(n353), .B(n437), .ZN(n516) );
  XNOR2_X1 U540 ( .A(KEYINPUT13), .B(G475), .ZN(n451) );
  XNOR2_X1 U541 ( .A(G140), .B(n438), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n439), .B(KEYINPUT10), .ZN(n713) );
  XNOR2_X1 U543 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U544 ( .A(n713), .B(n442), .ZN(n449) );
  XNOR2_X1 U545 ( .A(n443), .B(KEYINPUT12), .ZN(n447) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n445) );
  NAND2_X1 U547 ( .A1(G214), .A2(n475), .ZN(n444) );
  XNOR2_X1 U548 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U549 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U550 ( .A(n449), .B(n448), .ZN(n686) );
  NOR2_X1 U551 ( .A1(G902), .A2(n686), .ZN(n450) );
  XNOR2_X1 U552 ( .A(n451), .B(n450), .ZN(n515) );
  INV_X1 U553 ( .A(n515), .ZN(n452) );
  NAND2_X1 U554 ( .A1(n516), .A2(n452), .ZN(n453) );
  XNOR2_X1 U555 ( .A(KEYINPUT106), .B(n453), .ZN(n608) );
  NOR2_X1 U556 ( .A1(n594), .A2(n608), .ZN(n454) );
  NAND2_X1 U557 ( .A1(n512), .A2(n454), .ZN(n457) );
  XNOR2_X1 U558 ( .A(KEYINPUT22), .B(KEYINPUT75), .ZN(n455) );
  XNOR2_X1 U559 ( .A(n455), .B(KEYINPUT66), .ZN(n456) );
  XNOR2_X2 U560 ( .A(n457), .B(n456), .ZN(n493) );
  NAND2_X1 U561 ( .A1(n592), .A2(n493), .ZN(n488) );
  XNOR2_X1 U562 ( .A(n459), .B(n458), .ZN(n469) );
  XOR2_X1 U563 ( .A(KEYINPUT96), .B(KEYINPUT23), .Z(n461) );
  XNOR2_X1 U564 ( .A(n461), .B(n460), .ZN(n463) );
  XOR2_X1 U565 ( .A(KEYINPUT71), .B(KEYINPUT97), .Z(n462) );
  NAND2_X1 U566 ( .A1(n464), .A2(G221), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n467), .B(n713), .ZN(n468) );
  XNOR2_X1 U568 ( .A(n469), .B(n468), .ZN(n694) );
  NAND2_X1 U569 ( .A1(n470), .A2(G217), .ZN(n472) );
  INV_X1 U570 ( .A(KEYINPUT25), .ZN(n471) );
  INV_X1 U571 ( .A(n595), .ZN(n510) );
  NAND2_X1 U572 ( .A1(G210), .A2(n475), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U574 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U575 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U576 ( .A(n483), .B(n482), .ZN(n640) );
  OR2_X1 U577 ( .A1(n640), .A2(G902), .ZN(n486) );
  INV_X1 U578 ( .A(KEYINPUT74), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n484), .B(G472), .ZN(n485) );
  XNOR2_X2 U580 ( .A(n486), .B(n485), .ZN(n537) );
  XNOR2_X1 U581 ( .A(n537), .B(KEYINPUT6), .ZN(n566) );
  NAND2_X1 U582 ( .A1(n510), .A2(n361), .ZN(n487) );
  NOR2_X1 U583 ( .A1(n488), .A2(n487), .ZN(n654) );
  AND2_X1 U584 ( .A1(n595), .A2(n361), .ZN(n489) );
  AND2_X1 U585 ( .A1(n362), .A2(n489), .ZN(n490) );
  NAND2_X1 U586 ( .A1(n493), .A2(n490), .ZN(n492) );
  XOR2_X1 U587 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n491) );
  XNOR2_X1 U588 ( .A(n492), .B(n491), .ZN(n729) );
  AND2_X1 U589 ( .A1(n354), .A2(n493), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n494), .A2(n537), .ZN(n646) );
  AND2_X1 U591 ( .A1(n729), .A2(n646), .ZN(n503) );
  INV_X1 U592 ( .A(n516), .ZN(n495) );
  NAND2_X1 U593 ( .A1(n515), .A2(n495), .ZN(n496) );
  XNOR2_X1 U594 ( .A(KEYINPUT107), .B(n496), .ZN(n560) );
  XNOR2_X1 U595 ( .A(n560), .B(KEYINPUT82), .ZN(n501) );
  XOR2_X1 U596 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n498) );
  NAND2_X1 U597 ( .A1(n510), .A2(n538), .ZN(n591) );
  XNOR2_X1 U598 ( .A(n498), .B(n497), .ZN(n613) );
  NAND2_X1 U599 ( .A1(n512), .A2(n613), .ZN(n500) );
  NAND2_X1 U600 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U601 ( .A(KEYINPUT100), .B(n506), .Z(n602) );
  NAND2_X1 U602 ( .A1(n602), .A2(n512), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n507), .B(KEYINPUT101), .ZN(n508) );
  XNOR2_X1 U604 ( .A(KEYINPUT31), .B(n508), .ZN(n673) );
  NOR2_X1 U605 ( .A1(n509), .A2(n594), .ZN(n511) );
  NAND2_X1 U606 ( .A1(n526), .A2(n512), .ZN(n513) );
  XNOR2_X1 U607 ( .A(KEYINPUT99), .B(n513), .ZN(n514) );
  NAND2_X1 U608 ( .A1(n514), .A2(n537), .ZN(n662) );
  NAND2_X1 U609 ( .A1(n673), .A2(n662), .ZN(n519) );
  NOR2_X1 U610 ( .A1(n516), .A2(n515), .ZN(n661) );
  AND2_X1 U611 ( .A1(n516), .A2(n515), .ZN(n518) );
  INV_X1 U612 ( .A(KEYINPUT105), .ZN(n517) );
  NOR2_X1 U613 ( .A1(n661), .A2(n655), .ZN(n610) );
  INV_X1 U614 ( .A(n610), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n519), .A2(n552), .ZN(n520) );
  XOR2_X1 U616 ( .A(KEYINPUT88), .B(KEYINPUT45), .Z(n522) );
  NAND2_X1 U617 ( .A1(G953), .A2(G900), .ZN(n524) );
  AND2_X1 U618 ( .A1(n525), .A2(n524), .ZN(n540) );
  INV_X1 U619 ( .A(n605), .ZN(n527) );
  XNOR2_X1 U620 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n528) );
  NAND2_X1 U621 ( .A1(n388), .A2(n387), .ZN(n530) );
  XNOR2_X1 U622 ( .A(KEYINPUT76), .B(KEYINPUT38), .ZN(n531) );
  XNOR2_X1 U623 ( .A(n580), .B(n531), .ZN(n532) );
  NAND2_X1 U624 ( .A1(n533), .A2(n655), .ZN(n535) );
  INV_X1 U625 ( .A(KEYINPUT40), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n536), .B(KEYINPUT41), .ZN(n590) );
  INV_X1 U627 ( .A(n537), .ZN(n541) );
  AND2_X1 U628 ( .A1(n538), .A2(n595), .ZN(n539) );
  AND2_X1 U629 ( .A1(n540), .A2(n539), .ZN(n565) );
  INV_X1 U630 ( .A(KEYINPUT28), .ZN(n542) );
  XNOR2_X1 U631 ( .A(n543), .B(n542), .ZN(n544) );
  INV_X1 U632 ( .A(n551), .ZN(n546) );
  NOR2_X1 U633 ( .A1(n590), .A2(n546), .ZN(n547) );
  INV_X1 U634 ( .A(KEYINPUT90), .ZN(n548) );
  XNOR2_X1 U635 ( .A(n549), .B(n356), .ZN(n572) );
  NAND2_X1 U636 ( .A1(KEYINPUT84), .A2(n667), .ZN(n553) );
  AND2_X1 U637 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U638 ( .A1(n554), .A2(KEYINPUT47), .ZN(n559) );
  NOR2_X1 U639 ( .A1(n667), .A2(n610), .ZN(n557) );
  INV_X1 U640 ( .A(KEYINPUT47), .ZN(n555) );
  NAND2_X1 U641 ( .A1(n555), .A2(KEYINPUT84), .ZN(n556) );
  NAND2_X1 U642 ( .A1(n559), .A2(n558), .ZN(n564) );
  AND2_X1 U643 ( .A1(n560), .A2(n580), .ZN(n561) );
  AND2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n644) );
  NOR2_X1 U645 ( .A1(n389), .A2(n644), .ZN(n563) );
  NAND2_X1 U646 ( .A1(n655), .A2(n565), .ZN(n568) );
  NAND2_X1 U647 ( .A1(n566), .A2(n605), .ZN(n567) );
  NOR2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X2 U650 ( .A(n573), .B(KEYINPUT48), .ZN(n630) );
  INV_X1 U651 ( .A(n630), .ZN(n586) );
  AND2_X1 U652 ( .A1(n350), .A2(n661), .ZN(n645) );
  INV_X1 U653 ( .A(n645), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n574), .A2(KEYINPUT2), .ZN(n575) );
  XNOR2_X1 U655 ( .A(n575), .B(KEYINPUT83), .ZN(n584) );
  XOR2_X1 U656 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n578) );
  NAND2_X1 U657 ( .A1(n576), .A2(n592), .ZN(n577) );
  XNOR2_X1 U658 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U659 ( .A(n579), .B(KEYINPUT43), .ZN(n582) );
  INV_X1 U660 ( .A(n580), .ZN(n581) );
  AND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n679) );
  INV_X1 U662 ( .A(n679), .ZN(n583) );
  AND2_X1 U663 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U664 ( .A(KEYINPUT89), .ZN(n587) );
  INV_X1 U665 ( .A(n628), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT50), .B(n593), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n597) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n600), .A2(n541), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT51), .B(n603), .Z(n604) );
  NOR2_X1 U675 ( .A1(n590), .A2(n604), .ZN(n617) );
  NOR2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n612) );
  NOR2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U680 ( .A(n613), .ZN(n623) );
  NOR2_X1 U681 ( .A1(n614), .A2(n623), .ZN(n615) );
  XOR2_X1 U682 ( .A(KEYINPUT119), .B(n615), .Z(n616) );
  NOR2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U684 ( .A(KEYINPUT52), .B(n618), .Z(n619) );
  XOR2_X1 U685 ( .A(KEYINPUT120), .B(n619), .Z(n622) );
  NAND2_X1 U686 ( .A1(n620), .A2(G952), .ZN(n621) );
  OR2_X1 U687 ( .A1(n622), .A2(n621), .ZN(n626) );
  NOR2_X1 U688 ( .A1(n590), .A2(n623), .ZN(n624) );
  NOR2_X1 U689 ( .A1(G953), .A2(n624), .ZN(n625) );
  NAND2_X1 U690 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U691 ( .A1(n639), .A2(n627), .ZN(n632) );
  OR2_X1 U692 ( .A1(n645), .A2(n679), .ZN(n629) );
  NOR2_X1 U693 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U694 ( .A1(n632), .A2(n636), .ZN(n635) );
  INV_X1 U695 ( .A(KEYINPUT53), .ZN(n633) );
  XNOR2_X1 U696 ( .A(n633), .B(KEYINPUT121), .ZN(n634) );
  XOR2_X1 U697 ( .A(KEYINPUT86), .B(n637), .Z(n638) );
  NAND2_X1 U698 ( .A1(n685), .A2(G472), .ZN(n641) );
  INV_X1 U699 ( .A(G952), .ZN(n642) );
  AND2_X1 U700 ( .A1(n642), .A2(G953), .ZN(n697) );
  XOR2_X1 U701 ( .A(G143), .B(n644), .Z(G45) );
  XOR2_X1 U702 ( .A(G134), .B(n645), .Z(G36) );
  XNOR2_X1 U703 ( .A(n646), .B(G110), .ZN(G12) );
  XOR2_X1 U704 ( .A(G131), .B(n351), .Z(G33) );
  NAND2_X1 U705 ( .A1(n685), .A2(G210), .ZN(n651) );
  XNOR2_X1 U706 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n648) );
  XNOR2_X1 U707 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U708 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X2 U709 ( .A1(n652), .A2(n697), .ZN(n653) );
  XNOR2_X1 U710 ( .A(n653), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U711 ( .A(G101), .B(n654), .Z(G3) );
  INV_X1 U712 ( .A(n655), .ZN(n670) );
  NOR2_X1 U713 ( .A1(n662), .A2(n670), .ZN(n657) );
  XNOR2_X1 U714 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n656) );
  XNOR2_X1 U715 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U716 ( .A(G104), .B(n658), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n660) );
  XNOR2_X1 U718 ( .A(G107), .B(KEYINPUT26), .ZN(n659) );
  XNOR2_X1 U719 ( .A(n660), .B(n659), .ZN(n664) );
  INV_X1 U720 ( .A(n661), .ZN(n674) );
  NOR2_X1 U721 ( .A1(n662), .A2(n674), .ZN(n663) );
  XOR2_X1 U722 ( .A(n664), .B(n663), .Z(G9) );
  NOR2_X1 U723 ( .A1(n674), .A2(n667), .ZN(n666) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .ZN(n665) );
  XNOR2_X1 U725 ( .A(n666), .B(n665), .ZN(G30) );
  NOR2_X1 U726 ( .A1(n670), .A2(n667), .ZN(n669) );
  XNOR2_X1 U727 ( .A(G146), .B(KEYINPUT115), .ZN(n668) );
  XNOR2_X1 U728 ( .A(n669), .B(n668), .ZN(G48) );
  NOR2_X1 U729 ( .A1(n670), .A2(n673), .ZN(n671) );
  XOR2_X1 U730 ( .A(KEYINPUT116), .B(n671), .Z(n672) );
  XNOR2_X1 U731 ( .A(G113), .B(n672), .ZN(G15) );
  NOR2_X1 U732 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U733 ( .A(G116), .B(n675), .Z(G18) );
  XOR2_X1 U734 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n678) );
  XNOR2_X1 U735 ( .A(G125), .B(n676), .ZN(n677) );
  XNOR2_X1 U736 ( .A(n678), .B(n677), .ZN(G27) );
  XOR2_X1 U737 ( .A(G140), .B(n679), .Z(G42) );
  NAND2_X1 U738 ( .A1(n685), .A2(G469), .ZN(n683) );
  XOR2_X1 U739 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  NOR2_X1 U740 ( .A1(n697), .A2(n684), .ZN(G54) );
  NAND2_X1 U741 ( .A1(n685), .A2(G475), .ZN(n688) );
  XOR2_X1 U742 ( .A(n686), .B(KEYINPUT59), .Z(n687) );
  XNOR2_X1 U743 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X2 U744 ( .A1(n689), .A2(n697), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n685), .A2(G478), .ZN(n692) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n697), .A2(n693), .ZN(G63) );
  NAND2_X1 U749 ( .A1(n685), .A2(G217), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U751 ( .A1(n697), .A2(n696), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n721), .A2(n698), .ZN(n702) );
  NAND2_X1 U753 ( .A1(G953), .A2(G224), .ZN(n699) );
  XNOR2_X1 U754 ( .A(KEYINPUT61), .B(n699), .ZN(n700) );
  NAND2_X1 U755 ( .A1(n700), .A2(G898), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n710) );
  XOR2_X1 U757 ( .A(KEYINPUT122), .B(n703), .Z(n706) );
  XNOR2_X1 U758 ( .A(G101), .B(n704), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U760 ( .A1(G898), .A2(n721), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(G69) );
  XNOR2_X1 U763 ( .A(n712), .B(n711), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(n717) );
  XOR2_X1 U765 ( .A(n717), .B(n715), .Z(n716) );
  NOR2_X1 U766 ( .A1(G953), .A2(n716), .ZN(n724) );
  XNOR2_X1 U767 ( .A(G227), .B(n717), .ZN(n718) );
  NAND2_X1 U768 ( .A1(n718), .A2(G900), .ZN(n719) );
  XNOR2_X1 U769 ( .A(KEYINPUT123), .B(n719), .ZN(n720) );
  NOR2_X1 U770 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n722), .B(KEYINPUT124), .ZN(n723) );
  NOR2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U773 ( .A(KEYINPUT125), .B(n725), .ZN(G72) );
  XOR2_X1 U774 ( .A(G137), .B(KEYINPUT126), .Z(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(G39) );
  XOR2_X1 U776 ( .A(n728), .B(G122), .Z(G24) );
  XNOR2_X1 U777 ( .A(G119), .B(n729), .ZN(G21) );
endmodule

