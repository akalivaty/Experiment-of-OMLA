

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XOR2_X2 U324 ( .A(G92GAT), .B(G64GAT), .Z(n390) );
  INV_X1 U325 ( .A(n553), .ZN(n504) );
  XOR2_X2 U326 ( .A(KEYINPUT41), .B(n459), .Z(n564) );
  XNOR2_X1 U327 ( .A(n455), .B(n454), .ZN(n506) );
  XOR2_X1 U328 ( .A(n398), .B(n397), .Z(n553) );
  XNOR2_X1 U329 ( .A(n525), .B(n524), .ZN(n555) );
  XOR2_X1 U330 ( .A(n422), .B(n438), .Z(n292) );
  XNOR2_X1 U331 ( .A(n301), .B(KEYINPUT21), .ZN(n302) );
  XNOR2_X1 U332 ( .A(n303), .B(n302), .ZN(n305) );
  XNOR2_X1 U333 ( .A(n391), .B(G8GAT), .ZN(n392) );
  XNOR2_X1 U334 ( .A(n523), .B(KEYINPUT64), .ZN(n524) );
  XNOR2_X1 U335 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U336 ( .A(n329), .B(n328), .ZN(n330) );
  AND2_X1 U337 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U338 ( .A(n398), .B(n387), .Z(n561) );
  XNOR2_X1 U339 ( .A(n456), .B(G106GAT), .ZN(n457) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(G1339GAT) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U342 ( .A(G22GAT), .B(G155GAT), .Z(n434) );
  XNOR2_X1 U343 ( .A(n428), .B(n434), .ZN(n294) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(G78GAT), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n293), .B(G148GAT), .ZN(n325) );
  XNOR2_X1 U346 ( .A(n294), .B(n325), .ZN(n300) );
  XOR2_X1 U347 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n296) );
  XNOR2_X1 U348 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n362) );
  XOR2_X1 U350 ( .A(n362), .B(KEYINPUT23), .Z(n298) );
  NAND2_X1 U351 ( .A1(G228GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n310) );
  XNOR2_X1 U354 ( .A(G211GAT), .B(G218GAT), .ZN(n303) );
  INV_X1 U355 ( .A(KEYINPUT89), .ZN(n301) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n393) );
  XOR2_X1 U358 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n307) );
  XNOR2_X1 U359 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n393), .B(n308), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n557) );
  XNOR2_X1 U363 ( .A(n557), .B(KEYINPUT28), .ZN(n499) );
  INV_X1 U364 ( .A(n499), .ZN(n486) );
  INV_X1 U365 ( .A(KEYINPUT110), .ZN(n455) );
  INV_X1 U366 ( .A(KEYINPUT75), .ZN(n311) );
  NAND2_X1 U367 ( .A1(KEYINPUT77), .A2(n311), .ZN(n314) );
  INV_X1 U368 ( .A(KEYINPUT77), .ZN(n312) );
  NAND2_X1 U369 ( .A1(n312), .A2(KEYINPUT75), .ZN(n313) );
  NAND2_X1 U370 ( .A1(n314), .A2(n313), .ZN(n316) );
  XNOR2_X1 U371 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n315) );
  XOR2_X1 U372 ( .A(n316), .B(n315), .Z(n317) );
  XNOR2_X1 U373 ( .A(n317), .B(n390), .ZN(n319) );
  XNOR2_X1 U374 ( .A(G176GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U376 ( .A(G85GAT), .B(KEYINPUT78), .Z(n422) );
  XNOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n320), .B(KEYINPUT74), .ZN(n438) );
  NAND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n292), .B(n321), .ZN(n322) );
  XOR2_X1 U381 ( .A(n323), .B(n322), .Z(n331) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G71GAT), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n324), .B(G120GAT), .ZN(n376) );
  XNOR2_X1 U384 ( .A(n376), .B(n325), .ZN(n329) );
  XOR2_X1 U385 ( .A(KEYINPUT33), .B(KEYINPUT80), .Z(n327) );
  XNOR2_X1 U386 ( .A(KEYINPUT79), .B(KEYINPUT76), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X2 U388 ( .A(n331), .B(n330), .ZN(n459) );
  INV_X1 U389 ( .A(n564), .ZN(n508) );
  XOR2_X1 U390 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n333) );
  XNOR2_X1 U391 ( .A(KEYINPUT68), .B(KEYINPUT73), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n351) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(G197GAT), .Z(n335) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G22GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U396 ( .A(G43GAT), .B(G36GAT), .Z(n337) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G50GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n349) );
  XOR2_X1 U400 ( .A(G113GAT), .B(G15GAT), .Z(n384) );
  XNOR2_X1 U401 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n340), .B(G8GAT), .ZN(n435) );
  XOR2_X1 U403 ( .A(n384), .B(n435), .Z(n342) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U406 ( .A(n343), .B(KEYINPUT72), .Z(n347) );
  XOR2_X1 U407 ( .A(G29GAT), .B(KEYINPUT7), .Z(n345) );
  XNOR2_X1 U408 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n429) );
  XNOR2_X1 U410 ( .A(n429), .B(KEYINPUT69), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n519) );
  INV_X1 U414 ( .A(n519), .ZN(n579) );
  NOR2_X1 U415 ( .A1(n508), .A2(n579), .ZN(n490) );
  XOR2_X1 U416 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n353) );
  XNOR2_X1 U417 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n370) );
  XOR2_X1 U419 ( .A(G85GAT), .B(G162GAT), .Z(n355) );
  XNOR2_X1 U420 ( .A(G29GAT), .B(G134GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U422 ( .A(G148GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U423 ( .A(G113GAT), .B(G120GAT), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U425 ( .A(n359), .B(n358), .Z(n368) );
  XOR2_X1 U426 ( .A(G57GAT), .B(KEYINPUT93), .Z(n361) );
  XNOR2_X1 U427 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U429 ( .A(KEYINPUT0), .B(G127GAT), .Z(n383) );
  XOR2_X1 U430 ( .A(n362), .B(n383), .Z(n364) );
  NAND2_X1 U431 ( .A1(G225GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n575) );
  XOR2_X1 U436 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n372) );
  XNOR2_X1 U437 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U439 ( .A(n373), .B(G183GAT), .Z(n375) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(G176GAT), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n398) );
  XOR2_X1 U442 ( .A(G43GAT), .B(G134GAT), .Z(n423) );
  XOR2_X1 U443 ( .A(n423), .B(n376), .Z(n378) );
  NAND2_X1 U444 ( .A1(G227GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U446 ( .A(KEYINPUT85), .B(KEYINPUT65), .Z(n380) );
  XNOR2_X1 U447 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U449 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U452 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n389) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U455 ( .A(KEYINPUT94), .B(n390), .Z(n391) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G190GAT), .ZN(n426) );
  XNOR2_X1 U458 ( .A(n396), .B(n426), .ZN(n397) );
  NAND2_X1 U459 ( .A1(n561), .A2(n504), .ZN(n399) );
  XOR2_X1 U460 ( .A(KEYINPUT99), .B(n399), .Z(n400) );
  NAND2_X1 U461 ( .A1(n557), .A2(n400), .ZN(n401) );
  XOR2_X1 U462 ( .A(KEYINPUT25), .B(n401), .Z(n406) );
  NOR2_X1 U463 ( .A1(n557), .A2(n561), .ZN(n404) );
  XOR2_X1 U464 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n402) );
  XNOR2_X1 U465 ( .A(KEYINPUT97), .B(n402), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n577) );
  XOR2_X1 U467 ( .A(n553), .B(KEYINPUT27), .Z(n409) );
  NAND2_X1 U468 ( .A1(n577), .A2(n409), .ZN(n405) );
  NAND2_X1 U469 ( .A1(n406), .A2(n405), .ZN(n407) );
  NAND2_X1 U470 ( .A1(n575), .A2(n407), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n408), .B(KEYINPUT100), .ZN(n412) );
  INV_X1 U472 ( .A(n561), .ZN(n495) );
  XOR2_X1 U473 ( .A(n495), .B(KEYINPUT87), .Z(n410) );
  INV_X1 U474 ( .A(n575), .ZN(n502) );
  NAND2_X1 U475 ( .A1(n502), .A2(n409), .ZN(n540) );
  NOR2_X1 U476 ( .A1(n486), .A2(n540), .ZN(n526) );
  NAND2_X1 U477 ( .A1(n410), .A2(n526), .ZN(n411) );
  NAND2_X1 U478 ( .A1(n412), .A2(n411), .ZN(n463) );
  XOR2_X1 U479 ( .A(G92GAT), .B(G106GAT), .Z(n414) );
  NAND2_X1 U480 ( .A1(G232GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U482 ( .A(G99GAT), .B(n415), .ZN(n433) );
  XOR2_X1 U483 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n417) );
  XNOR2_X1 U484 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U486 ( .A(KEYINPUT66), .B(KEYINPUT82), .Z(n419) );
  XNOR2_X1 U487 ( .A(KEYINPUT81), .B(KEYINPUT83), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U489 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U495 ( .A(n433), .B(n432), .Z(n460) );
  INV_X1 U496 ( .A(n460), .ZN(n570) );
  XOR2_X1 U497 ( .A(KEYINPUT36), .B(n570), .Z(n590) );
  XOR2_X1 U498 ( .A(n434), .B(G183GAT), .Z(n437) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n442) );
  XOR2_X1 U501 ( .A(n438), .B(KEYINPUT15), .Z(n440) );
  NAND2_X1 U502 ( .A1(G231GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U504 ( .A(n442), .B(n441), .Z(n450) );
  XOR2_X1 U505 ( .A(G78GAT), .B(G211GAT), .Z(n444) );
  XNOR2_X1 U506 ( .A(G127GAT), .B(G71GAT), .ZN(n443) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U508 ( .A(KEYINPUT14), .B(KEYINPUT84), .Z(n446) );
  XNOR2_X1 U509 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U511 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U512 ( .A(n450), .B(n449), .Z(n515) );
  INV_X1 U513 ( .A(n515), .ZN(n586) );
  NOR2_X1 U514 ( .A1(n590), .A2(n586), .ZN(n451) );
  NAND2_X1 U515 ( .A1(n463), .A2(n451), .ZN(n452) );
  XNOR2_X1 U516 ( .A(KEYINPUT37), .B(n452), .ZN(n453) );
  XOR2_X1 U517 ( .A(KEYINPUT105), .B(n453), .Z(n475) );
  NAND2_X1 U518 ( .A1(n490), .A2(n475), .ZN(n454) );
  NAND2_X1 U519 ( .A1(n486), .A2(n506), .ZN(n458) );
  XOR2_X1 U520 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n456) );
  NOR2_X1 U521 ( .A1(n519), .A2(n459), .ZN(n474) );
  NAND2_X1 U522 ( .A1(n586), .A2(n460), .ZN(n461) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n461), .Z(n462) );
  AND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n489) );
  NAND2_X1 U525 ( .A1(n474), .A2(n489), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n575), .A2(n471), .ZN(n464) );
  XOR2_X1 U527 ( .A(KEYINPUT34), .B(n464), .Z(n465) );
  XNOR2_X1 U528 ( .A(G1GAT), .B(n465), .ZN(G1324GAT) );
  NOR2_X1 U529 ( .A1(n553), .A2(n471), .ZN(n466) );
  XOR2_X1 U530 ( .A(G8GAT), .B(n466), .Z(G1325GAT) );
  NOR2_X1 U531 ( .A1(n471), .A2(n495), .ZN(n470) );
  XOR2_X1 U532 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n468) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n467) );
  XNOR2_X1 U534 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U535 ( .A(n470), .B(n469), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n499), .A2(n471), .ZN(n473) );
  XNOR2_X1 U537 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n472) );
  XNOR2_X1 U538 ( .A(n473), .B(n472), .ZN(G1327GAT) );
  INV_X1 U539 ( .A(KEYINPUT38), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n487) );
  NAND2_X1 U542 ( .A1(n502), .A2(n487), .ZN(n479) );
  XOR2_X1 U543 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n478) );
  XNOR2_X1 U544 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n480), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n482) );
  NAND2_X1 U547 ( .A1(n504), .A2(n487), .ZN(n481) );
  XNOR2_X1 U548 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U549 ( .A(G36GAT), .B(n483), .ZN(G1329GAT) );
  NAND2_X1 U550 ( .A1(n487), .A2(n561), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n484), .B(KEYINPUT40), .ZN(n485) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n485), .ZN(G1330GAT) );
  NAND2_X1 U553 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n488), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U555 ( .A1(n490), .A2(n489), .ZN(n498) );
  NOR2_X1 U556 ( .A1(n575), .A2(n498), .ZN(n492) );
  XNOR2_X1 U557 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U559 ( .A(G57GAT), .B(n493), .Z(G1332GAT) );
  NOR2_X1 U560 ( .A1(n553), .A2(n498), .ZN(n494) );
  XOR2_X1 U561 ( .A(G64GAT), .B(n494), .Z(G1333GAT) );
  NOR2_X1 U562 ( .A1(n495), .A2(n498), .ZN(n497) );
  XNOR2_X1 U563 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n497), .B(n496), .ZN(G1334GAT) );
  NOR2_X1 U565 ( .A1(n499), .A2(n498), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(G1335GAT) );
  NAND2_X1 U568 ( .A1(n502), .A2(n506), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G85GAT), .B(n503), .ZN(G1336GAT) );
  NAND2_X1 U570 ( .A1(n506), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U572 ( .A1(n506), .A2(n561), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n529) );
  NOR2_X1 U575 ( .A1(n508), .A2(n519), .ZN(n510) );
  XNOR2_X1 U576 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(n511) );
  NOR2_X1 U578 ( .A1(n511), .A2(n586), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(KEYINPUT113), .ZN(n513) );
  NOR2_X1 U580 ( .A1(n570), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT47), .ZN(n522) );
  NOR2_X1 U582 ( .A1(n590), .A2(n515), .ZN(n516) );
  XOR2_X1 U583 ( .A(KEYINPUT45), .B(n516), .Z(n517) );
  NOR2_X1 U584 ( .A1(n459), .A2(n517), .ZN(n518) );
  XNOR2_X1 U585 ( .A(KEYINPUT114), .B(n518), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n525) );
  INV_X1 U588 ( .A(KEYINPUT48), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n561), .A2(n526), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n555), .A2(n527), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n536), .A2(n579), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U595 ( .A1(n536), .A2(n564), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U598 ( .A1(n536), .A2(n586), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U602 ( .A1(n536), .A2(n570), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n555), .A2(n540), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n541), .A2(n577), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT119), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n579), .A2(n550), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT120), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U612 ( .A1(n550), .A2(n564), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT121), .Z(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n586), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n550), .A2(n570), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT122), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  XOR2_X1 U621 ( .A(n553), .B(KEYINPUT123), .Z(n554) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT54), .ZN(n574) );
  AND2_X1 U624 ( .A1(n575), .A2(n557), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n574), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT55), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT124), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n571), .A2(n579), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n566) );
  NAND2_X1 U631 ( .A1(n571), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n567), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT125), .Z(n569) );
  NAND2_X1 U635 ( .A1(n586), .A2(n571), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT58), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n573), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(n578), .ZN(n589) );
  INV_X1 U644 ( .A(n589), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n585), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n459), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

