//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G116), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(KEYINPUT65), .A3(G119), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(new_n189), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT2), .B(G113), .Z(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n200), .A2(new_n202), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G101), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n198), .A2(new_n201), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n198), .A2(new_n201), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n217), .A2(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n216), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n216), .B(new_n227), .C1(new_n222), .C2(new_n225), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(KEYINPUT6), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n232), .B2(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(G146), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G143), .ZN(new_n236));
  OAI211_X1 g050(.A(G128), .B(new_n233), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G125), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(G146), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n239), .B(new_n240), .C1(KEYINPUT1), .C2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT0), .A4(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n234), .A2(new_n236), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n247), .B2(new_n238), .ZN(new_n248));
  INV_X1    g062(.A(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G224), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n226), .A2(new_n252), .A3(new_n228), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n231), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n248), .A2(new_n255), .A3(KEYINPUT7), .A4(new_n250), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n230), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n220), .B1(new_n199), .B2(new_n193), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n193), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n215), .A2(new_n202), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n258), .A2(new_n215), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n227), .B(KEYINPUT8), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n250), .A2(KEYINPUT7), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n255), .B1(new_n248), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n250), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n262), .A2(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(G902), .B1(new_n257), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G210), .B1(G237), .B2(G902), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT80), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n254), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n254), .B2(new_n268), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n187), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT11), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(G137), .ZN(new_n279));
  INV_X1    g093(.A(G137), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT11), .A3(G134), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(G137), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n279), .A2(new_n281), .A3(new_n285), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n237), .A2(new_n242), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n237), .A2(KEYINPUT67), .A3(new_n242), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(KEYINPUT10), .A3(new_n295), .A4(new_n215), .ZN(new_n296));
  INV_X1    g110(.A(new_n247), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n219), .C1(new_n223), .C2(new_n224), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n237), .A2(new_n210), .A3(new_n213), .A4(new_n242), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n291), .A2(new_n296), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G110), .B(G140), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n249), .A2(G227), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT77), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n296), .A2(new_n298), .A3(new_n301), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n284), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT66), .B1(new_n284), .B2(new_n286), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n309), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n292), .A2(new_n214), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n299), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT12), .A3(new_n287), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  AOI211_X1 g135(.A(new_n321), .B(KEYINPUT12), .C1(new_n315), .C2(new_n319), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n290), .A3(new_n289), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT76), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n320), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(new_n302), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n305), .B(KEYINPUT75), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n317), .B(G469), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(G469), .A2(G902), .ZN(new_n330));
  INV_X1    g144(.A(G469), .ZN(new_n331));
  INV_X1    g145(.A(G902), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n323), .A2(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n321), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(KEYINPUT76), .A3(new_n324), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n307), .B1(new_n336), .B2(new_n320), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n306), .B1(new_n316), .B2(new_n302), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n331), .B(new_n332), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n330), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G221), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT9), .B(G234), .Z(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(new_n332), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT81), .B(new_n187), .C1(new_n272), .C2(new_n273), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n276), .A2(new_n340), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G475), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT16), .ZN(new_n350));
  INV_X1    g164(.A(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G125), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n352), .A2(KEYINPUT16), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(G146), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G146), .B1(new_n350), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n348), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n350), .A2(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n235), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT85), .A3(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n232), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n285), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n365), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G131), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n366), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n361), .B(new_n367), .C1(KEYINPUT17), .C2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(KEYINPUT18), .A3(G131), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT18), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n364), .B(new_n365), .C1(new_n374), .C2(new_n285), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n238), .A2(G140), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n352), .A2(new_n377), .A3(KEYINPUT72), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT72), .B1(new_n352), .B2(new_n377), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n378), .A2(new_n379), .A3(G146), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n349), .A2(new_n235), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT82), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT72), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n238), .A2(G140), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n351), .A2(G125), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n352), .A2(new_n377), .A3(KEYINPUT72), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n235), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n388), .B(new_n389), .C1(new_n235), .C2(new_n349), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n376), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n372), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n203), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n372), .A2(new_n392), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n347), .B1(new_n399), .B2(new_n332), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT19), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n386), .A2(new_n401), .A3(new_n387), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT19), .B1(new_n384), .B2(new_n385), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n235), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n354), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n370), .B1(new_n405), .B2(KEYINPUT83), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n407), .A3(new_n354), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n391), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT84), .B1(new_n409), .B2(new_n395), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n404), .A2(new_n407), .A3(new_n354), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n407), .B1(new_n404), .B2(new_n354), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n412), .A2(new_n413), .A3(new_n370), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n411), .B(new_n396), .C1(new_n414), .C2(new_n391), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n415), .A3(new_n398), .ZN(new_n416));
  NOR2_X1   g230(.A1(G475), .A2(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT20), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n420), .A3(new_n417), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n400), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n232), .A2(G128), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n241), .A2(G143), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n424), .A2(new_n425), .A3(new_n278), .ZN(new_n426));
  INV_X1    g240(.A(G122), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G116), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n191), .A2(G122), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G107), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n206), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT13), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n424), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n425), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n424), .A2(new_n434), .ZN(new_n437));
  OAI21_X1  g251(.A(G134), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n440));
  OAI211_X1 g254(.A(G107), .B(new_n440), .C1(new_n430), .C2(KEYINPUT14), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n278), .B1(new_n424), .B2(new_n425), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n441), .B(new_n432), .C1(new_n426), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT70), .B(G217), .Z(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n342), .A3(new_n249), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n446), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n452), .A3(new_n446), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n332), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n454), .A2(new_n456), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n423), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT88), .A3(new_n457), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(G234), .A2(G237), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n465), .A2(G902), .A3(G953), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n249), .A2(G952), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n465), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT89), .Z(new_n472));
  NAND3_X1  g286(.A1(new_n422), .A2(new_n464), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n346), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n289), .A2(new_n297), .A3(new_n290), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n280), .A2(KEYINPUT64), .A3(G134), .ZN(new_n477));
  INV_X1    g291(.A(new_n282), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT64), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n278), .B2(G137), .ZN(new_n480));
  OAI211_X1 g294(.A(G131), .B(new_n477), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n294), .A2(new_n286), .A3(new_n481), .A4(new_n295), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n220), .A2(new_n221), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n284), .A2(new_n286), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n286), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n486), .A2(new_n247), .B1(new_n487), .B2(new_n292), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n362), .A2(G210), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT27), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G101), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n476), .A2(new_n484), .A3(new_n482), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT31), .ZN(new_n498));
  INV_X1    g312(.A(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n488), .A2(new_n485), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n496), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT31), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n491), .A2(new_n506), .A3(new_n495), .A4(new_n496), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n498), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  NOR2_X1   g323(.A1(G472), .A2(G902), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G472), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n515));
  INV_X1    g329(.A(new_n496), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n484), .B1(new_n476), .B2(new_n482), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n515), .B(KEYINPUT28), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n500), .B1(new_n519), .B2(new_n496), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n501), .A2(KEYINPUT68), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n499), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n502), .A2(new_n504), .A3(new_n499), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n491), .A2(new_n496), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n499), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n514), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n475), .B1(new_n513), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n508), .A2(new_n510), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT32), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n525), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G472), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(KEYINPUT69), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT22), .B(G137), .ZN(new_n540));
  INV_X1    g354(.A(G234), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n341), .A2(new_n541), .A3(G953), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n540), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT23), .B1(new_n241), .B2(G119), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT71), .B1(new_n241), .B2(G119), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT24), .B(G110), .Z(new_n549));
  OAI22_X1  g363(.A1(new_n547), .A2(G110), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n354), .A3(new_n388), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(G110), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n548), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n552), .B(new_n553), .C1(new_n355), .C2(new_n356), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n551), .A2(KEYINPUT73), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT73), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n544), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n543), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n539), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n559), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n567), .B2(new_n544), .ZN(new_n568));
  OAI211_X1 g382(.A(KEYINPUT74), .B(KEYINPUT25), .C1(new_n568), .C2(G902), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n445), .B1(new_n541), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n562), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n568), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n474), .A2(new_n531), .A3(new_n538), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  AOI21_X1  g393(.A(new_n514), .B1(new_n508), .B2(new_n332), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n532), .B1(new_n581), .B2(KEYINPUT90), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n340), .A2(new_n344), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(new_n576), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n399), .A2(new_n332), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G475), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n416), .A2(new_n420), .A3(new_n417), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n420), .B1(new_n416), .B2(new_n417), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n450), .A2(new_n453), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n332), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT91), .B(G478), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n447), .A2(KEYINPUT33), .A3(new_n449), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n455), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n472), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n605), .A2(new_n606), .A3(new_n274), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n588), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G104), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  AOI21_X1  g425(.A(new_n400), .B1(new_n592), .B2(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n419), .A2(new_n421), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(KEYINPUT93), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n464), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n472), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n614), .A2(new_n464), .A3(new_n606), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n274), .B1(new_n619), .B2(KEYINPUT94), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n620), .A3(new_n588), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NOR2_X1   g437(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n567), .B(new_n624), .Z(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n574), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n572), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n474), .A2(new_n585), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  INV_X1    g444(.A(new_n470), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n466), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n614), .A2(new_n464), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n187), .ZN(new_n636));
  INV_X1    g450(.A(new_n273), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n254), .A2(new_n268), .A3(new_n271), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n340), .A2(new_n639), .A3(new_n344), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n531), .A2(new_n538), .A3(new_n627), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n241), .ZN(G30));
  XOR2_X1   g457(.A(new_n633), .B(KEYINPUT39), .Z(new_n644));
  NAND3_X1  g458(.A1(new_n340), .A2(new_n344), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT40), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n646), .A2(KEYINPUT97), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(KEYINPUT97), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n499), .B1(new_n516), .B2(new_n517), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n497), .A2(new_n649), .A3(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n332), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT95), .B1(new_n497), .B2(new_n649), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n511), .B2(new_n512), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n535), .A2(KEYINPUT96), .A3(new_n653), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n627), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n637), .A2(new_n638), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT38), .Z(new_n660));
  NOR4_X1   g474(.A1(new_n660), .A2(new_n422), .A3(new_n464), .A4(new_n636), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n647), .A2(new_n648), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  AND4_X1   g477(.A1(new_n531), .A2(new_n538), .A3(new_n627), .A4(new_n640), .ZN(new_n664));
  INV_X1    g478(.A(new_n604), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n613), .B2(new_n590), .ZN(new_n666));
  INV_X1    g480(.A(new_n633), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT98), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n593), .A2(KEYINPUT98), .A3(new_n604), .A4(new_n667), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AOI21_X1  g487(.A(new_n338), .B1(new_n326), .B2(new_n308), .ZN(new_n674));
  OAI21_X1  g488(.A(G469), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n339), .A3(new_n344), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT99), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n339), .A3(new_n678), .A4(new_n344), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n531), .A2(new_n680), .A3(new_n538), .A4(new_n577), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n607), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND3_X1  g498(.A1(new_n618), .A2(new_n620), .A3(new_n681), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  AND2_X1   g500(.A1(new_n531), .A2(new_n538), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n677), .A2(new_n639), .A3(new_n679), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n473), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n687), .A2(KEYINPUT100), .A3(new_n627), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n531), .A2(new_n538), .A3(new_n627), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n593), .A2(new_n463), .A3(new_n606), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n639), .A3(new_n679), .A4(new_n677), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND2_X1  g511(.A1(new_n508), .A2(new_n332), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT101), .B(G472), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n498), .B(new_n507), .C1(new_n522), .C2(new_n495), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n510), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n577), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n677), .A2(new_n472), .A3(new_n639), .A4(new_n679), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n422), .B2(new_n464), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n593), .A2(KEYINPUT102), .A3(new_n463), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n668), .B2(new_n670), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n593), .A2(new_n604), .A3(new_n667), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n669), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n703), .A2(new_n627), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n688), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n713), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  AND3_X1   g536(.A1(new_n531), .A2(new_n538), .A3(new_n577), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n586), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n340), .A2(KEYINPUT104), .A3(new_n344), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n659), .A2(new_n636), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n713), .A2(new_n723), .A3(new_n718), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n716), .A2(new_n717), .A3(new_n669), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n717), .B1(new_n716), .B2(new_n669), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n726), .A4(new_n727), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n576), .B1(new_n535), .B2(new_n537), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n729), .A2(new_n730), .B1(new_n733), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n285), .ZN(G33));
  NAND3_X1  g555(.A1(new_n723), .A2(new_n634), .A3(new_n728), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND2_X1  g557(.A1(new_n422), .A2(new_n604), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n585), .B1(new_n572), .B2(new_n626), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT44), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT108), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n317), .B1(new_n327), .B2(new_n328), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n331), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n330), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(KEYINPUT106), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n339), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n343), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT44), .B1(new_n749), .B2(new_n750), .ZN(new_n764));
  INV_X1    g578(.A(new_n727), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n752), .A2(new_n644), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  INV_X1    g582(.A(new_n762), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n344), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n774));
  OAI22_X1  g588(.A1(new_n762), .A2(new_n343), .B1(new_n774), .B2(new_n771), .ZN(new_n775));
  INV_X1    g589(.A(new_n671), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n776), .A2(new_n687), .A3(new_n577), .A4(new_n765), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  NAND2_X1  g593(.A1(new_n664), .A2(new_n634), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n340), .A2(new_n344), .A3(new_n667), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n658), .A2(new_n710), .A3(new_n639), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n721), .A2(new_n780), .A3(new_n672), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n639), .A2(new_n782), .A3(new_n708), .A4(new_n709), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n664), .A2(new_n671), .B1(new_n787), .B2(new_n658), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(KEYINPUT52), .A3(new_n780), .A4(new_n721), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n681), .A2(new_n607), .B1(new_n710), .B2(new_n706), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n696), .A2(new_n791), .A3(new_n685), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n461), .A2(new_n457), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n727), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n614), .A3(new_n781), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n687), .A2(new_n627), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n742), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n627), .A2(new_n702), .A3(new_n700), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n731), .A2(new_n732), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n605), .B1(new_n593), .B2(new_n794), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n276), .A2(new_n472), .A3(new_n345), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n585), .A2(new_n802), .A3(new_n587), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n578), .A2(new_n628), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n798), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n729), .A2(new_n730), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n733), .A2(new_n739), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n792), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n790), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n680), .A2(new_n799), .A3(new_n639), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n731), .A2(new_n732), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT110), .B1(new_n813), .B2(new_n642), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n721), .A2(new_n815), .A3(new_n780), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n672), .A2(new_n783), .A3(KEYINPUT52), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n786), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n811), .A2(KEYINPUT53), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n792), .A2(new_n824), .A3(new_n809), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n696), .A2(new_n791), .A3(new_n685), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT111), .B1(new_n740), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n819), .A2(new_n823), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n790), .B2(new_n810), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT112), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n830), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(KEYINPUT54), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n822), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n680), .A2(new_n727), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n749), .A2(new_n631), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n656), .A2(new_n657), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n577), .A3(new_n839), .A4(new_n631), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n422), .A2(new_n665), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n838), .A2(new_n719), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n704), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n749), .A2(new_n631), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n660), .A2(new_n680), .A3(new_n636), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT113), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n842), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n675), .A2(new_n339), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n344), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n773), .B2(new_n775), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n844), .A2(new_n765), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n852), .B(KEYINPUT51), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n737), .A2(new_n738), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n838), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT48), .ZN(new_n863));
  OAI221_X1 g677(.A(new_n469), .B1(new_n605), .B2(new_n840), .C1(new_n844), .C2(new_n688), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n858), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n855), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n852), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n860), .B(new_n865), .C1(new_n868), .C2(KEYINPUT51), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n836), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n660), .A2(new_n577), .A3(new_n344), .A4(new_n187), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n853), .B(KEYINPUT49), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n744), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n839), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(G75));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n249), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n332), .B1(new_n828), .B2(new_n830), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(new_n270), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n231), .A2(new_n253), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n251), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n878), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n883), .B(KEYINPUT116), .Z(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(KEYINPUT56), .B(new_n887), .C1(new_n879), .C2(new_n270), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n876), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n834), .A2(G902), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n271), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n883), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n880), .A2(new_n886), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(KEYINPUT117), .A3(new_n894), .A4(new_n878), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n895), .ZN(G51));
  XNOR2_X1  g710(.A(new_n674), .B(KEYINPUT118), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n834), .B(new_n831), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n330), .B(KEYINPUT57), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n891), .A2(new_n756), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n877), .B1(new_n900), .B2(new_n901), .ZN(G54));
  AND2_X1   g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n879), .A2(new_n416), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n416), .B1(new_n879), .B2(new_n903), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n878), .B(new_n904), .C1(new_n905), .C2(KEYINPUT119), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n834), .A2(G902), .A3(new_n903), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n416), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT120), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n907), .B2(new_n416), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n877), .B1(new_n907), .B2(new_n416), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n905), .A2(KEYINPUT119), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n915), .ZN(G60));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT59), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n599), .A2(new_n600), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n878), .B1(new_n898), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n836), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n601), .ZN(G63));
  NAND2_X1  g736(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n923));
  OR2_X1    g737(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n828), .B2(new_n830), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n625), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n878), .B1(new_n927), .B2(new_n573), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n923), .B(new_n924), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(G66));
  INV_X1    g747(.A(G224), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n467), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n826), .A2(new_n805), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n881), .B1(G898), .B2(new_n249), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n937), .B(new_n939), .ZN(G69));
  INV_X1    g754(.A(new_n752), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n766), .A2(new_n763), .A3(new_n644), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n814), .A2(new_n816), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n672), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n710), .A2(new_n639), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n861), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n763), .A2(new_n947), .A3(new_n644), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n778), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n943), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n809), .A2(new_n742), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT124), .Z(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n249), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n483), .A2(new_n490), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n402), .A2(new_n403), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(G900), .B2(G953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n249), .B1(G227), .B2(G900), .ZN(new_n959));
  AOI22_X1  g773(.A1(new_n953), .A2(new_n958), .B1(KEYINPUT125), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n944), .A2(new_n662), .A3(new_n672), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n765), .A2(new_n645), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n723), .A2(new_n802), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n767), .A2(new_n778), .A3(new_n965), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n957), .B1(new_n967), .B2(G953), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n960), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n960), .B2(new_n968), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(new_n527), .A2(new_n495), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n967), .A2(new_n936), .ZN(new_n974));
  XOR2_X1   g788(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n975));
  NOR2_X1   g789(.A1(new_n514), .A2(new_n332), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  AOI21_X1  g792(.A(new_n973), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n950), .A2(new_n936), .A3(new_n952), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n495), .B(new_n527), .C1(new_n980), .C2(new_n978), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n528), .A2(new_n497), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n821), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n878), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n979), .A2(new_n981), .A3(new_n984), .ZN(G57));
endmodule


