

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595;

  NOR2_X2 U321 ( .A1(n424), .A2(n532), .ZN(n577) );
  XNOR2_X1 U322 ( .A(n390), .B(n290), .ZN(n391) );
  XNOR2_X1 U323 ( .A(G106GAT), .B(G78GAT), .ZN(n348) );
  NOR2_X1 U324 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U325 ( .A(n365), .B(n364), .ZN(n489) );
  XNOR2_X1 U326 ( .A(n486), .B(KEYINPUT104), .ZN(n487) );
  XNOR2_X1 U327 ( .A(n392), .B(n391), .ZN(n399) );
  XOR2_X1 U328 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n289) );
  XOR2_X1 U329 ( .A(n389), .B(n388), .Z(n290) );
  INV_X1 U330 ( .A(KEYINPUT45), .ZN(n346) );
  XNOR2_X1 U331 ( .A(n347), .B(n346), .ZN(n366) );
  INV_X1 U332 ( .A(KEYINPUT47), .ZN(n375) );
  XNOR2_X1 U333 ( .A(n448), .B(n447), .ZN(n449) );
  OR2_X1 U334 ( .A1(n356), .A2(n355), .ZN(n357) );
  INV_X1 U335 ( .A(KEYINPUT37), .ZN(n486) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U337 ( .A1(n536), .A2(n474), .ZN(n475) );
  INV_X1 U338 ( .A(KEYINPUT48), .ZN(n380) );
  NOR2_X1 U339 ( .A1(n460), .A2(n473), .ZN(n461) );
  NOR2_X1 U340 ( .A1(n552), .A2(n539), .ZN(n542) );
  XNOR2_X1 U341 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U342 ( .A(KEYINPUT119), .B(n461), .ZN(n462) );
  XNOR2_X1 U343 ( .A(n459), .B(n458), .ZN(n473) );
  XNOR2_X1 U344 ( .A(n489), .B(n369), .ZN(n571) );
  XNOR2_X1 U345 ( .A(KEYINPUT38), .B(n493), .ZN(n516) );
  XNOR2_X1 U346 ( .A(n463), .B(G190GAT), .ZN(n464) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U348 ( .A(n497), .B(n496), .ZN(G1348GAT) );
  XOR2_X1 U349 ( .A(G29GAT), .B(G43GAT), .Z(n292) );
  XNOR2_X1 U350 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U351 ( .A(n292), .B(n291), .ZN(n310) );
  XOR2_X1 U352 ( .A(G141GAT), .B(G22GAT), .Z(n433) );
  XNOR2_X1 U353 ( .A(n310), .B(n433), .ZN(n293) );
  XOR2_X1 U354 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XNOR2_X1 U355 ( .A(n293), .B(n385), .ZN(n296) );
  XOR2_X1 U356 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n295) );
  NAND2_X1 U357 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U358 ( .A(n295), .B(n294), .Z(n297) );
  NAND2_X1 U359 ( .A1(n296), .A2(n297), .ZN(n301) );
  INV_X1 U360 ( .A(n296), .ZN(n299) );
  INV_X1 U361 ( .A(n297), .ZN(n298) );
  NAND2_X1 U362 ( .A1(n299), .A2(n298), .ZN(n300) );
  NAND2_X1 U363 ( .A1(n301), .A2(n300), .ZN(n306) );
  XOR2_X1 U364 ( .A(KEYINPUT68), .B(G197GAT), .Z(n303) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U367 ( .A(n304), .B(KEYINPUT66), .Z(n305) );
  XNOR2_X1 U368 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U369 ( .A(KEYINPUT67), .B(G1GAT), .Z(n341) );
  XNOR2_X1 U370 ( .A(n307), .B(n341), .ZN(n309) );
  XNOR2_X1 U371 ( .A(G50GAT), .B(G36GAT), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n309), .B(n308), .ZN(n490) );
  XOR2_X1 U373 ( .A(G92GAT), .B(n310), .Z(n312) );
  NAND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n317) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .Z(n386) );
  XNOR2_X1 U378 ( .A(n427), .B(n386), .ZN(n315) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n313), .B(KEYINPUT70), .ZN(n349) );
  INV_X1 U381 ( .A(n349), .ZN(n314) );
  XNOR2_X1 U382 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U383 ( .A(n317), .B(n316), .ZN(n325) );
  XOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n319) );
  XNOR2_X1 U385 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n318) );
  XNOR2_X1 U386 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U387 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n321) );
  XNOR2_X1 U388 ( .A(G134GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U389 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U390 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U391 ( .A(n325), .B(n324), .ZN(n565) );
  XOR2_X1 U392 ( .A(KEYINPUT36), .B(n565), .Z(n592) );
  XOR2_X1 U393 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n327) );
  XNOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT80), .ZN(n326) );
  XNOR2_X1 U395 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U396 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n329) );
  XNOR2_X1 U397 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n328) );
  XNOR2_X1 U398 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U399 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U400 ( .A(G155GAT), .B(G78GAT), .Z(n333) );
  XNOR2_X1 U401 ( .A(G183GAT), .B(G71GAT), .ZN(n332) );
  XNOR2_X1 U402 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U403 ( .A(G64GAT), .B(G211GAT), .Z(n335) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G8GAT), .ZN(n334) );
  XNOR2_X1 U405 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U406 ( .A(n337), .B(n336), .Z(n343) );
  XOR2_X1 U407 ( .A(KEYINPUT13), .B(G57GAT), .Z(n355) );
  XOR2_X1 U408 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XOR2_X1 U409 ( .A(n355), .B(n442), .Z(n339) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U411 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U412 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U413 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n345), .B(n344), .ZN(n588) );
  NOR2_X1 U415 ( .A1(n592), .A2(n588), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n348), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U417 ( .A(n429), .B(n349), .ZN(n354) );
  NAND2_X1 U418 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n289), .B(n350), .ZN(n352) );
  INV_X1 U420 ( .A(KEYINPUT69), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n356) );
  NAND2_X1 U423 ( .A1(n356), .A2(n355), .ZN(n358) );
  NAND2_X1 U424 ( .A1(n358), .A2(n357), .ZN(n361) );
  XOR2_X1 U425 ( .A(G120GAT), .B(G71GAT), .Z(n443) );
  XNOR2_X1 U426 ( .A(G176GAT), .B(G92GAT), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n359), .B(G64GAT), .ZN(n387) );
  XOR2_X1 U428 ( .A(n443), .B(n387), .Z(n360) );
  XNOR2_X1 U429 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U430 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n363) );
  XNOR2_X1 U431 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  NOR2_X1 U433 ( .A1(n366), .A2(n489), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n367), .B(KEYINPUT113), .ZN(n368) );
  NOR2_X1 U435 ( .A1(n490), .A2(n368), .ZN(n379) );
  INV_X1 U436 ( .A(KEYINPUT41), .ZN(n369) );
  NAND2_X1 U437 ( .A1(n490), .A2(n571), .ZN(n371) );
  XNOR2_X1 U438 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n372) );
  AND2_X1 U440 ( .A1(n372), .A2(n588), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n373), .B(KEYINPUT111), .ZN(n374) );
  NOR2_X1 U442 ( .A1(n374), .A2(n565), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U444 ( .A(KEYINPUT112), .B(n377), .ZN(n378) );
  NOR2_X1 U445 ( .A1(n379), .A2(n378), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n554) );
  XOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U448 ( .A(KEYINPUT83), .B(G183GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U450 ( .A(KEYINPUT19), .B(n384), .ZN(n457) );
  XOR2_X1 U451 ( .A(n385), .B(n457), .Z(n392) );
  XOR2_X1 U452 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U453 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n389) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XOR2_X1 U455 ( .A(KEYINPUT21), .B(G204GAT), .Z(n394) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(G211GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U458 ( .A(G218GAT), .B(KEYINPUT87), .Z(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n438) );
  INV_X1 U460 ( .A(n438), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n397), .B(KEYINPUT91), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n534) );
  NAND2_X1 U463 ( .A1(n554), .A2(n534), .ZN(n401) );
  XOR2_X1 U464 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n424) );
  XOR2_X1 U466 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n403) );
  XNOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n402) );
  XOR2_X1 U468 ( .A(n403), .B(n402), .Z(n422) );
  XOR2_X1 U469 ( .A(G162GAT), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U470 ( .A(G120GAT), .B(G127GAT), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U472 ( .A(KEYINPUT90), .B(G57GAT), .Z(n407) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G141GAT), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U475 ( .A(n409), .B(n408), .Z(n415) );
  XNOR2_X1 U476 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n410), .B(KEYINPUT2), .ZN(n428) );
  XOR2_X1 U478 ( .A(G85GAT), .B(n428), .Z(n412) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n413), .B(G29GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U483 ( .A(n416), .B(KEYINPUT6), .Z(n420) );
  XOR2_X1 U484 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n418) );
  XNOR2_X1 U485 ( .A(G113GAT), .B(G134GAT), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n450) );
  XNOR2_X1 U487 ( .A(n450), .B(KEYINPUT88), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n466) );
  INV_X1 U490 ( .A(n466), .ZN(n423) );
  INV_X1 U491 ( .A(n423), .ZN(n532) );
  XOR2_X1 U492 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n437) );
  XOR2_X1 U495 ( .A(n428), .B(n427), .Z(n435) );
  XOR2_X1 U496 ( .A(n429), .B(KEYINPUT23), .Z(n431) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n474) );
  NAND2_X1 U503 ( .A1(n577), .A2(n474), .ZN(n441) );
  XOR2_X1 U504 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n460) );
  XOR2_X1 U506 ( .A(KEYINPUT20), .B(G190GAT), .Z(n445) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U509 ( .A(n446), .B(G99GAT), .Z(n453) );
  NAND2_X1 U510 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  INV_X1 U511 ( .A(G169GAT), .ZN(n447) );
  XNOR2_X1 U512 ( .A(G43GAT), .B(n451), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n455) );
  XNOR2_X1 U515 ( .A(G176GAT), .B(KEYINPUT64), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U517 ( .A(n473), .ZN(n536) );
  INV_X1 U518 ( .A(n462), .ZN(n574) );
  NAND2_X1 U519 ( .A1(n574), .A2(n565), .ZN(n465) );
  XOR2_X1 U520 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n463) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  INV_X1 U522 ( .A(n588), .ZN(n575) );
  XNOR2_X1 U523 ( .A(n534), .B(KEYINPUT27), .ZN(n476) );
  NAND2_X1 U524 ( .A1(n466), .A2(n476), .ZN(n552) );
  XNOR2_X1 U525 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(n474), .ZN(n539) );
  XNOR2_X1 U527 ( .A(KEYINPUT94), .B(n542), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n468), .A2(n473), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT95), .ZN(n482) );
  NAND2_X1 U530 ( .A1(n536), .A2(n534), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT97), .B(n470), .Z(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n474), .ZN(n472) );
  XNOR2_X1 U533 ( .A(KEYINPUT25), .B(n472), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT26), .B(n475), .Z(n553) );
  INV_X1 U535 ( .A(n553), .ZN(n578) );
  AND2_X1 U536 ( .A1(n578), .A2(n476), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT96), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n532), .A2(n480), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT98), .ZN(n500) );
  NOR2_X1 U541 ( .A1(n575), .A2(n500), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(KEYINPUT103), .ZN(n485) );
  NOR2_X1 U543 ( .A1(n485), .A2(n592), .ZN(n488) );
  XNOR2_X1 U544 ( .A(n488), .B(n487), .ZN(n529) );
  INV_X1 U545 ( .A(n489), .ZN(n585) );
  INV_X1 U546 ( .A(n490), .ZN(n579) );
  INV_X1 U547 ( .A(n579), .ZN(n557) );
  NAND2_X1 U548 ( .A1(n585), .A2(n557), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(KEYINPUT73), .ZN(n502) );
  NAND2_X1 U550 ( .A1(n529), .A2(n502), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT105), .ZN(n493) );
  NAND2_X1 U552 ( .A1(n516), .A2(n536), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n574), .A2(n557), .ZN(n497) );
  XNOR2_X1 U555 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n496) );
  NOR2_X1 U556 ( .A1(n565), .A2(n588), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT16), .B(n498), .Z(n499) );
  NOR2_X1 U558 ( .A1(n500), .A2(n499), .ZN(n501) );
  XOR2_X1 U559 ( .A(KEYINPUT99), .B(n501), .Z(n519) );
  AND2_X1 U560 ( .A1(n502), .A2(n519), .ZN(n510) );
  NAND2_X1 U561 ( .A1(n510), .A2(n532), .ZN(n506) );
  XOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n504) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(G1324GAT) );
  NAND2_X1 U566 ( .A1(n510), .A2(n534), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT35), .Z(n509) );
  NAND2_X1 U569 ( .A1(n510), .A2(n536), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  NAND2_X1 U571 ( .A1(n539), .A2(n510), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n511), .B(KEYINPUT102), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G22GAT), .B(n512), .ZN(G1327GAT) );
  XOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT39), .Z(n514) );
  NAND2_X1 U575 ( .A1(n532), .A2(n516), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1328GAT) );
  NAND2_X1 U577 ( .A1(n516), .A2(n534), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n539), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n517), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U581 ( .A1(n571), .A2(n579), .ZN(n518) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(n518), .Z(n530) );
  AND2_X1 U583 ( .A1(n519), .A2(n530), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n532), .A2(n526), .ZN(n520) );
  XNOR2_X1 U585 ( .A(KEYINPUT42), .B(n520), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  XOR2_X1 U587 ( .A(G64GAT), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U588 ( .A1(n526), .A2(n534), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1333GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n536), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT108), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G71GAT), .B(n525), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U594 ( .A1(n526), .A2(n539), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT109), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n532), .A2(n538), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n533), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n534), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n536), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(KEYINPUT44), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  NAND2_X1 U607 ( .A1(n554), .A2(n542), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n473), .A2(n543), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n549), .A2(n557), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U612 ( .A1(n549), .A2(n571), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U614 ( .A1(n575), .A2(n549), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U618 ( .A1(n549), .A2(n565), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT114), .B(n556), .Z(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(n561), .Z(n563) );
  NAND2_X1 U629 ( .A1(n566), .A2(n571), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n575), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(n570), .Z(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U643 ( .A1(n577), .A2(n578), .ZN(n591) );
  NOR2_X1 U644 ( .A1(n579), .A2(n591), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT124), .B(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n591), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n591), .ZN(n589) );
  XOR2_X1 U654 ( .A(KEYINPUT126), .B(n589), .Z(n590) );
  XNOR2_X1 U655 ( .A(G211GAT), .B(n590), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U657 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

