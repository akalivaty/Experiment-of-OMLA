//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1046, new_n1047;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT67), .B1(new_n206), .B2(G113gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n204), .B(new_n205), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G127gat), .B(G134gat), .Z(new_n213));
  XNOR2_X1  g012(.A(G113gat), .B(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(KEYINPUT1), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT68), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n212), .A2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n226), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n223), .B(new_n225), .C1(new_n227), .C2(new_n222), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n230), .A2(new_n231), .A3(new_n224), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n221), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  OR3_X1    g032(.A1(new_n230), .A2(new_n231), .A3(new_n224), .ZN(new_n234));
  INV_X1    g033(.A(new_n222), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n235), .A2(new_n237), .B1(new_n230), .B2(new_n224), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n234), .A2(new_n238), .A3(KEYINPUT25), .A4(new_n223), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n222), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(KEYINPUT66), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n243), .A2(new_n236), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n229), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  INV_X1    g049(.A(G183gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(KEYINPUT27), .ZN(new_n252));
  INV_X1    g051(.A(G190gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT27), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n254), .B2(G183gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(KEYINPUT64), .A3(KEYINPUT27), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n249), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT28), .A3(new_n253), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n248), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n217), .B(new_n220), .C1(new_n240), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G227gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n263), .ZN(new_n269));
  INV_X1    g068(.A(new_n248), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n233), .A2(new_n239), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT68), .A4(new_n216), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n265), .A2(KEYINPUT69), .A3(new_n268), .A4(new_n273), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n203), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT33), .B1(new_n276), .B2(new_n277), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G71gat), .ZN(new_n281));
  INV_X1    g080(.A(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n278), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  AOI221_X4 g084(.A(new_n203), .B1(KEYINPUT33), .B2(new_n283), .C1(new_n276), .C2(new_n277), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT70), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n273), .ZN(new_n288));
  INV_X1    g087(.A(new_n268), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n288), .A2(KEYINPUT34), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT34), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n284), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n278), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n278), .B1(new_n279), .B2(new_n284), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n287), .A2(new_n292), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n292), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT36), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n202), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n292), .B1(new_n285), .B2(new_n286), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(new_n303), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT36), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n297), .A2(new_n302), .A3(KEYINPUT72), .A4(new_n299), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n287), .A2(new_n292), .A3(new_n300), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n312), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n303), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G155gat), .B(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(G148gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G141gat), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G148gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n317), .A2(new_n319), .B1(KEYINPUT2), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n318), .A2(G148gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n316), .A2(G141gat), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT79), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331));
  OAI211_X1 g130(.A(KEYINPUT78), .B(new_n315), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n216), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n212), .A2(new_n215), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n322), .B1(new_n321), .B2(KEYINPUT79), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n322), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n339));
  XOR2_X1   g138(.A(G155gat), .B(G162gat), .Z(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n332), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n333), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT5), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n342), .B2(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n329), .A2(KEYINPUT3), .A3(new_n332), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n337), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n332), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n218), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n352), .A2(new_n356), .A3(new_n346), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n333), .B(new_n355), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(KEYINPUT5), .A3(new_n346), .A4(new_n352), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n359), .A2(new_n364), .A3(new_n366), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n364), .B1(new_n359), .B2(new_n366), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT6), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(KEYINPUT87), .ZN(new_n374));
  OR3_X1    g173(.A1(new_n367), .A2(KEYINPUT87), .A3(new_n368), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT37), .ZN(new_n376));
  NAND2_X1  g175(.A1(G211gat), .A2(G218gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G197gat), .B(G204gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(G211gat), .A2(G218gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT75), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G211gat), .ZN(new_n389));
  INV_X1    g188(.A(G218gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n377), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n394), .B2(KEYINPUT74), .ZN(new_n395));
  AND2_X1   g194(.A1(G197gat), .A2(G204gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(G197gat), .A2(G204gat), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n381), .A2(new_n382), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n388), .A2(new_n393), .A3(KEYINPUT74), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n271), .A2(new_n272), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(new_n405), .A3(G226gat), .A4(G233gat), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n269), .A2(new_n270), .B1(new_n233), .B2(new_n239), .ZN(new_n407));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT76), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n407), .B2(KEYINPUT29), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n403), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(G226gat), .A3(G233gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n413), .A3(new_n403), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n376), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G92gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT77), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n419), .B(G64gat), .Z(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n406), .A2(new_n409), .B1(new_n422), .B2(new_n408), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n414), .B(KEYINPUT37), .C1(new_n423), .C2(new_n403), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n414), .B1(new_n423), .B2(new_n403), .ZN(new_n426));
  INV_X1    g225(.A(new_n420), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n425), .A2(KEYINPUT38), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n403), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n413), .A2(new_n411), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n429), .B(KEYINPUT37), .C1(new_n403), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT38), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n431), .A3(new_n432), .A4(new_n420), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n374), .A2(new_n375), .A3(new_n428), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n427), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n414), .B(new_n420), .C1(new_n423), .C2(new_n403), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(new_n438), .A3(new_n427), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(G225gat), .A3(G233gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n345), .A2(new_n346), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT39), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(new_n363), .C1(KEYINPUT39), .C2(new_n443), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT40), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(KEYINPUT86), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n448), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n441), .A2(new_n449), .A3(new_n367), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n421), .B1(new_n395), .B2(new_n402), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT84), .B(new_n351), .C1(new_n452), .C2(new_n353), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n394), .A2(KEYINPUT74), .A3(new_n385), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n400), .A2(new_n401), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT29), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n344), .B(new_n454), .C1(new_n457), .C2(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G228gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(new_n267), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n350), .A2(new_n421), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n403), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n403), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n350), .B2(new_n421), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n400), .A2(new_n394), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n400), .A2(new_n394), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n421), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n353), .B1(new_n469), .B2(new_n349), .ZN(new_n470));
  OAI22_X1  g269(.A1(new_n466), .A2(new_n470), .B1(new_n460), .B2(new_n267), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G22gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474));
  XOR2_X1   g273(.A(G78gat), .B(G106gat), .Z(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT31), .ZN(new_n476));
  INV_X1    g275(.A(G50gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G22gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n471), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n473), .A2(new_n474), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n472), .A2(G22gat), .A3(new_n478), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n464), .A2(new_n471), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(new_n480), .C1(KEYINPUT85), .C2(new_n478), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n434), .A2(new_n451), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n359), .A2(new_n366), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT6), .B1(new_n489), .B2(new_n363), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n371), .B1(new_n490), .B2(KEYINPUT82), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n372), .B2(KEYINPUT6), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n369), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n494), .A2(new_n495), .A3(new_n441), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n363), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT82), .A3(new_n368), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n367), .A3(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n370), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT83), .B1(new_n500), .B2(new_n440), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n488), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n314), .A2(new_n487), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n285), .A2(new_n292), .A3(new_n286), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(new_n488), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n506), .A2(new_n507), .A3(new_n312), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n506), .B2(new_n312), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n496), .A2(new_n501), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT87), .B1(new_n490), .B2(new_n367), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n375), .B1(new_n513), .B2(new_n369), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n514), .A2(new_n504), .A3(new_n486), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n441), .B1(new_n308), .B2(new_n310), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n503), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G57gat), .B(G64gat), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT9), .ZN(new_n523));
  INV_X1    g322(.A(G71gat), .ZN(new_n524));
  INV_X1    g323(.A(G78gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G71gat), .B(G78gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n522), .A2(new_n528), .A3(new_n526), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n530), .A2(KEYINPUT94), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT94), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(G1gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(G1gat), .B2(new_n540), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n251), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n251), .B1(new_n539), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT95), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n546), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n549), .A2(new_n552), .A3(G231gat), .A4(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n549), .A2(new_n552), .B1(G231gat), .B2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n389), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n552), .ZN(new_n560));
  INV_X1    g359(.A(G231gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(new_n267), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n562), .B2(new_n553), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n538), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n557), .B1(new_n554), .B2(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n553), .A3(new_n559), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n537), .ZN(new_n567));
  INV_X1    g366(.A(G232gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(new_n267), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  INV_X1    g373(.A(G29gat), .ZN(new_n575));
  INV_X1    g374(.A(G36gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n577), .A2(new_n578), .B1(G29gat), .B2(G36gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT15), .ZN(new_n580));
  XOR2_X1   g379(.A(G43gat), .B(G50gat), .Z(new_n581));
  OR3_X1    g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n580), .ZN(new_n583));
  XNOR2_X1  g382(.A(G43gat), .B(G50gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n585), .A3(new_n579), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT91), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n582), .A2(KEYINPUT91), .A3(new_n586), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n586), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT17), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n597), .B2(new_n598), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n595), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n569), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT96), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n592), .A2(new_n611), .A3(new_n593), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n587), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n605), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n610), .B1(new_n607), .B2(new_n615), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n573), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n607), .A2(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n609), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n572), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n564), .A2(new_n567), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G113gat), .B(G141gat), .Z(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n545), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n591), .B2(new_n594), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n613), .A2(new_n545), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT92), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n639));
  INV_X1    g438(.A(new_n637), .ZN(new_n640));
  NOR4_X1   g439(.A1(new_n634), .A2(new_n635), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n638), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(new_n645));
  INV_X1    g444(.A(new_n635), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n613), .A2(new_n545), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n637), .B(KEYINPUT13), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n645), .A2(KEYINPUT18), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n632), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n595), .A2(new_n545), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n646), .A3(new_n637), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n639), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n645), .A2(KEYINPUT92), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n642), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n651), .A3(new_n631), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  INV_X1    g460(.A(G176gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n530), .A2(new_n531), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n605), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n604), .A2(new_n667), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n532), .A2(new_n533), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(new_n606), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n606), .B(new_n672), .C1(new_n532), .C2(new_n533), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT97), .B1(new_n534), .B2(new_n605), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n670), .B1(new_n682), .B2(new_n675), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT99), .B1(new_n683), .B2(new_n679), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT10), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n686), .B(new_n671), .C1(new_n674), .C2(new_n676), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n673), .A2(new_n686), .A3(new_n606), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n680), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n665), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT10), .B(new_n670), .C1(new_n682), .C2(new_n675), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n679), .B1(new_n692), .B2(new_n688), .ZN(new_n693));
  INV_X1    g492(.A(new_n665), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n681), .A4(new_n684), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n660), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n625), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n521), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n500), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n440), .ZN(new_n703));
  NAND2_X1  g502(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n541), .A2(new_n544), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n707), .B(new_n708), .C1(new_n544), .C2(new_n703), .ZN(G1325gat));
  INV_X1    g508(.A(G15gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n308), .A2(new_n310), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n700), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT100), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n700), .A2(new_n710), .A3(new_n314), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n486), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  NAND4_X1  g518(.A1(new_n303), .A2(new_n483), .A3(new_n482), .A4(new_n485), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT89), .B1(new_n301), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n495), .B1(new_n494), .B2(new_n441), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n500), .A2(KEYINPUT83), .A3(new_n440), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n506), .A2(new_n507), .A3(new_n312), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT35), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n488), .B1(new_n374), .B2(new_n375), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n727), .A3(new_n504), .A4(new_n440), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT88), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n486), .B1(new_n722), .B2(new_n723), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n434), .A2(new_n486), .A3(new_n451), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n726), .A2(new_n731), .B1(new_n314), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n564), .A2(new_n567), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n698), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n735), .A2(new_n624), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n575), .A3(new_n494), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n731), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n503), .A2(KEYINPUT102), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n734), .A2(new_n746), .A3(new_n314), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n623), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n619), .A2(new_n622), .A3(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT44), .B1(new_n735), .B2(new_n624), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n738), .ZN(new_n758));
  OAI21_X1  g557(.A(G29gat), .B1(new_n758), .B2(new_n500), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n759), .ZN(G1328gat));
  NAND3_X1  g559(.A1(new_n740), .A2(new_n576), .A3(new_n441), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT46), .Z(new_n762));
  OAI21_X1  g561(.A(G36gat), .B1(new_n758), .B2(new_n440), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1329gat));
  INV_X1    g563(.A(new_n314), .ZN(new_n765));
  INV_X1    g564(.A(new_n754), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n746), .A2(new_n314), .A3(new_n487), .A4(new_n502), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n746), .B1(new_n734), .B2(new_n314), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(new_n744), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n521), .B2(new_n623), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n765), .B(new_n738), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n521), .A2(new_n711), .A3(new_n623), .A4(new_n738), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(G43gat), .ZN(new_n776));
  INV_X1    g575(.A(G43gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n740), .A2(KEYINPUT105), .A3(new_n777), .A4(new_n711), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n773), .A2(G43gat), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n779), .A2(KEYINPUT104), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n776), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n314), .B(new_n739), .C1(new_n755), .C2(new_n756), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n777), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT47), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n781), .A2(new_n786), .ZN(G1330gat));
  OAI21_X1  g586(.A(G50gat), .B1(new_n758), .B2(new_n486), .ZN(new_n788));
  NAND2_X1  g587(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n789));
  OR2_X1    g588(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n740), .A2(new_n477), .A3(new_n488), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n739), .B1(new_n755), .B2(new_n756), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n477), .B1(new_n793), .B2(new_n488), .ZN(new_n794));
  INV_X1    g593(.A(new_n791), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT106), .B(KEYINPUT48), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n792), .A2(new_n796), .ZN(G1331gat));
  NOR2_X1   g596(.A1(new_n625), .A2(new_n660), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n748), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n494), .A3(new_n696), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n441), .A3(new_n696), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n803));
  XOR2_X1   g602(.A(KEYINPUT49), .B(G64gat), .Z(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(G1333gat));
  AND3_X1   g604(.A1(new_n799), .A2(new_n711), .A3(new_n696), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n799), .A2(G71gat), .A3(new_n696), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n806), .A2(G71gat), .B1(new_n314), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g608(.A1(new_n799), .A2(new_n488), .A3(new_n696), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g610(.A1(new_n737), .A2(new_n624), .A3(new_n660), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n748), .B2(new_n812), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n696), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n597), .B1(new_n815), .B2(new_n500), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n737), .A2(new_n660), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n757), .A2(new_n696), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n494), .A2(G85gat), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n816), .B(KEYINPUT107), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT107), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n748), .A2(new_n812), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n812), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n697), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(G85gat), .B1(new_n826), .B2(new_n494), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n818), .A2(new_n819), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n821), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n820), .A2(new_n829), .ZN(G1336gat));
  NAND4_X1  g629(.A1(new_n757), .A2(new_n441), .A3(new_n696), .A4(new_n817), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G92gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n697), .A2(G92gat), .A3(new_n440), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT108), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n813), .B2(new_n814), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT109), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(new_n834), .C1(new_n813), .C2(new_n814), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n833), .B1(new_n813), .B2(new_n814), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n832), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(G1337gat));
  AOI21_X1  g643(.A(G99gat), .B1(new_n826), .B2(new_n711), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n818), .A2(new_n282), .A3(new_n314), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(G1338gat));
  XNOR2_X1  g646(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n488), .A2(G106gat), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n488), .B(new_n696), .C1(new_n813), .C2(new_n814), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI221_X1 g650(.A(new_n848), .B1(new_n818), .B2(new_n849), .C1(new_n851), .C2(G106gat), .ZN(new_n852));
  INV_X1    g651(.A(new_n848), .ZN(new_n853));
  AOI21_X1  g652(.A(G106gat), .B1(new_n826), .B2(new_n488), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n818), .A2(new_n849), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(G1339gat));
  NOR3_X1   g656(.A1(new_n625), .A2(new_n696), .A3(new_n660), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n687), .A2(new_n680), .A3(new_n689), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n693), .A2(new_n859), .A3(KEYINPUT54), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n694), .B1(new_n690), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n695), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT55), .B1(new_n860), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n630), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n636), .A2(new_n637), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n648), .A2(new_n650), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n659), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n752), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n696), .A2(new_n659), .A3(new_n870), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n866), .B2(new_n660), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n872), .B1(new_n874), .B2(new_n752), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n858), .B1(new_n875), .B2(new_n736), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT112), .B1(new_n876), .B2(new_n488), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n863), .A2(new_n695), .ZN(new_n878));
  INV_X1    g677(.A(new_n865), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n660), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n873), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n752), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n866), .A2(new_n752), .A3(new_n871), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n736), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n858), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n486), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n877), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(new_n494), .A3(new_n516), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n208), .B1(new_n890), .B2(new_n660), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n500), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n510), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(new_n441), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n893), .A2(KEYINPUT113), .A3(new_n440), .A4(new_n510), .ZN(new_n896));
  INV_X1    g695(.A(new_n660), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(G113gat), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n891), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n891), .B2(new_n899), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1340gat));
  NAND4_X1  g702(.A1(new_n895), .A2(new_n206), .A3(new_n696), .A4(new_n896), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n696), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(G120gat), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT115), .B(new_n206), .C1(new_n890), .C2(new_n696), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G1341gat));
  AND3_X1   g708(.A1(new_n890), .A2(G127gat), .A3(new_n737), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n441), .ZN(new_n911));
  AOI21_X1  g710(.A(G127gat), .B1(new_n911), .B2(new_n737), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n910), .A2(new_n912), .ZN(G1342gat));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n624), .A2(G134gat), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n911), .B2(new_n915), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n890), .ZN(new_n920));
  OAI21_X1  g719(.A(G134gat), .B1(new_n920), .B2(new_n624), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n916), .B2(new_n917), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(G1343gat));
  NOR2_X1   g722(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n860), .A2(new_n862), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n653), .A2(new_n659), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n873), .B1(new_n928), .B2(new_n878), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT118), .B1(new_n929), .B2(new_n623), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n927), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n878), .A2(new_n660), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n881), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n624), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n935), .A3(new_n872), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n858), .B1(new_n936), .B2(new_n736), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n486), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT119), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n876), .B2(new_n486), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n623), .B1(new_n932), .B2(new_n881), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n883), .B1(new_n944), .B2(new_n934), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n737), .B1(new_n945), .B2(new_n930), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n943), .B(new_n939), .C1(new_n946), .C2(new_n858), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n941), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n765), .A2(new_n500), .A3(new_n441), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n660), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G141gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n876), .A2(new_n486), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n952), .A2(new_n318), .A3(new_n660), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n925), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g756(.A(new_n924), .B(new_n955), .C1(new_n950), .C2(G141gat), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(G1344gat));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n948), .A2(new_n949), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n960), .B(G148gat), .C1(new_n961), .C2(new_n697), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n866), .A2(new_n623), .A3(new_n871), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n929), .B2(new_n623), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n858), .B1(new_n964), .B2(new_n736), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n938), .B1(new_n965), .B2(new_n486), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n886), .A2(KEYINPUT57), .A3(new_n488), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n697), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n316), .B1(new_n968), .B2(new_n949), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n962), .B1(new_n969), .B2(new_n960), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n952), .A2(new_n949), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n316), .A3(new_n696), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1345gat));
  INV_X1    g772(.A(G155gat), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n961), .A2(new_n974), .A3(new_n736), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n737), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT121), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n975), .B1(new_n974), .B2(new_n977), .ZN(G1346gat));
  OAI21_X1  g777(.A(G162gat), .B1(new_n961), .B2(new_n753), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n952), .A2(new_n494), .A3(new_n314), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n980), .A2(G162gat), .A3(new_n624), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n441), .B2(new_n981), .ZN(G1347gat));
  INV_X1    g781(.A(G169gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n494), .A2(new_n440), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n889), .A2(new_n711), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n983), .B1(new_n985), .B2(new_n660), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n876), .A2(new_n494), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n508), .A2(new_n509), .A3(new_n440), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n989), .A2(G169gat), .A3(new_n897), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n986), .A2(new_n990), .ZN(G1348gat));
  NAND3_X1  g790(.A1(new_n985), .A2(G176gat), .A3(new_n696), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n662), .B1(new_n989), .B2(new_n697), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n992), .A2(new_n993), .ZN(G1349gat));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n889), .A2(new_n711), .A3(new_n737), .A4(new_n984), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G183gat), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n987), .A2(new_n262), .A3(new_n737), .A4(new_n988), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n995), .B1(new_n999), .B2(KEYINPUT60), .ZN(new_n1000));
  INV_X1    g799(.A(new_n998), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n1001), .B1(new_n996), .B2(G183gat), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT60), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n1002), .A2(KEYINPUT122), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n1005));
  AND4_X1   g804(.A1(new_n1005), .A2(new_n997), .A3(new_n1003), .A4(new_n998), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1005), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1007));
  OAI22_X1  g806(.A1(new_n1000), .A2(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1350gat));
  NAND4_X1  g807(.A1(new_n889), .A2(new_n711), .A3(new_n623), .A4(new_n984), .ZN(new_n1009));
  NAND2_X1  g808(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1009), .A2(G190gat), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g810(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n1012));
  OR2_X1    g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n987), .A2(new_n253), .A3(new_n752), .A4(new_n988), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(G1351gat));
  NOR3_X1   g815(.A1(new_n876), .A2(new_n494), .A3(new_n765), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n486), .A2(new_n440), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g818(.A1(new_n1019), .A2(G197gat), .A3(new_n897), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n314), .A2(new_n984), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1021), .B1(new_n966), .B2(new_n967), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(new_n660), .ZN(new_n1023));
  AOI21_X1  g822(.A(new_n1020), .B1(G197gat), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g823(.A(new_n1024), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g824(.A(new_n1019), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1026), .A2(new_n664), .A3(new_n696), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1028));
  OR3_X1    g827(.A1(new_n1027), .A2(new_n1028), .A3(KEYINPUT62), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1030));
  INV_X1    g829(.A(new_n1021), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n968), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1032), .A2(G204gat), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n1028), .B1(new_n1027), .B2(KEYINPUT62), .ZN(new_n1034));
  NAND4_X1  g833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .A4(new_n1034), .ZN(G1353gat));
  NAND3_X1  g834(.A1(new_n1026), .A2(new_n389), .A3(new_n737), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n966), .A2(new_n967), .ZN(new_n1037));
  NAND3_X1  g836(.A1(new_n1037), .A2(new_n737), .A3(new_n1031), .ZN(new_n1038));
  AND3_X1   g837(.A1(new_n1038), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1039));
  AOI21_X1  g838(.A(KEYINPUT63), .B1(new_n1038), .B2(G211gat), .ZN(new_n1040));
  OAI21_X1  g839(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1041), .A2(KEYINPUT127), .ZN(new_n1042));
  INV_X1    g841(.A(KEYINPUT127), .ZN(new_n1043));
  OAI211_X1 g842(.A(new_n1036), .B(new_n1043), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n1042), .A2(new_n1044), .ZN(G1354gat));
  AOI21_X1  g844(.A(G218gat), .B1(new_n1026), .B2(new_n752), .ZN(new_n1046));
  NOR2_X1   g845(.A1(new_n624), .A2(new_n390), .ZN(new_n1047));
  AOI21_X1  g846(.A(new_n1046), .B1(new_n1022), .B2(new_n1047), .ZN(G1355gat));
endmodule


