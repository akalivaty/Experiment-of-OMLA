//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT2), .A2(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n189), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(new_n195), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n187), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n196), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n195), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(KEYINPUT70), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(KEYINPUT0), .B2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n207), .A2(G146), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT66), .B1(new_n205), .B2(G143), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n207), .A3(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT0), .A3(G128), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n206), .A2(new_n208), .B1(new_n213), .B2(KEYINPUT64), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .A3(new_n210), .A4(new_n212), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n217), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G134), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n233), .A3(G137), .ZN(new_n234));
  NOR2_X1   g048(.A1(G134), .A2(G137), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n229), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT11), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n228), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT67), .B(G134), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n229), .A3(new_n238), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n235), .B1(new_n242), .B2(G137), .ZN(new_n244));
  OAI211_X1 g058(.A(G131), .B(new_n243), .C1(new_n244), .C2(new_n229), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n219), .A2(new_n221), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n249), .A3(new_n206), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n218), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n209), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n230), .A2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n239), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n250), .A2(new_n253), .B1(new_n255), .B2(G131), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n241), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n227), .A2(new_n246), .B1(new_n257), .B2(KEYINPUT68), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n241), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n204), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n227), .A2(new_n246), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n241), .A3(KEYINPUT71), .ZN(new_n265));
  AND4_X1   g079(.A1(new_n204), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT28), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n204), .A2(new_n257), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n270), .B2(new_n262), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n262), .A2(new_n273), .A3(new_n260), .ZN(new_n274));
  INV_X1    g088(.A(new_n204), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n262), .A2(new_n264), .A3(new_n204), .A4(new_n265), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT73), .A3(KEYINPUT28), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n269), .A2(new_n272), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(G101), .ZN(new_n282));
  NOR2_X1   g096(.A1(G237), .A2(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G210), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n282), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n266), .B2(new_n286), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT30), .A4(new_n265), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n226), .B1(new_n241), .B2(new_n245), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n256), .A2(new_n241), .A3(new_n259), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n259), .B1(new_n256), .B2(new_n241), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n275), .B(new_n289), .C1(new_n293), .C2(KEYINPUT30), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n277), .A2(KEYINPUT72), .A3(new_n285), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n288), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n288), .A2(new_n294), .A3(KEYINPUT31), .A4(new_n295), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n280), .A2(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G472), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT74), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(G472), .B2(G902), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT32), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT73), .B1(new_n278), .B2(KEYINPUT28), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n311));
  AOI211_X1 g125(.A(new_n268), .B(new_n311), .C1(new_n276), .C2(new_n277), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n285), .B1(new_n313), .B2(new_n272), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n277), .A2(KEYINPUT72), .A3(new_n285), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT72), .B1(new_n277), .B2(new_n285), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT31), .B1(new_n317), .B2(new_n294), .ZN(new_n318));
  AND4_X1   g132(.A1(KEYINPUT31), .A2(new_n288), .A3(new_n294), .A4(new_n295), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n309), .B(new_n306), .C1(new_n314), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n294), .A2(new_n277), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n286), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n322), .B(new_n324), .C1(new_n280), .C2(new_n286), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n275), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n311), .B1(new_n327), .B2(new_n277), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n328), .A2(new_n322), .A3(new_n271), .ZN(new_n329));
  AOI21_X1  g143(.A(G902), .B1(new_n329), .B2(new_n285), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n308), .A2(new_n321), .B1(G472), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n248), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT24), .B(G110), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT75), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G125), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n342), .B2(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT16), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT16), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(new_n341), .A3(KEYINPUT76), .A4(G125), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n205), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n346), .A3(G146), .A4(new_n348), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G110), .ZN(new_n353));
  OR3_X1    g167(.A1(new_n333), .A2(KEYINPUT23), .A3(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n354), .A2(new_n355), .B1(new_n333), .B2(G128), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n339), .B(new_n352), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n356), .A2(new_n353), .B1(new_n336), .B2(new_n337), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n342), .A2(new_n345), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n351), .B1(G146), .B2(new_n359), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G953), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(G221), .A3(G234), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT22), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n238), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT77), .B1(new_n357), .B2(new_n361), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI211_X1 g183(.A(KEYINPUT77), .B(new_n366), .C1(new_n357), .C2(new_n361), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n302), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT25), .ZN(new_n372));
  INV_X1    g186(.A(G217), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(G234), .B2(new_n302), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n375), .B(new_n302), .C1(new_n369), .C2(new_n370), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n372), .A2(KEYINPUT78), .A3(new_n374), .A4(new_n376), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n369), .A2(new_n370), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n374), .A2(G902), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G469), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n387), .A2(new_n390), .A3(new_n394), .A4(new_n391), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(G101), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(G101), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT81), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n392), .A2(new_n401), .A3(new_n398), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n396), .B(KEYINPUT4), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n393), .A2(new_n404), .A3(G101), .A4(new_n395), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n227), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n222), .B(new_n249), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n397), .A2(KEYINPUT81), .A3(new_n399), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n401), .B1(new_n392), .B2(new_n398), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n391), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n386), .A2(G107), .ZN(new_n412));
  OAI21_X1  g226(.A(G101), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n246), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n250), .A2(new_n253), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n410), .A2(KEYINPUT10), .A3(new_n413), .A4(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n406), .A2(new_n416), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT82), .B1(new_n241), .B2(new_n245), .ZN(new_n421));
  INV_X1    g235(.A(new_n414), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n410), .B2(new_n413), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT12), .ZN(new_n425));
  XOR2_X1   g239(.A(G110), .B(G140), .Z(new_n426));
  INV_X1    g240(.A(G227), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G953), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n426), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n431));
  AND4_X1   g245(.A1(new_n420), .A2(new_n425), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n406), .A2(new_n416), .A3(new_n419), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n246), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n429), .B1(new_n434), .B2(new_n420), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n385), .B(new_n302), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(G469), .A2(G902), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n420), .A3(new_n429), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n425), .A2(new_n420), .A3(new_n431), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n429), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n436), .B(new_n437), .C1(new_n385), .C2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT9), .B(G234), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G221), .B1(new_n443), .B2(G902), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n332), .A2(new_n384), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n250), .A2(new_n253), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(new_n344), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n226), .A2(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n363), .A2(G224), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n226), .A2(new_n451), .A3(G125), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n455), .B2(new_n457), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n403), .A2(new_n203), .A3(new_n200), .A4(new_n405), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n333), .A2(G116), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(G113), .C1(KEYINPUT5), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n202), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n410), .A3(new_n413), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n462), .A2(KEYINPUT83), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT83), .B1(new_n462), .B2(new_n468), .ZN(new_n470));
  XOR2_X1   g284(.A(G110), .B(G122), .Z(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT84), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT85), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n472), .A3(new_n468), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT6), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n462), .A2(new_n468), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n462), .A2(KEYINPUT83), .A3(new_n468), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n461), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n456), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n458), .B2(new_n459), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n455), .A2(new_n457), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n487), .A3(new_n456), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n410), .A2(new_n413), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n466), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n468), .A2(new_n494), .A3(KEYINPUT87), .ZN(new_n495));
  OR3_X1    g309(.A1(new_n493), .A2(KEYINPUT87), .A3(new_n466), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n472), .B(KEYINPUT8), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n492), .A2(new_n476), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n302), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n450), .B1(new_n486), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n484), .B1(new_n483), .B2(new_n476), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n469), .A2(new_n470), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT6), .B1(new_n503), .B2(new_n473), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n460), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n498), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n489), .B2(new_n491), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n507), .B2(new_n476), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n508), .A3(new_n449), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n448), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n363), .A2(G952), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(G234), .B2(G237), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT21), .B(G898), .Z(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT94), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n302), .B(new_n363), .C1(G234), .C2(G237), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G475), .ZN(new_n522));
  INV_X1    g336(.A(G237), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n363), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n207), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n283), .A2(G143), .A3(G214), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(KEYINPUT88), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT18), .A3(G131), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n359), .B(G146), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT18), .A4(G131), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n386), .ZN(new_n537));
  INV_X1    g351(.A(new_n526), .ZN(new_n538));
  AOI21_X1  g352(.A(G143), .B1(new_n283), .B2(G214), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n525), .A2(new_n228), .A3(new_n526), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n529), .A2(KEYINPUT17), .A3(G131), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n351), .A3(new_n350), .A4(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n535), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n542), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n205), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n550), .A3(new_n351), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n537), .B1(new_n535), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n522), .B(new_n302), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n546), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n535), .A2(new_n545), .ZN(new_n560));
  INV_X1    g374(.A(new_n537), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI211_X1 g376(.A(KEYINPUT89), .B(new_n537), .C1(new_n535), .C2(new_n545), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n302), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G478), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n570));
  INV_X1    g384(.A(G122), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G116), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT90), .ZN(new_n573));
  INV_X1    g387(.A(G116), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G122), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT14), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n575), .B(KEYINPUT91), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT14), .ZN(new_n581));
  OAI21_X1  g395(.A(G107), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n573), .A2(new_n580), .A3(new_n389), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(G128), .B(G143), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(new_n242), .Z(new_n587));
  NAND3_X1  g401(.A1(new_n573), .A2(new_n580), .A3(new_n389), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT92), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n582), .A2(new_n585), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(KEYINPUT13), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n248), .A2(KEYINPUT13), .A3(G143), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n230), .ZN(new_n593));
  INV_X1    g407(.A(new_n242), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n591), .A2(new_n593), .B1(new_n594), .B2(new_n586), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n389), .B1(new_n573), .B2(new_n580), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n583), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n443), .A2(new_n373), .A3(G953), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n590), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n590), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n302), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n570), .B1(new_n601), .B2(KEYINPUT93), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(KEYINPUT93), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n604), .B(new_n302), .C1(new_n599), .C2(new_n600), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n606), .B2(new_n570), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n568), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n446), .A2(new_n521), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n398), .ZN(G3));
  OAI21_X1  g425(.A(G472), .B1(new_n300), .B2(G902), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(new_n307), .B2(new_n300), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n613), .A2(new_n384), .A3(new_n445), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT33), .B1(new_n599), .B2(new_n600), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n590), .A2(new_n597), .ZN(new_n616));
  INV_X1    g430(.A(new_n598), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n590), .A2(new_n597), .A3(new_n598), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n621), .A3(G478), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n569), .B(new_n302), .C1(new_n599), .C2(new_n600), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n569), .A2(new_n302), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT95), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n568), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n520), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n614), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n565), .B2(G475), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT97), .B(new_n522), .C1(new_n564), .C2(new_n302), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT96), .B1(new_n553), .B2(KEYINPUT20), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n554), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n553), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n638));
  OAI22_X1  g452(.A1(new_n634), .A2(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n520), .A2(new_n607), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n614), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n613), .A2(new_n445), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n366), .A2(KEYINPUT36), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n357), .A2(new_n361), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n647), .B(new_n648), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n382), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n379), .A2(new_n380), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n644), .A2(new_n521), .A3(new_n609), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT37), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n353), .ZN(G12));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n505), .A2(new_n449), .A3(new_n508), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n449), .B1(new_n505), .B2(new_n508), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n447), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n634), .A2(new_n635), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n637), .A2(new_n638), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n514), .B1(G900), .B2(new_n518), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n608), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT100), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n331), .A2(G472), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n280), .A2(new_n286), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n298), .A2(new_n299), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n309), .B1(new_n668), .B2(new_n306), .ZN(new_n669));
  AOI211_X1 g483(.A(KEYINPUT32), .B(new_n307), .C1(new_n666), .C2(new_n667), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n664), .A2(new_n671), .A3(new_n652), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n501), .A2(new_n509), .ZN(new_n673));
  INV_X1    g487(.A(new_n662), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n639), .A2(new_n607), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n673), .A2(new_n675), .A3(new_n676), .A4(new_n447), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n441), .A2(new_n444), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n656), .B1(new_n672), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n308), .A2(new_n321), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n651), .B1(new_n682), .B2(new_n665), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n681), .A2(KEYINPUT101), .A3(new_n664), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n662), .B(KEYINPUT39), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT40), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n690), .A2(new_n448), .A3(new_n652), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n673), .B(KEYINPUT38), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n567), .A2(new_n607), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n327), .A2(new_n277), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n296), .B1(new_n285), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(new_n302), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n682), .B1(new_n301), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n691), .A2(new_n692), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND3_X1  g513(.A1(new_n627), .A2(new_n568), .A3(new_n662), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n659), .A3(new_n445), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n683), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  OAI21_X1  g517(.A(new_n302), .B1(new_n432), .B2(new_n435), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n436), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n444), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n332), .A2(new_n384), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n629), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n640), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  OAI21_X1  g527(.A(KEYINPUT102), .B1(new_n659), .B2(new_n707), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n705), .A2(new_n444), .A3(new_n436), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n510), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n519), .A3(new_n609), .A4(new_n683), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  XNOR2_X1  g534(.A(new_n306), .B(KEYINPUT103), .ZN(new_n721));
  OR3_X1    g535(.A1(new_n328), .A2(KEYINPUT104), .A3(new_n271), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT104), .B1(new_n328), .B2(new_n271), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n722), .A2(new_n286), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n721), .B1(new_n724), .B2(new_n320), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n612), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n384), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n510), .A2(new_n693), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n519), .A4(new_n716), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  INV_X1    g544(.A(new_n700), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n726), .A2(new_n651), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n659), .A2(new_n707), .A3(KEYINPUT102), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n715), .B1(new_n510), .B2(new_n716), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  INV_X1    g551(.A(new_n384), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n673), .A2(new_n448), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n671), .A2(new_n738), .A3(new_n678), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n737), .B1(new_n740), .B2(new_n700), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT105), .B(new_n737), .C1(new_n740), .C2(new_n700), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n682), .A2(KEYINPUT106), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n308), .A2(new_n321), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n665), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n700), .A2(new_n445), .ZN(new_n749));
  AND4_X1   g563(.A1(KEYINPUT42), .A2(new_n748), .A3(new_n738), .A4(new_n749), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n743), .A2(new_n744), .B1(new_n750), .B2(new_n739), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n228), .ZN(G33));
  NOR2_X1   g566(.A1(new_n740), .A2(new_n663), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n230), .ZN(G36));
  INV_X1    g568(.A(new_n739), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n627), .A2(new_n567), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n613), .A3(new_n652), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n440), .B(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(G469), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n437), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n765), .B(G469), .C1(new_n762), .C2(G902), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n436), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n444), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n687), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n761), .B(new_n769), .C1(new_n760), .C2(new_n759), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n444), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n700), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n332), .A3(new_n384), .A4(new_n739), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  AND3_X1   g591(.A1(new_n758), .A2(new_n513), .A3(new_n727), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n692), .A2(new_n447), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n716), .A3(new_n779), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n780), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n781));
  INV_X1    g595(.A(new_n706), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n773), .B(new_n774), .C1(new_n444), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n739), .A3(new_n778), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n755), .A2(new_n707), .A3(new_n514), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n697), .A2(new_n384), .ZN(new_n786));
  INV_X1    g600(.A(new_n627), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n567), .A4(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n789));
  AND4_X1   g603(.A1(new_n513), .A2(new_n758), .A3(new_n716), .A4(new_n739), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n780), .A2(new_n789), .B1(new_n732), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n781), .A2(new_n784), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n512), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n748), .A2(new_n738), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n785), .A2(new_n786), .A3(new_n568), .A4(new_n627), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n794), .A2(new_n795), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n778), .A2(new_n718), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n719), .A2(new_n712), .A3(new_n709), .A4(new_n729), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n743), .A2(new_n744), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n750), .A2(new_n739), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n610), .A2(new_n653), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n608), .A2(new_n639), .A3(new_n674), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n445), .B1(new_n812), .B2(KEYINPUT108), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n671), .C1(KEYINPUT108), .C2(new_n812), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n749), .A2(new_n612), .A3(new_n725), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n652), .A3(new_n739), .ZN(new_n817));
  INV_X1    g631(.A(new_n753), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n609), .B1(new_n787), .B2(new_n568), .ZN(new_n819));
  MUX2_X1   g633(.A(new_n628), .B(new_n819), .S(KEYINPUT107), .Z(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n521), .A3(new_n614), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n811), .A2(new_n817), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n735), .A2(new_n702), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n680), .B2(new_n684), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n662), .B(KEYINPUT109), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n652), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n697), .A3(new_n678), .A4(new_n728), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT52), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n700), .B1(new_n714), .B2(new_n717), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n830), .A2(new_n732), .B1(new_n683), .B2(new_n701), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n685), .A2(KEYINPUT52), .A3(new_n831), .A4(new_n828), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n810), .B(new_n823), .C1(new_n829), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n810), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n676), .B1(new_n510), .B2(new_n675), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n332), .A3(new_n651), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT101), .B1(new_n840), .B2(new_n681), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n672), .A2(new_n656), .A3(new_n679), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n831), .B(new_n828), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n822), .B1(new_n845), .B2(new_n832), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT110), .B1(new_n751), .B2(new_n807), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n838), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n810), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n836), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n801), .A2(KEYINPUT113), .A3(new_n803), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n806), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  INV_X1    g671(.A(new_n692), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n786), .A2(new_n858), .A3(new_n447), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n860));
  INV_X1    g674(.A(new_n756), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n444), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n856), .A2(new_n857), .B1(new_n859), .B2(new_n863), .ZN(G75));
  NOR2_X1   g678(.A1(new_n502), .A2(new_n504), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(new_n460), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT55), .Z(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n302), .B1(new_n836), .B2(new_n848), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n869), .B2(G210), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n363), .A2(G952), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT115), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  INV_X1    g689(.A(G210), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n876), .B(new_n302), .C1(new_n836), .C2(new_n848), .ZN(new_n877));
  OAI211_X1 g691(.A(KEYINPUT114), .B(new_n867), .C1(new_n877), .C2(KEYINPUT56), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n872), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT116), .A4(new_n878), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(G51));
  XNOR2_X1  g697(.A(new_n849), .B(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n437), .A2(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n437), .A2(KEYINPUT57), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n886), .A2(new_n887), .B1(new_n435), .B2(new_n432), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n869), .A2(G469), .A3(new_n762), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n873), .B1(new_n888), .B2(new_n889), .ZN(G54));
  NAND3_X1  g704(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n546), .A2(new_n552), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n873), .ZN(G60));
  XNOR2_X1  g708(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n624), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n615), .A2(new_n621), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT117), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n884), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n850), .B2(new_n853), .ZN(new_n901));
  INV_X1    g715(.A(new_n898), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n874), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n884), .A2(new_n904), .A3(new_n896), .A4(new_n898), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n900), .A2(new_n903), .A3(new_n905), .ZN(G63));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT60), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n849), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n849), .B2(new_n909), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n649), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n849), .A2(new_n909), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n915));
  INV_X1    g729(.A(new_n381), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n910), .ZN(new_n917));
  INV_X1    g731(.A(new_n874), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n913), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n913), .A2(new_n917), .A3(KEYINPUT61), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(G66));
  NAND2_X1  g737(.A1(new_n516), .A2(G224), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G953), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n811), .A2(new_n821), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n807), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n927), .B2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n865), .B1(G898), .B2(new_n363), .ZN(new_n929));
  XOR2_X1   g743(.A(KEYINPUT121), .B(KEYINPUT122), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n928), .B(new_n931), .ZN(G69));
  OAI21_X1  g746(.A(new_n289), .B1(new_n293), .B2(KEYINPUT30), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n548), .A2(new_n549), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n776), .A2(new_n818), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n751), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n796), .A2(new_n769), .A3(new_n728), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n770), .A2(new_n825), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n937), .B(new_n938), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n939), .B(KEYINPUT123), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n944), .A2(new_n945), .A3(new_n937), .A4(new_n938), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n935), .B1(new_n947), .B2(new_n363), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n427), .A2(G900), .A3(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n698), .A2(new_n825), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n332), .A2(new_n384), .ZN(new_n954));
  INV_X1    g768(.A(new_n689), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n820), .A2(new_n954), .A3(new_n955), .A4(new_n739), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n953), .A2(new_n770), .A3(new_n776), .A4(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n951), .B(new_n935), .C1(new_n957), .C2(G953), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n950), .A2(new_n958), .ZN(G72));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  INV_X1    g775(.A(new_n927), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n323), .B(KEYINPUT125), .Z(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n285), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n836), .A2(new_n852), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n324), .A2(new_n296), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n961), .A3(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n965), .B(new_n968), .C1(G952), .C2(new_n363), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n943), .A2(new_n927), .A3(new_n946), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n971), .A3(new_n961), .ZN(new_n972));
  INV_X1    g786(.A(new_n964), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n972), .A2(new_n286), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n961), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n969), .B1(new_n974), .B2(new_n976), .ZN(G57));
endmodule


