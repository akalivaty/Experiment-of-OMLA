//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n438, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G132), .A4(new_n438), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  INV_X1    g036(.A(G2106), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(new_n455), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n468), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n472), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n476), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(new_n488));
  INV_X1    g063(.A(new_n473), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n468), .A2(new_n470), .A3(G2105), .A4(new_n472), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT70), .Z(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(G114), .B2(new_n471), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n473), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n503));
  AND4_X1   g078(.A1(new_n471), .A2(new_n503), .A3(new_n477), .A4(new_n472), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n502), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT72), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n518), .A3(new_n514), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n507), .A2(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n522), .B1(new_n528), .B2(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n522), .A3(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n521), .B1(new_n530), .B2(new_n531), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n518), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n524), .B2(new_n525), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT74), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n509), .A2(new_n512), .B1(new_n508), .B2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G51), .A3(G543), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT75), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT75), .B1(new_n538), .B2(new_n540), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n513), .A2(G89), .A3(new_n518), .A4(new_n514), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n544), .A2(new_n543), .A3(new_n546), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n541), .A2(new_n542), .B1(new_n547), .B2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND4_X1  g125(.A1(new_n513), .A2(G52), .A3(G543), .A4(new_n514), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n513), .A2(G90), .A3(new_n518), .A4(new_n514), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n516), .B2(new_n517), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT77), .B(new_n557), .C1(new_n526), .C2(new_n555), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(G651), .A3(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n553), .A2(KEYINPUT78), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT78), .B1(new_n553), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  NAND2_X1  g140(.A1(G68), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G56), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n526), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n539), .A2(G43), .A3(G543), .ZN(new_n570));
  INV_X1    g145(.A(G81), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n519), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G188));
  AOI22_X1  g154(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n511), .ZN(new_n581));
  INV_X1    g156(.A(G91), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT79), .B1(new_n519), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n539), .A2(new_n584), .A3(G91), .A4(new_n518), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n514), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT9), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(new_n515), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G50), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n513), .A2(new_n518), .A3(new_n514), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G88), .ZN(new_n593));
  INV_X1    g168(.A(new_n531), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n591), .B(new_n593), .C1(new_n594), .C2(new_n529), .ZN(G303));
  NAND4_X1  g170(.A1(new_n513), .A2(G87), .A3(new_n518), .A4(new_n514), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n513), .A2(G49), .A3(G543), .A4(new_n514), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G288));
  AND2_X1   g175(.A1(G48), .A2(G543), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n513), .A2(new_n514), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT81), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n539), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(G61), .B1(new_n524), .B2(new_n525), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT80), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G61), .C1(new_n524), .C2(new_n525), .ZN(new_n610));
  NAND2_X1  g185(.A1(G73), .A2(G543), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n592), .A2(G86), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n606), .A2(new_n613), .A3(new_n614), .ZN(G305));
  NAND2_X1  g190(.A1(new_n590), .A2(G47), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT82), .B(G85), .Z(new_n618));
  OAI221_X1 g193(.A(new_n616), .B1(new_n511), .B2(new_n617), .C1(new_n519), .C2(new_n618), .ZN(G290));
  INV_X1    g194(.A(G92), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n621));
  OR3_X1    g196(.A1(new_n519), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n519), .B2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n526), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G651), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n539), .A2(G54), .A3(G543), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n622), .A2(new_n623), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G171), .B2(G868), .ZN(G284));
  XOR2_X1   g206(.A(G284), .B(KEYINPUT84), .Z(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(G299), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G168), .B2(new_n633), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(G168), .B2(new_n633), .ZN(G280));
  INV_X1    g211(.A(new_n629), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G860), .ZN(G148));
  OAI21_X1  g214(.A(KEYINPUT85), .B1(new_n573), .B2(G868), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n629), .A2(G559), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(new_n633), .ZN(new_n642));
  MUX2_X1   g217(.A(new_n640), .B(KEYINPUT85), .S(new_n642), .Z(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n489), .A2(G135), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n471), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n492), .A2(KEYINPUT87), .A3(G123), .ZN(new_n648));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n492), .B2(G123), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n645), .B1(new_n646), .B2(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT12), .Z(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT13), .Z(new_n655));
  NAND2_X1  g230(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(KEYINPUT86), .B2(G2100), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n657), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n651), .A2(new_n652), .A3(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT89), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2430), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(KEYINPUT14), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT90), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2451), .B(G2454), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G14), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n675), .B2(new_n678), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(G401));
  XNOR2_X1  g258(.A(G2084), .B(G2090), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT92), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n687), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT17), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G2072), .A2(G2078), .ZN(new_n694));
  OAI22_X1  g269(.A1(new_n688), .A2(new_n692), .B1(new_n444), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G2096), .B(G2100), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n701), .B2(new_n707), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1991), .B(G1996), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n711), .ZN(new_n715));
  INV_X1    g290(.A(new_n713), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n710), .A2(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1981), .B(G1986), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n714), .B2(new_n718), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(G229));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G22), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1971), .ZN(new_n726));
  MUX2_X1   g301(.A(G6), .B(G305), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT32), .B(G1981), .Z(new_n729));
  AOI21_X1  g304(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n723), .A2(G23), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n599), .B2(new_n723), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT96), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT33), .ZN(new_n735));
  INV_X1    g310(.A(G1976), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(KEYINPUT33), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR3_X1    g315(.A1(new_n731), .A2(new_n740), .A3(KEYINPUT34), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT34), .B1(new_n731), .B2(new_n740), .ZN(new_n742));
  OR2_X1    g317(.A1(G16), .A2(G24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G290), .B2(new_n723), .ZN(new_n744));
  INV_X1    g319(.A(G1986), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  OR3_X1    g322(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT97), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n492), .A2(G119), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G107), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n489), .B2(G131), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT93), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n749), .A2(KEYINPUT93), .A3(new_n753), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G25), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n758), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT35), .B(G1991), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n766), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n762), .A2(new_n768), .A3(new_n764), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n748), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n741), .A2(new_n742), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n772), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n741), .A2(new_n774), .A3(new_n742), .A4(new_n770), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n492), .A2(G129), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n489), .A2(G141), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT100), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(new_n759), .ZN(new_n783));
  OAI21_X1  g358(.A(KEYINPUT101), .B1(G29), .B2(G32), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT102), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n782), .A2(KEYINPUT101), .A3(new_n759), .ZN(new_n788));
  OR3_X1    g363(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(new_n785), .B2(new_n788), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT30), .B(G28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(new_n759), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(new_n650), .C2(new_n759), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT104), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n789), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n723), .A2(G19), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n573), .B2(new_n723), .ZN(new_n798));
  INV_X1    g373(.A(G2084), .ZN(new_n799));
  INV_X1    g374(.A(G34), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n800), .B2(KEYINPUT24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT24), .B2(new_n800), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n484), .B2(new_n759), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n798), .A2(G1341), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n723), .A2(G4), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n637), .B2(new_n723), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1348), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n804), .B(new_n807), .C1(G1341), .C2(new_n798), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n759), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT28), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n492), .A2(G128), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(G116), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n489), .B2(G140), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(G29), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G2067), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n759), .A2(G35), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G162), .B2(new_n759), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT29), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G2090), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n803), .A2(new_n799), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT105), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n759), .A2(G33), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT25), .Z(new_n827));
  INV_X1    g402(.A(G139), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n473), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n477), .A2(new_n472), .A3(G127), .ZN(new_n830));
  INV_X1    g405(.A(G115), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n467), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n471), .B1(new_n832), .B2(KEYINPUT99), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n825), .B1(new_n835), .B2(new_n759), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2072), .ZN(new_n837));
  NOR2_X1   g412(.A1(G27), .A2(G29), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G164), .B2(G29), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2078), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n824), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n808), .A2(new_n818), .A3(new_n822), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(G5), .A2(G16), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G171), .B2(G16), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1961), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n723), .A2(G21), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G168), .B2(new_n723), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT103), .B(G1966), .Z(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(new_n848), .Z(new_n849));
  NOR2_X1   g424(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n723), .A2(G20), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT23), .Z(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G299), .B2(G16), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G1956), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n850), .B(new_n854), .C1(G2090), .C2(new_n821), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n796), .A2(new_n842), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n773), .A2(new_n775), .A3(new_n856), .ZN(G311));
  NAND3_X1  g432(.A1(new_n773), .A2(new_n775), .A3(new_n856), .ZN(G150));
  NAND2_X1  g433(.A1(new_n572), .A2(KEYINPUT107), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n592), .A2(G81), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n570), .A4(new_n569), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n511), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n592), .A2(G93), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT106), .B(G55), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n590), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n859), .A2(new_n867), .A3(new_n869), .A4(new_n862), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n637), .A2(G559), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g452(.A(G860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n870), .A2(G860), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(new_n650), .B(new_n494), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n484), .B(KEYINPUT108), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n816), .A2(G164), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n492), .A2(G130), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n489), .A2(G142), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n470), .A2(new_n472), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(G138), .A3(new_n471), .A4(new_n468), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n504), .B1(new_n893), .B2(KEYINPUT4), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n811), .B(new_n815), .C1(new_n894), .C2(new_n500), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n886), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n891), .B1(new_n886), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n900));
  INV_X1    g475(.A(new_n756), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n754), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n756), .ZN(new_n903));
  INV_X1    g478(.A(new_n654), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n654), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n898), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n781), .A2(new_n835), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n782), .B2(new_n835), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n907), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n907), .B2(new_n911), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n885), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n913), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n883), .B(new_n884), .Z(new_n920));
  NAND3_X1  g495(.A1(new_n907), .A2(new_n911), .A3(new_n914), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g500(.A1(new_n873), .A2(new_n641), .ZN(new_n926));
  NAND2_X1  g501(.A1(G299), .A2(new_n629), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n623), .A2(new_n627), .A3(new_n628), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n928), .A2(new_n588), .A3(new_n586), .A4(new_n622), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n873), .A2(new_n641), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n926), .A2(new_n935), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT41), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n936), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(G288), .ZN(new_n944));
  XNOR2_X1  g519(.A(G166), .B(G305), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n944), .B(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n943), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n943), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n870), .A2(new_n633), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n538), .A2(new_n540), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT75), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT75), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n548), .A2(new_n547), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n960), .B(new_n961), .C1(new_n562), .C2(new_n563), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n553), .A2(KEYINPUT78), .A3(new_n561), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n553), .A2(new_n561), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT78), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(G286), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n873), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n962), .A2(new_n871), .A3(new_n967), .A4(new_n872), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(KEYINPUT112), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n871), .A2(new_n872), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n962), .A4(new_n967), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n930), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n941), .B1(new_n970), .B2(new_n969), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n947), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n934), .A2(new_n969), .A3(new_n970), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n939), .A2(new_n940), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n983), .A3(new_n974), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n934), .A2(new_n969), .A3(KEYINPUT113), .A4(new_n970), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n946), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n978), .A2(new_n979), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n946), .B1(new_n975), .B2(new_n976), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n979), .B1(new_n978), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n955), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n976), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n971), .A2(new_n974), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n992), .B(new_n947), .C1(new_n993), .C2(new_n930), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n987), .A2(new_n923), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n978), .A2(new_n979), .A3(new_n989), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(KEYINPUT44), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n995), .B2(KEYINPUT43), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n991), .B1(new_n999), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n1002), .A2(new_n606), .A3(new_n613), .A4(new_n614), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n612), .A2(G651), .B1(new_n592), .B2(G86), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1005), .B2(new_n606), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1002), .A3(new_n606), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(KEYINPUT49), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n502), .A2(new_n505), .ZN(new_n1012));
  INV_X1    g587(.A(new_n500), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  NOR4_X1   g590(.A1(new_n475), .A2(new_n480), .A3(new_n1015), .A4(new_n482), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1011), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1007), .A2(new_n1010), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1007), .A2(new_n1010), .A3(KEYINPUT119), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n599), .A2(new_n736), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT120), .Z(new_n1024));
  AOI21_X1  g599(.A(new_n1003), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1017), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n599), .A2(G1976), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1017), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n599), .B2(G1976), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n1032));
  AOI221_X4 g607(.A(new_n1011), .B1(new_n599), .B2(G1976), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(KEYINPUT118), .A3(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1022), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(G164), .B2(G1384), .ZN(new_n1039));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT45), .B(new_n1040), .C1(new_n894), .C2(new_n500), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1041), .A3(new_n1016), .ZN(new_n1042));
  INV_X1    g617(.A(G1971), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1040), .C1(new_n894), .C2(new_n500), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n1016), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n1051));
  NOR3_X1   g626(.A1(G166), .A2(new_n1051), .A3(new_n1011), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT117), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(G166), .B2(new_n1011), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1050), .A2(G8), .A3(new_n1054), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1025), .A2(new_n1026), .B1(new_n1037), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1045), .A2(new_n1016), .A3(new_n1047), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1062), .A2(new_n1048), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1063), .B2(new_n1011), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1022), .A2(new_n1064), .A3(new_n1036), .A4(new_n1059), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1042), .A2(new_n848), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1045), .A2(new_n1047), .A3(new_n799), .A4(new_n1016), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1011), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G168), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT121), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT63), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT121), .B(new_n1072), .C1(new_n1065), .C2(new_n1069), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1060), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1039), .A2(new_n1041), .A3(new_n1076), .A4(new_n1016), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1045), .A2(new_n1047), .A3(new_n1016), .ZN(new_n1078));
  INV_X1    g653(.A(G1961), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1075), .A2(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n476), .A2(G40), .A3(new_n481), .A4(new_n483), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1040), .B1(new_n894), .B2(new_n500), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1038), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(KEYINPUT53), .A3(new_n1076), .A4(new_n1041), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1065), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1066), .A2(new_n1088), .A3(new_n1067), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1089), .A2(new_n1090), .A3(G286), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n1011), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G286), .A2(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1092), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1091), .A2(new_n1094), .B1(new_n1068), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT125), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1066), .A2(new_n1088), .A3(new_n1067), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT62), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1068), .A2(new_n1096), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(G168), .A3(new_n1100), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1093), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1101), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1087), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n586), .A2(new_n588), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n586), .B2(new_n588), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1083), .A2(new_n1041), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1956), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1078), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1113), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1111), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1081), .B1(new_n1082), .B2(KEYINPUT50), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1956), .B1(new_n1122), .B2(new_n1047), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1041), .A2(new_n1039), .A3(new_n1016), .A4(new_n1115), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G2067), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1014), .A2(new_n1128), .A3(new_n1016), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1348), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1078), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n629), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1119), .B1(new_n1126), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1131), .A2(new_n629), .A3(new_n1133), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT60), .B1(new_n1136), .B2(new_n1134), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n629), .A2(KEYINPUT60), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1131), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1125), .A2(new_n1140), .A3(new_n1119), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n1125), .B2(new_n1119), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1137), .B(new_n1139), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1129), .A2(new_n1130), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1042), .A2(G1996), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n573), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1144), .B(new_n1145), .C1(new_n1150), .C2(KEYINPUT124), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT59), .B1(new_n1150), .B2(new_n1144), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1014), .A2(new_n1128), .A3(new_n1016), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n1146), .ZN(new_n1155));
  INV_X1    g730(.A(G1996), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1083), .A2(new_n1156), .A3(new_n1041), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n572), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1151), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1135), .B1(new_n1143), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(KEYINPUT54), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1080), .A2(G301), .A3(new_n1084), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1086), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1077), .A2(new_n1075), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT127), .B1(new_n562), .B2(new_n563), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1084), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT54), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1166), .A2(new_n1065), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1162), .A2(new_n1163), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1074), .A2(new_n1109), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1039), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1016), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n757), .B(new_n766), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n1180), .B2(new_n1179), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n816), .B(new_n1127), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n781), .A2(G1996), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1178), .A2(G1996), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT115), .ZN(new_n1187));
  INV_X1    g762(.A(new_n782), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1185), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1182), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1178), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G290), .B(G1986), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1176), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n757), .A2(new_n768), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n816), .A2(G2067), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1191), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1178), .A2(G1986), .A3(G290), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT48), .Z(new_n1200));
  NAND3_X1  g775(.A1(new_n1182), .A2(new_n1189), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1187), .B(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT47), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1183), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1191), .B1(new_n1205), .B2(new_n781), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1204), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1198), .B(new_n1201), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1194), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g786(.A1(G227), .A2(new_n464), .ZN(new_n1213));
  OAI21_X1  g787(.A(new_n1213), .B1(new_n720), .B2(new_n721), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1214), .B1(new_n680), .B2(new_n682), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n924), .B(new_n1215), .C1(new_n988), .C2(new_n990), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


