

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587;

  XNOR2_X1 U321 ( .A(n335), .B(n334), .ZN(n580) );
  XNOR2_X1 U322 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X2 U323 ( .A1(n533), .A2(n446), .ZN(n563) );
  XNOR2_X1 U324 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U325 ( .A(KEYINPUT38), .B(n475), .ZN(n499) );
  XNOR2_X1 U326 ( .A(n415), .B(n307), .ZN(n533) );
  INV_X1 U327 ( .A(KEYINPUT25), .ZN(n457) );
  XOR2_X1 U328 ( .A(G99GAT), .B(G85GAT), .Z(n371) );
  INV_X1 U329 ( .A(KEYINPUT20), .ZN(n297) );
  XNOR2_X1 U330 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U331 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U332 ( .A(n328), .B(n327), .ZN(n330) );
  XNOR2_X1 U333 ( .A(n300), .B(n299), .ZN(n304) );
  OR2_X1 U334 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U335 ( .A(n386), .B(n385), .ZN(n390) );
  XNOR2_X1 U336 ( .A(n471), .B(KEYINPUT91), .ZN(n484) );
  INV_X1 U337 ( .A(G43GAT), .ZN(n476) );
  XNOR2_X1 U338 ( .A(n447), .B(G190GAT), .ZN(n448) );
  XNOR2_X1 U339 ( .A(n476), .B(KEYINPUT40), .ZN(n477) );
  XNOR2_X1 U340 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT80), .B(G134GAT), .Z(n290) );
  XNOR2_X1 U343 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n289) );
  XNOR2_X1 U344 ( .A(n290), .B(n289), .ZN(n291) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(n291), .ZN(n415) );
  XOR2_X1 U346 ( .A(KEYINPUT81), .B(G183GAT), .Z(n293) );
  XNOR2_X1 U347 ( .A(G15GAT), .B(G176GAT), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n357) );
  XOR2_X1 U350 ( .A(G99GAT), .B(KEYINPUT83), .Z(n295) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U353 ( .A(n357), .B(n296), .Z(n300) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XOR2_X1 U355 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n302) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n315) );
  XNOR2_X1 U358 ( .A(n315), .B(KEYINPUT82), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n306), .B(n305), .Z(n307) );
  XOR2_X1 U361 ( .A(G36GAT), .B(G190GAT), .Z(n372) );
  XOR2_X1 U362 ( .A(G64GAT), .B(G92GAT), .Z(n309) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G204GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n359) );
  XOR2_X1 U365 ( .A(n372), .B(n359), .Z(n311) );
  NAND2_X1 U366 ( .A1(G226GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U368 ( .A(G8GAT), .B(G183GAT), .Z(n320) );
  XOR2_X1 U369 ( .A(n312), .B(n320), .Z(n317) );
  XOR2_X1 U370 ( .A(G211GAT), .B(KEYINPUT21), .Z(n314) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n429) );
  XNOR2_X1 U373 ( .A(n315), .B(n429), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n521) );
  XOR2_X1 U375 ( .A(G211GAT), .B(G71GAT), .Z(n319) );
  XNOR2_X1 U376 ( .A(G22GAT), .B(G127GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n335) );
  XOR2_X1 U378 ( .A(G57GAT), .B(KEYINPUT13), .Z(n356) );
  XNOR2_X1 U379 ( .A(n356), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(G78GAT), .B(G155GAT), .Z(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n328) );
  XOR2_X1 U382 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n324) );
  XNOR2_X1 U383 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n326) );
  AND2_X1 U385 ( .A1(G231GAT), .A2(G233GAT), .ZN(n325) );
  INV_X1 U386 ( .A(KEYINPUT14), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n333) );
  XNOR2_X1 U388 ( .A(G15GAT), .B(G1GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n331), .B(KEYINPUT71), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(KEYINPUT15), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G22GAT), .Z(n426) );
  XOR2_X1 U393 ( .A(n336), .B(n426), .Z(n338) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G50GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n351) );
  XOR2_X1 U396 ( .A(G8GAT), .B(G113GAT), .Z(n340) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G197GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U399 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n342) );
  XNOR2_X1 U400 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U403 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n346) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT73), .B(n347), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U409 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n353) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(G29GAT), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U412 ( .A(KEYINPUT7), .B(n354), .ZN(n384) );
  XNOR2_X1 U413 ( .A(n355), .B(n384), .ZN(n570) );
  INV_X1 U414 ( .A(n570), .ZN(n536) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n368) );
  XNOR2_X1 U416 ( .A(G106GAT), .B(G78GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n358), .B(G148GAT), .ZN(n437) );
  XNOR2_X1 U418 ( .A(n437), .B(n359), .ZN(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n361) );
  XNOR2_X1 U420 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n371), .B(n362), .Z(n364) );
  NAND2_X1 U423 ( .A1(G230GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n575) );
  XNOR2_X1 U427 ( .A(n575), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U428 ( .A1(n536), .A2(n555), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT46), .ZN(n370) );
  NOR2_X1 U430 ( .A1(n580), .A2(n370), .ZN(n387) );
  XOR2_X1 U431 ( .A(KEYINPUT10), .B(n371), .Z(n374) );
  XNOR2_X1 U432 ( .A(G218GAT), .B(n372), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U434 ( .A(KEYINPUT76), .B(G92GAT), .Z(n376) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U437 ( .A(n378), .B(n377), .Z(n380) );
  XOR2_X1 U438 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XNOR2_X1 U439 ( .A(G106GAT), .B(n428), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n382) );
  XNOR2_X1 U442 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U444 ( .A(n390), .ZN(n392) );
  INV_X1 U445 ( .A(n392), .ZN(n546) );
  NAND2_X1 U446 ( .A1(n387), .A2(n546), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n388), .B(KEYINPUT47), .ZN(n389) );
  XNOR2_X1 U448 ( .A(KEYINPUT106), .B(n389), .ZN(n401) );
  INV_X1 U449 ( .A(n580), .ZN(n541) );
  NAND2_X1 U450 ( .A1(n390), .A2(KEYINPUT36), .ZN(n394) );
  INV_X1 U451 ( .A(KEYINPUT36), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n392), .A2(n391), .ZN(n393) );
  NAND2_X1 U453 ( .A1(n394), .A2(n393), .ZN(n454) );
  NOR2_X1 U454 ( .A1(n541), .A2(n454), .ZN(n395) );
  XOR2_X1 U455 ( .A(KEYINPUT45), .B(n395), .Z(n396) );
  NOR2_X1 U456 ( .A1(n575), .A2(n396), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n397), .B(KEYINPUT107), .ZN(n398) );
  NOR2_X1 U458 ( .A1(n398), .A2(n570), .ZN(n399) );
  XNOR2_X1 U459 ( .A(KEYINPUT108), .B(n399), .ZN(n400) );
  NOR2_X1 U460 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U461 ( .A(KEYINPUT48), .B(n402), .ZN(n530) );
  NOR2_X1 U462 ( .A1(n521), .A2(n530), .ZN(n403) );
  XNOR2_X1 U463 ( .A(KEYINPUT54), .B(n403), .ZN(n424) );
  XOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT84), .Z(n405) );
  XNOR2_X1 U465 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n436) );
  XOR2_X1 U467 ( .A(G162GAT), .B(n436), .Z(n407) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(n408), .ZN(n423) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G148GAT), .Z(n410) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(G120GAT), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n412) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(G57GAT), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U477 ( .A(n414), .B(n413), .Z(n421) );
  INV_X1 U478 ( .A(n415), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT87), .B(KEYINPUT5), .Z(n417) );
  XNOR2_X1 U480 ( .A(KEYINPUT6), .B(KEYINPUT88), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n519) );
  NAND2_X1 U485 ( .A1(n424), .A2(n519), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n425), .B(KEYINPUT64), .ZN(n569) );
  XNOR2_X1 U487 ( .A(n426), .B(KEYINPUT22), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n427), .B(G204GAT), .ZN(n441) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U493 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n465) );
  NOR2_X1 U499 ( .A1(n569), .A2(n465), .ZN(n445) );
  XNOR2_X1 U500 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n443) );
  INV_X1 U501 ( .A(KEYINPUT55), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U503 ( .A1(n563), .A2(n392), .ZN(n449) );
  XOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n447) );
  NAND2_X1 U505 ( .A1(n563), .A2(n570), .ZN(n452) );
  XOR2_X1 U506 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n450) );
  XNOR2_X1 U507 ( .A(n450), .B(G169GAT), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(G1348GAT) );
  NOR2_X1 U509 ( .A1(n536), .A2(n575), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT75), .B(n453), .Z(n485) );
  INV_X1 U511 ( .A(n519), .ZN(n464) );
  NOR2_X1 U512 ( .A1(n533), .A2(n521), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT90), .ZN(n456) );
  NOR2_X1 U514 ( .A1(n465), .A2(n456), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(n457), .ZN(n462) );
  XOR2_X1 U516 ( .A(KEYINPUT89), .B(KEYINPUT26), .Z(n460) );
  NAND2_X1 U517 ( .A1(n533), .A2(n465), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n568) );
  XNOR2_X1 U519 ( .A(n521), .B(KEYINPUT27), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n568), .A2(n467), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n470) );
  XNOR2_X1 U523 ( .A(KEYINPUT66), .B(KEYINPUT28), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n493) );
  NOR2_X1 U525 ( .A1(n519), .A2(n467), .ZN(n531) );
  NAND2_X1 U526 ( .A1(n531), .A2(n533), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n493), .A2(n468), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n454), .A2(n484), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n541), .A2(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT37), .B(n473), .ZN(n518) );
  NAND2_X1 U531 ( .A1(n485), .A2(n518), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT94), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n499), .A2(n533), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n580), .A2(n563), .ZN(n480) );
  XNOR2_X1 U535 ( .A(KEYINPUT120), .B(G183GAT), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n480), .B(n479), .ZN(G1350GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n482) );
  NAND2_X1 U538 ( .A1(n580), .A2(n546), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n502) );
  NAND2_X1 U541 ( .A1(n485), .A2(n502), .ZN(n494) );
  NOR2_X1 U542 ( .A1(n519), .A2(n494), .ZN(n486) );
  XOR2_X1 U543 ( .A(G1GAT), .B(n486), .Z(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT34), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U545 ( .A1(n521), .A2(n494), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT92), .B(n488), .Z(n489) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n533), .A2(n494), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT35), .B(KEYINPUT93), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n492), .Z(G1326GAT) );
  INV_X1 U552 ( .A(n493), .ZN(n535) );
  NOR2_X1 U553 ( .A1(n535), .A2(n494), .ZN(n495) );
  XOR2_X1 U554 ( .A(G22GAT), .B(n495), .Z(G1327GAT) );
  NOR2_X1 U555 ( .A1(n519), .A2(n499), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n521), .A2(n499), .ZN(n498) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  NOR2_X1 U560 ( .A1(n535), .A2(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT95), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U563 ( .A1(n570), .A2(n555), .ZN(n517) );
  NAND2_X1 U564 ( .A1(n502), .A2(n517), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT97), .B(n503), .Z(n512) );
  NOR2_X1 U566 ( .A1(n512), .A2(n519), .ZN(n507) );
  XOR2_X1 U567 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n505) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n521), .A2(n512), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT99), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n533), .A2(n512), .ZN(n510) );
  XOR2_X1 U575 ( .A(KEYINPUT100), .B(n510), .Z(n511) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n535), .ZN(n516) );
  XOR2_X1 U578 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT102), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n519), .A2(n527), .ZN(n520) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n533), .A2(n527), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT103), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT104), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n535), .A2(n527), .ZN(n528) );
  XOR2_X1 U594 ( .A(n529), .B(n528), .Z(G1339GAT) );
  INV_X1 U595 ( .A(n530), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n549) );
  NOR2_X1 U597 ( .A1(n533), .A2(n549), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n545) );
  NOR2_X1 U599 ( .A1(n536), .A2(n545), .ZN(n537) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  NOR2_X1 U601 ( .A1(n555), .A2(n545), .ZN(n539) );
  XNOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT109), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  NOR2_X1 U605 ( .A1(n541), .A2(n545), .ZN(n543) );
  XNOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT110), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n544), .Z(G1342GAT) );
  NOR2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n568), .A2(n549), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT111), .B(n550), .Z(n560) );
  NAND2_X1 U614 ( .A1(n560), .A2(n570), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT113), .Z(n553) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT112), .B(n554), .Z(n557) );
  INV_X1 U620 ( .A(n555), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n560), .A2(n562), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n580), .A2(n560), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT114), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n392), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XNOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT122), .ZN(n574) );
  XOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .Z(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n584) );
  NAND2_X1 U636 ( .A1(n584), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n577) );
  NAND2_X1 U640 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT123), .Z(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n584), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n587) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n454), .A2(n585), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

