//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n642, new_n643, new_n644, new_n646, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n465), .A2(new_n466), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n464), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n478), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT67), .ZN(G162));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n464), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT69), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n490), .A2(new_n493), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n496), .B(new_n487), .C1(new_n497), .C2(new_n489), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n464), .A2(G138), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n479), .B2(new_n480), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT71), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n501), .B2(KEYINPUT70), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n464), .A2(G138), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(KEYINPUT70), .C1(new_n466), .C2(new_n465), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n476), .B2(new_n500), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n510), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(new_n506), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n499), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT73), .B1(new_n517), .B2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n518), .B1(new_n522), .B2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  AOI211_X1 g099(.A(KEYINPUT73), .B(new_n524), .C1(new_n519), .C2(new_n521), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n516), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n518), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT72), .B(KEYINPUT6), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n530), .B2(new_n524), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n522), .A2(new_n532), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n528), .A2(G88), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G62), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n514), .B2(new_n515), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(G75), .A2(G543), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n531), .B2(new_n533), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n542), .A2(G651), .B1(new_n544), .B2(G50), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n536), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G166));
  NAND2_X1  g125(.A1(new_n528), .A2(new_n535), .ZN(new_n551));
  INV_X1    g126(.A(G89), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n544), .A2(G51), .ZN(new_n554));
  NAND3_X1  g129(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT7), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n553), .A2(new_n558), .ZN(G168));
  AOI21_X1  g134(.A(KEYINPUT74), .B1(new_n534), .B2(new_n516), .ZN(new_n560));
  INV_X1    g135(.A(new_n516), .ZN(new_n561));
  AOI211_X1 g136(.A(new_n527), .B(new_n561), .C1(new_n531), .C2(new_n533), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G90), .ZN(new_n564));
  NAND2_X1  g139(.A1(G77), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G64), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n524), .B1(new_n567), .B2(KEYINPUT77), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(new_n569), .B1(G52), .B2(new_n544), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n564), .A2(new_n570), .ZN(G171));
  NAND2_X1  g146(.A1(new_n563), .A2(G81), .ZN(new_n572));
  NAND2_X1  g147(.A1(G68), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G56), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n561), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n544), .A2(G43), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  NAND4_X1  g154(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(G188));
  AOI22_X1  g159(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n524), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  AND2_X1   g162(.A1(KEYINPUT79), .A2(G53), .ZN(new_n588));
  AND4_X1   g163(.A1(new_n587), .A2(new_n534), .A3(G543), .A4(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n587), .B1(new_n544), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G91), .ZN(new_n592));
  NOR3_X1   g167(.A1(new_n560), .A2(new_n562), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G299));
  NAND2_X1  g170(.A1(new_n564), .A2(new_n570), .ZN(G301));
  INV_X1    g171(.A(G168), .ZN(G286));
  AND3_X1   g172(.A1(new_n536), .A2(new_n548), .A3(new_n545), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n548), .B1(new_n536), .B2(new_n545), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(G303));
  OAI21_X1  g175(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n602));
  AND2_X1   g177(.A1(G49), .A2(G543), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n534), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n602), .B1(new_n534), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n563), .B2(G87), .ZN(new_n610));
  INV_X1    g185(.A(G87), .ZN(new_n611));
  NOR4_X1   g186(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT80), .A4(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n608), .B1(new_n610), .B2(new_n612), .ZN(G288));
  AOI22_X1  g188(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n614), .A2(new_n615), .A3(new_n524), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n614), .B2(new_n524), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n616), .A2(new_n617), .B1(new_n544), .B2(G48), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n528), .A2(G86), .A3(new_n535), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(G305));
  NAND2_X1  g195(.A1(new_n563), .A2(G85), .ZN(new_n621));
  NAND2_X1  g196(.A1(G72), .A2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G60), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n561), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n544), .A2(G47), .B1(G651), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(G301), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n544), .A2(G54), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n524), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n631));
  INV_X1    g206(.A(G92), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n551), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n563), .A2(KEYINPUT10), .A3(G92), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n627), .B1(new_n635), .B2(G868), .ZN(G284));
  OAI21_X1  g211(.A(new_n627), .B1(new_n635), .B2(G868), .ZN(G321));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(G299), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(G168), .ZN(G297));
  OAI21_X1  g215(.A(new_n639), .B1(new_n638), .B2(G168), .ZN(G280));
  INV_X1    g216(.A(new_n635), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n642), .A2(G559), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(G860), .B2(new_n635), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT83), .Z(G148));
  NAND2_X1  g220(.A1(new_n577), .A2(new_n638), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n643), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g222(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g223(.A1(new_n477), .A2(G123), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n481), .A2(G135), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n464), .A2(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT85), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n476), .A2(new_n471), .A3(G2105), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  XOR2_X1   g233(.A(KEYINPUT13), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n660), .ZN(G156));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n675), .A3(G14), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(G401));
  XNOR2_X1  g252(.A(G2084), .B(G2090), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(KEYINPUT18), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT17), .B1(new_n679), .B2(new_n681), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n679), .B2(new_n681), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(KEYINPUT18), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2096), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n693), .A2(new_n694), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(new_n697), .A3(new_n695), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n702), .C1(new_n697), .C2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n706), .A2(new_n707), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n706), .A2(new_n707), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(G229));
  NOR2_X1   g290(.A1(G29), .A2(G35), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G162), .B2(G29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2090), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G32), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT26), .Z(new_n724));
  INV_X1    g299(.A(new_n477), .ZN(new_n725));
  INV_X1    g300(.A(G129), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n722), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n721), .B1(new_n728), .B2(new_n720), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT27), .ZN(new_n730));
  INV_X1    g305(.A(G1996), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n512), .A2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n720), .A2(G27), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n732), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n720), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n477), .A2(G128), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n481), .A2(G140), .ZN(new_n741));
  OR2_X1    g316(.A1(G104), .A2(G2105), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n742), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G2067), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n736), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(G2078), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G168), .A2(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT96), .B2(new_n752), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n737), .B(new_n751), .C1(G1966), .C2(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n719), .B(new_n755), .C1(G1966), .C2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(G16), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n757), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n635), .B2(new_n757), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G171), .A2(new_n757), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G5), .B2(new_n757), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT99), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n481), .A2(G139), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  INV_X1    g348(.A(new_n476), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n774), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n771), .B(new_n773), .C1(new_n775), .C2(new_n464), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT95), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G33), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT94), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  INV_X1    g357(.A(KEYINPUT24), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n720), .B1(new_n783), .B2(G34), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n783), .B2(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G160), .B2(G29), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(G2084), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G2084), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G28), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(new_n720), .C1(new_n790), .C2(G28), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n788), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n654), .A2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT97), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n782), .A2(new_n787), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n767), .A2(new_n768), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n757), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n578), .B2(new_n757), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1341), .Z(new_n801));
  AND4_X1   g376(.A1(new_n770), .A2(new_n797), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n756), .A2(new_n761), .A3(new_n765), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G290), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(new_n757), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n757), .B2(G24), .ZN(new_n806));
  INV_X1    g381(.A(G1986), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n720), .A2(G25), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n477), .A2(G119), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n481), .A2(G131), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n720), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n808), .A2(new_n809), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n618), .A2(new_n619), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G16), .ZN(new_n823));
  OR2_X1    g398(.A1(G6), .A2(G16), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT32), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n823), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1981), .ZN(new_n830));
  NAND2_X1  g405(.A1(G303), .A2(G16), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n757), .A2(G22), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT91), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G1971), .ZN(new_n835));
  INV_X1    g410(.A(G1971), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n835), .A2(KEYINPUT92), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n757), .A2(G23), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT80), .B1(new_n551), .B2(new_n611), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n563), .A2(new_n609), .A3(G87), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n607), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n842), .B1(new_n845), .B2(new_n757), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT33), .B(G1976), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n830), .A2(new_n840), .A3(new_n841), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n821), .B1(new_n849), .B2(KEYINPUT34), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT36), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT36), .B1(new_n855), .B2(new_n850), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n803), .B1(new_n854), .B2(new_n856), .ZN(G311));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n856), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n756), .A2(new_n802), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(new_n761), .A3(new_n765), .A4(new_n859), .ZN(G150));
  NAND2_X1  g435(.A1(new_n635), .A2(G559), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT38), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n563), .A2(G93), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT100), .B(G55), .Z(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n561), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n544), .A2(new_n864), .B1(G651), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n577), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n572), .A2(new_n863), .A3(new_n576), .A4(new_n868), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n862), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  AOI21_X1  g450(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(G145));
  NAND2_X1  g456(.A1(new_n477), .A2(G130), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n481), .A2(G142), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n464), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n815), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT103), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n508), .A2(new_n511), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n488), .A2(new_n494), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n746), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n744), .B(KEYINPUT93), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n508), .A2(new_n511), .A3(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n728), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n728), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n777), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n776), .A3(new_n896), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT102), .ZN(new_n902));
  INV_X1    g477(.A(new_n658), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n904), .B(new_n777), .C1(new_n897), .C2(new_n898), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n889), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n658), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n888), .A3(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n654), .B(G160), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(G162), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT40), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G395));
  NAND2_X1  g496(.A1(G166), .A2(G305), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(G166), .A2(G305), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n922), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G288), .A2(KEYINPUT105), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n845), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G290), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(G290), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n925), .B(new_n928), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT106), .ZN(new_n936));
  INV_X1    g511(.A(new_n932), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n643), .B(new_n873), .Z(new_n941));
  NAND2_X1  g516(.A1(new_n635), .A2(new_n594), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n635), .A2(new_n594), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n943), .A2(KEYINPUT41), .A3(new_n944), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n642), .A2(G299), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n942), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n941), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n940), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n869), .A2(new_n638), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(G295));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n956), .ZN(G331));
  NAND2_X1  g533(.A1(new_n577), .A2(new_n869), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g535(.A1(G301), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n961), .A3(new_n871), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n959), .B2(new_n871), .ZN(new_n964));
  OAI21_X1  g539(.A(G168), .B1(G301), .B2(new_n960), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n965), .ZN(new_n967));
  INV_X1    g542(.A(new_n961), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n870), .B2(new_n872), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n969), .B2(new_n962), .ZN(new_n970));
  OAI22_X1  g545(.A1(new_n966), .A2(new_n970), .B1(new_n947), .B2(new_n950), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n965), .B1(new_n963), .B2(new_n964), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n967), .A3(new_n962), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n945), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(new_n938), .A3(new_n935), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n971), .A2(new_n974), .B1(new_n935), .B2(new_n938), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n966), .A2(new_n970), .ZN(new_n981));
  INV_X1    g556(.A(new_n948), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n949), .A2(new_n942), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n945), .B2(KEYINPUT41), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n974), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n939), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n976), .A4(new_n975), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n979), .A2(new_n980), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n975), .A2(new_n976), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n971), .A2(new_n974), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n939), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n990), .A2(KEYINPUT108), .A3(new_n987), .A4(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n987), .A3(new_n976), .A4(new_n975), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n986), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n997), .B2(new_n977), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n989), .B1(KEYINPUT44), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  NAND4_X1  g576(.A1(G303), .A2(new_n1001), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n547), .A2(G8), .A3(new_n549), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n894), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n470), .A2(new_n473), .ZN(new_n1013));
  INV_X1    g588(.A(G125), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n479), .B2(new_n480), .ZN(new_n1015));
  INV_X1    g590(.A(new_n468), .ZN(new_n1016));
  OAI21_X1  g591(.A(G2105), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1017), .A3(G40), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1011), .A2(new_n1012), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n894), .B2(new_n1009), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n512), .A2(new_n1024), .A3(new_n1009), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1023), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n894), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1022), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n512), .B2(new_n1009), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n836), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1008), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n512), .A2(new_n1009), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n894), .A2(new_n1024), .A3(new_n1009), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1022), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1034), .B1(new_n1042), .B2(G2090), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(G8), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G288), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1010), .A2(new_n1026), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(G1976), .B(new_n608), .C1(new_n610), .C2(new_n612), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1050), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n618), .B2(new_n619), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n618), .A2(new_n619), .A3(new_n1055), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1058), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(new_n1056), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1062), .A3(new_n1050), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1052), .A2(new_n1054), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT45), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1010), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(new_n1022), .A3(new_n1067), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n1068), .A2(G1966), .B1(new_n1042), .B2(G2084), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(G8), .A3(G168), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1037), .A2(new_n1044), .A3(new_n1064), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1044), .A2(new_n1064), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1043), .A2(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1008), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1078), .A2(KEYINPUT117), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1044), .A4(new_n1064), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1075), .A2(new_n1077), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1026), .B1(new_n1010), .B2(new_n1065), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1966), .B1(new_n1087), .B2(new_n1067), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1041), .A2(new_n1022), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1024), .B1(new_n512), .B2(new_n1009), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1089), .A2(G2084), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(G8), .B(G286), .C1(new_n1088), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(G8), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1095), .B(new_n1096), .C1(new_n1049), .C2(G168), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(KEYINPUT51), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(new_n1099), .C1(new_n1069), .C2(G286), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n733), .A2(KEYINPUT53), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(G160), .A2(G40), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1010), .B2(new_n1065), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1031), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(KEYINPUT123), .A3(new_n1031), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n768), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1033), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(new_n733), .A3(new_n1022), .A4(new_n1031), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1112), .A2(G301), .A3(new_n1113), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1087), .A2(new_n1067), .A3(new_n1105), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1032), .A2(G2078), .A3(new_n1033), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1116), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1119), .B(new_n1113), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G171), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1103), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1037), .A2(new_n1044), .A3(new_n1064), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1102), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT57), .B1(new_n591), .B2(new_n593), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n544), .A2(new_n588), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT9), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n544), .A2(new_n587), .A3(new_n588), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n528), .A2(G91), .A3(new_n535), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n586), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1129), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1032), .A2(new_n1033), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1023), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1141));
  INV_X1    g716(.A(G1956), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1137), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1029), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1026), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n1012), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1956), .B1(new_n1147), .B2(new_n1027), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1137), .B1(new_n1148), .B2(new_n1140), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1048), .A2(new_n748), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n764), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n642), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1144), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1048), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT58), .B(G1341), .Z(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1114), .A2(new_n731), .A3(new_n1022), .A4(new_n1031), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n577), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(KEYINPUT118), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1149), .B1(new_n1143), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1163), .ZN(new_n1165));
  NOR4_X1   g740(.A1(new_n1148), .A2(new_n1137), .A3(new_n1140), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT60), .B1(new_n1152), .B2(new_n1151), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n1151), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n635), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n642), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1168), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1154), .B1(new_n1167), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1113), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1179));
  OAI21_X1  g754(.A(G171), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(KEYINPUT125), .B(G171), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1122), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1125), .B1(new_n1185), .B2(G301), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT54), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1184), .A2(new_n1186), .B1(new_n1103), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1128), .A2(new_n1177), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1052), .A2(new_n1063), .A3(new_n1054), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1155), .A2(G8), .ZN(new_n1191));
  NOR2_X1   g766(.A1(G288), .A2(G1976), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1061), .B1(new_n1063), .B2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1044), .A2(new_n1190), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT114), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT62), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n1094), .C2(new_n1101), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1102), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1127), .A2(new_n1123), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1086), .A2(new_n1189), .A3(new_n1195), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT110), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(new_n1066), .B2(new_n1026), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1022), .A2(new_n1010), .A3(KEYINPUT110), .A4(new_n1065), .ZN(new_n1207));
  AND2_X1   g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n746), .B(G2067), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1210), .A2(KEYINPUT111), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(KEYINPUT111), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n727), .B(G1996), .ZN(new_n1213));
  AOI22_X1  g788(.A1(new_n1211), .A2(new_n1212), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n815), .B(new_n818), .ZN(new_n1215));
  XOR2_X1   g790(.A(new_n1215), .B(KEYINPUT112), .Z(new_n1216));
  NAND2_X1  g791(.A1(new_n1208), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(G290), .B(G1986), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1218), .B1(new_n1208), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1204), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1208), .A2(new_n731), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT46), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT47), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1208), .B1(new_n727), .B2(new_n1209), .ZN(new_n1225));
  AND3_X1   g800(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1224), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1208), .A2(new_n807), .A3(new_n804), .ZN(new_n1228));
  XOR2_X1   g803(.A(new_n1228), .B(KEYINPUT48), .Z(new_n1229));
  OAI22_X1  g804(.A1(new_n1226), .A2(new_n1227), .B1(new_n1218), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n816), .A2(new_n818), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1231), .ZN(new_n1232));
  AOI22_X1  g807(.A1(new_n1214), .A2(new_n1232), .B1(new_n748), .B2(new_n893), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1230), .B1(new_n1235), .B2(new_n1208), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1221), .A2(new_n1236), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g812(.A1(new_n917), .A2(new_n918), .ZN(new_n1239));
  OR3_X1    g813(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1240), .B1(new_n711), .B2(new_n714), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n979), .A2(new_n988), .ZN(new_n1242));
  AND3_X1   g816(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .ZN(G308));
  NAND3_X1  g817(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .ZN(G225));
endmodule


