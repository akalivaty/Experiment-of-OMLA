//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  AOI22_X1  g0004(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n204), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT1), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n204), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n212), .B(new_n215), .C1(new_n218), .C2(new_n220), .ZN(G361));
  XNOR2_X1  g0021(.A(G238), .B(G244), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(G232), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT2), .B(G226), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n225), .B(new_n228), .ZN(G358));
  XOR2_X1   g0029(.A(G50), .B(G68), .Z(new_n230));
  XNOR2_X1  g0030(.A(G58), .B(G77), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XNOR2_X1  g0033(.A(G107), .B(G116), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G351));
  INV_X1    g0036(.A(KEYINPUT66), .ZN(new_n237));
  NOR2_X1   g0037(.A1(G41), .A2(G45), .ZN(new_n238));
  OAI21_X1  g0038(.A(new_n237), .B1(new_n238), .B2(G1), .ZN(new_n239));
  INV_X1    g0039(.A(G1), .ZN(new_n240));
  OAI211_X1 g0040(.A(new_n240), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G274), .ZN(new_n243));
  AND2_X1   g0043(.A1(G1), .A2(G13), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT73), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n242), .A2(KEYINPUT73), .A3(new_n246), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT67), .B(G1), .ZN(new_n252));
  INV_X1    g0052(.A(new_n238), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n252), .A2(new_n253), .B1(new_n244), .B2(new_n245), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G238), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(G226), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n267), .A2(KEYINPUT72), .A3(G226), .A4(new_n257), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n262), .A2(new_n268), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n244), .A2(new_n245), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT13), .B1(new_n256), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n249), .A2(new_n250), .B1(G238), .B2(new_n254), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n271), .A2(new_n273), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n264), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(G68), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(G77), .B1(G20), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G50), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n291), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n216), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT11), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G1), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n297), .A2(new_n299), .A3(G13), .A4(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(KEYINPUT12), .A3(new_n283), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT12), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n300), .B2(G68), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n296), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n293), .B1(G20), .B2(new_n252), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G68), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n295), .B2(new_n294), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n275), .A2(G190), .A3(new_n279), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n281), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT14), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n275), .A2(G179), .A3(new_n279), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n309), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n311), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n247), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(G226), .B2(new_n254), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n267), .A2(G222), .A3(new_n257), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n267), .A2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n325), .B1(new_n326), .B2(new_n267), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n273), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n315), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G58), .A2(G68), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n217), .B1(new_n333), .B2(new_n285), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT69), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n287), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n293), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n306), .A2(G50), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n301), .A2(new_n285), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n332), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  INV_X1    g0146(.A(new_n331), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n341), .A2(KEYINPUT9), .A3(new_n342), .A4(new_n343), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT70), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n324), .B2(new_n330), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n347), .A2(G190), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n344), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT10), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n349), .B(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n331), .A2(new_n362), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n363), .A2(new_n352), .A3(new_n353), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT10), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(new_n364), .A3(new_n365), .A4(new_n357), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n348), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n323), .B1(G244), .B2(new_n254), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n267), .A2(G232), .A3(new_n257), .ZN(new_n369));
  INV_X1    g0169(.A(G107), .ZN(new_n370));
  INV_X1    g0170(.A(G238), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n369), .B1(new_n370), .B2(new_n267), .C1(new_n327), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n273), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G200), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n306), .A2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n282), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n379), .B1(new_n217), .B2(new_n326), .C1(new_n287), .C2(new_n336), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n293), .B1(new_n326), .B2(new_n301), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n368), .A2(new_n373), .A3(G190), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n375), .A2(new_n376), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n374), .A2(new_n315), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n376), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n368), .A2(new_n373), .A3(new_n346), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n322), .A2(new_n367), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n337), .A2(new_n300), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n306), .B2(new_n337), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n283), .ZN(new_n395));
  OAI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n333), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n286), .A2(G159), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT74), .B(G33), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n263), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n266), .A2(new_n217), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n259), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n265), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n403), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n402), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n399), .B1(new_n411), .B2(new_n283), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n290), .A2(new_n216), .A3(new_n292), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n217), .B(new_n265), .C1(new_n401), .C2(new_n263), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT7), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT74), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G33), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n264), .A2(KEYINPUT74), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT3), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n421), .A2(new_n403), .A3(new_n217), .A4(new_n265), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(G68), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n398), .A2(new_n413), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n393), .B1(new_n414), .B2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n254), .A2(G232), .B1(new_n242), .B2(new_n246), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n265), .B1(new_n401), .B2(new_n263), .ZN(new_n428));
  MUX2_X1   g0228(.A(G223), .B(G226), .S(G1698), .Z(new_n429));
  AOI22_X1  g0229(.A1(new_n428), .A2(new_n429), .B1(G33), .B2(G87), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n427), .B(new_n362), .C1(new_n430), .C2(new_n272), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n264), .A2(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n418), .A2(G33), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n263), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n429), .B1(new_n435), .B2(new_n259), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G87), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n272), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n252), .A2(new_n253), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(G232), .A3(new_n272), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n247), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n351), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n436), .A2(new_n437), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n273), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n362), .A4(new_n427), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n432), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n426), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n426), .B2(new_n447), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT17), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(G68), .B1(new_n416), .B2(KEYINPUT7), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n433), .A2(new_n434), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n259), .B1(new_n453), .B2(KEYINPUT3), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n403), .B1(new_n454), .B2(new_n217), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n424), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(KEYINPUT7), .B(new_n408), .C1(new_n453), .C2(KEYINPUT3), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT75), .B1(new_n409), .B2(new_n403), .ZN(new_n458));
  AOI211_X1 g0258(.A(new_n406), .B(KEYINPUT7), .C1(new_n265), .C2(new_n408), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n398), .B1(new_n460), .B2(G68), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n293), .B(new_n456), .C1(new_n461), .C2(KEYINPUT16), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n392), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n315), .B1(new_n438), .B2(new_n441), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n427), .B(new_n346), .C1(new_n430), .C2(new_n272), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT76), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT76), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n444), .A2(new_n467), .A3(new_n346), .A4(new_n427), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n463), .B2(new_n469), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT17), .B1(new_n426), .B2(new_n447), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n451), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT79), .B1(new_n390), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n348), .B(new_n388), .C1(new_n359), .C2(new_n366), .ZN(new_n478));
  INV_X1    g0278(.A(new_n476), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n322), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  MUX2_X1   g0284(.A(G257), .B(G264), .S(G1698), .Z(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n435), .B2(new_n259), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n258), .A2(new_n259), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G303), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n272), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n297), .A2(new_n299), .A3(G45), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(G270), .B(new_n272), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n246), .A2(new_n252), .A3(new_n495), .A4(G45), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n297), .A2(new_n299), .A3(G33), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n415), .A2(G116), .A3(new_n300), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n301), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(G20), .B1(G33), .B2(G283), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n264), .A2(G97), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n503), .A2(new_n504), .B1(G20), .B2(new_n501), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n293), .A2(KEYINPUT20), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT20), .B1(new_n293), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n500), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND4_X1   g0308(.A1(new_n484), .A2(new_n498), .A3(G179), .A4(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n489), .A2(new_n497), .A3(new_n346), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n484), .B1(new_n510), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  INV_X1    g0313(.A(new_n508), .ZN(new_n514));
  OAI21_X1  g0314(.A(G169), .B1(new_n489), .B2(new_n497), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n428), .A2(new_n485), .B1(G303), .B2(new_n487), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n496), .B(new_n494), .C1(new_n517), .C2(new_n272), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n508), .A3(KEYINPUT21), .A4(G169), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n498), .A2(G190), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n489), .B2(new_n497), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n512), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G264), .B(new_n272), .C1(new_n490), .C2(new_n493), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n496), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G250), .A2(G1698), .ZN(new_n527));
  INV_X1    g0327(.A(G257), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(G1698), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n435), .B2(new_n259), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n453), .A2(G294), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n272), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n526), .B1(new_n532), .B2(KEYINPUT85), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT85), .ZN(new_n534));
  INV_X1    g0334(.A(G294), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n401), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n428), .B2(new_n529), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n537), .B2(new_n272), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n315), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n496), .B(new_n525), .C1(new_n537), .C2(new_n272), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n346), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n217), .B(new_n544), .C1(new_n435), .C2(new_n259), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n217), .A2(G87), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n542), .B1(new_n487), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n453), .A2(new_n217), .A3(G116), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n217), .B2(G107), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n370), .A2(KEYINPUT23), .A3(G20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT24), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n501), .B1(new_n433), .B2(new_n434), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n217), .B1(new_n551), .B2(new_n552), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT24), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n545), .A2(new_n557), .A3(new_n558), .A4(new_n548), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n415), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n370), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT25), .B1(new_n301), .B2(new_n370), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n292), .A2(new_n216), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n300), .A3(new_n290), .A4(new_n499), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n561), .A2(new_n562), .B1(new_n370), .B2(new_n564), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n539), .A2(new_n541), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n555), .A2(new_n559), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n567), .B2(new_n293), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n528), .A2(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G250), .B2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n421), .B2(new_n265), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT85), .B(new_n273), .C1(new_n571), .C2(new_n536), .ZN(new_n572));
  INV_X1    g0372(.A(new_n526), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n538), .A2(new_n362), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n540), .A2(new_n351), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G257), .B(new_n272), .C1(new_n490), .C2(new_n493), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n496), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n582));
  AND2_X1   g0382(.A1(KEYINPUT4), .A2(G244), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n257), .B(new_n583), .C1(new_n258), .C2(new_n259), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  INV_X1    g0387(.A(G244), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G1698), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n435), .B2(new_n259), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n581), .B(new_n346), .C1(new_n591), .C2(new_n272), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT4), .B1(new_n428), .B2(new_n589), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n273), .B1(new_n595), .B2(new_n586), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT81), .A3(new_n346), .A4(new_n581), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT80), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n287), .A2(new_n326), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT6), .ZN(new_n603));
  INV_X1    g0403(.A(G97), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n602), .A2(new_n603), .B1(new_n370), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n599), .B(new_n601), .C1(new_n606), .C2(new_n217), .ZN(new_n607));
  AND2_X1   g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G97), .A2(G107), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n370), .A2(KEYINPUT6), .A3(G97), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n217), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT80), .B1(new_n612), .B2(new_n600), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n607), .B(new_n613), .C1(new_n411), .C2(new_n370), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n293), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n301), .A2(new_n604), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n564), .B2(new_n604), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n596), .A2(new_n581), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n615), .A2(new_n618), .B1(new_n619), .B2(new_n315), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n590), .A2(new_n587), .ZN(new_n621));
  INV_X1    g0421(.A(new_n586), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n272), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n623), .A2(new_n362), .A3(new_n580), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n351), .B1(new_n596), .B2(new_n581), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n617), .B1(new_n614), .B2(new_n293), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n598), .A2(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n371), .A2(new_n257), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n588), .A2(G1698), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n421), .B2(new_n265), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n273), .B1(new_n632), .B2(new_n556), .ZN(new_n633));
  AND2_X1   g0433(.A1(G33), .A2(G41), .ZN(new_n634));
  OAI21_X1  g0434(.A(G274), .B1(new_n634), .B2(new_n216), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT82), .B1(new_n490), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT82), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n246), .A2(new_n637), .A3(new_n252), .A4(G45), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n272), .A2(G250), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n636), .A2(new_n638), .B1(new_n490), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT19), .B1(new_n282), .B2(G97), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT19), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n217), .B1(new_n269), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n609), .A2(new_n543), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n217), .B(G68), .C1(new_n435), .C2(new_n259), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n415), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n564), .A2(new_n543), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n378), .A2(new_n300), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n633), .A2(new_n640), .A3(G190), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n642), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n564), .A2(new_n377), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n649), .A2(new_n655), .A3(new_n651), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n636), .A2(new_n638), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n639), .A2(new_n490), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n629), .B(new_n630), .C1(new_n435), .C2(new_n259), .ZN(new_n660));
  INV_X1    g0460(.A(new_n556), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n272), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(G169), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n633), .A2(new_n640), .A3(G179), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n656), .B1(new_n665), .B2(KEYINPUT83), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT83), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n663), .A2(new_n667), .A3(new_n664), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n654), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n524), .A2(new_n578), .A3(new_n628), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n483), .A2(new_n670), .ZN(G372));
  NAND3_X1  g0471(.A1(new_n281), .A2(new_n309), .A3(new_n310), .ZN(new_n672));
  INV_X1    g0472(.A(new_n387), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n320), .A2(new_n321), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n451), .A2(new_n475), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n473), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n359), .A2(new_n366), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n348), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n620), .A2(new_n598), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n669), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n656), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n665), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n642), .A2(new_n652), .A3(new_n653), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n620), .A2(new_n684), .A3(new_n598), .A4(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT86), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n633), .A2(G179), .A3(new_n640), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n315), .B1(new_n633), .B2(new_n640), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT83), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n668), .A3(new_n683), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n685), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT26), .B1(new_n693), .B2(new_n680), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n656), .B1(new_n663), .B2(new_n664), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n654), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n681), .A2(new_n696), .A3(new_n679), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT86), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n694), .A2(new_n697), .A3(new_n698), .A4(new_n684), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n577), .A2(new_n685), .A3(new_n684), .ZN(new_n700));
  INV_X1    g0500(.A(new_n566), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n498), .A2(new_n508), .A3(G179), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT84), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n510), .A2(new_n484), .A3(new_n508), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n516), .A3(new_n519), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n700), .B(new_n628), .C1(new_n701), .C2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n688), .A2(new_n699), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n678), .B1(new_n483), .B2(new_n709), .ZN(G369));
  INV_X1    g0510(.A(G13), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n252), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G213), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G343), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n508), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT87), .B1(new_n706), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n521), .A2(new_n514), .A3(new_n522), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n705), .A2(new_n516), .A3(new_n519), .A4(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n706), .A2(KEYINPUT87), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT88), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n727), .B(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n578), .B1(new_n568), .B2(new_n718), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n566), .B2(new_n718), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(G330), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n706), .A2(new_n718), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n566), .A2(new_n577), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n701), .A2(new_n718), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT89), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(KEYINPUT89), .A3(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n732), .A2(new_n741), .ZN(G399));
  INV_X1    g0542(.A(new_n213), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G41), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n646), .A2(G116), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n744), .A2(new_n240), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n220), .B2(new_n744), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n708), .A2(new_n750), .A3(new_n718), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n669), .A2(new_n681), .A3(new_n679), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n695), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n707), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n718), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n623), .A2(new_n580), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n659), .A2(new_n662), .ZN(new_n759));
  INV_X1    g0559(.A(new_n525), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n532), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n758), .A2(new_n759), .A3(new_n761), .A4(new_n510), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT30), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n759), .A2(new_n498), .A3(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n619), .A3(new_n540), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n641), .A2(new_n532), .A3(new_n760), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n767), .A2(KEYINPUT30), .A3(new_n758), .A4(new_n510), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n764), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n719), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT31), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT90), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n670), .B2(new_n719), .ZN(new_n776));
  INV_X1    g0576(.A(new_n625), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n777), .B(new_n627), .C1(new_n362), .C2(new_n619), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n680), .A2(new_n692), .A3(new_n778), .A4(new_n685), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n724), .A2(new_n734), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT90), .A4(new_n718), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n774), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G330), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n757), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n749), .B1(new_n786), .B2(G1), .ZN(G364));
  OR2_X1    g0587(.A1(new_n729), .A2(G330), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n729), .A2(G330), .ZN(new_n789));
  INV_X1    g0589(.A(G45), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n711), .A2(new_n790), .A3(G20), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n240), .B1(new_n791), .B2(KEYINPUT91), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(KEYINPUT91), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n744), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n788), .A2(new_n789), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n217), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n362), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n370), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n267), .B1(new_n800), .B2(new_n543), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT93), .Z(new_n802));
  NOR2_X1   g0602(.A1(G179), .A2(G200), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n217), .B1(new_n803), .B2(G190), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n604), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n217), .A2(G190), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n803), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G159), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n805), .B1(new_n809), .B2(KEYINPUT32), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n346), .A2(G200), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(G20), .A3(G190), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n806), .A2(new_n811), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n813), .A2(G58), .B1(new_n815), .B2(G77), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n810), .B(new_n816), .C1(KEYINPUT32), .C2(new_n809), .ZN(new_n817));
  NAND3_X1  g0617(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G190), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n362), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n283), .B1(new_n822), .B2(new_n285), .ZN(new_n823));
  OR4_X1    g0623(.A1(new_n799), .A2(new_n802), .A3(new_n817), .A4(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT94), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n814), .A2(new_n826), .B1(new_n804), .B2(new_n535), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G326), .B2(new_n821), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT95), .Z(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT33), .B(G317), .Z(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n820), .A2(new_n830), .B1(new_n798), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G322), .ZN(new_n833));
  INV_X1    g0633(.A(G303), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n487), .B1(new_n812), .B2(new_n833), .C1(new_n834), .C2(new_n800), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n832), .B(new_n835), .C1(new_n839), .C2(G329), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n824), .A2(new_n825), .B1(new_n829), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n825), .B2(new_n824), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n216), .B1(G20), .B2(new_n315), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n213), .A2(G355), .A3(new_n267), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n743), .A2(new_n428), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(G45), .B2(new_n219), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n232), .A2(new_n790), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n845), .B1(G116), .B2(new_n213), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(G13), .A2(G33), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT92), .Z(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(G20), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n843), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n795), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT97), .Z(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n727), .B2(new_n852), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n796), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G396));
  NAND2_X1  g0659(.A1(new_n385), .A2(new_n719), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n383), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n387), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n673), .A2(new_n718), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n709), .B2(new_n719), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n388), .A2(new_n719), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n708), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n785), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n794), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  INV_X1    g0671(.A(new_n851), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n843), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT98), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n795), .B1(new_n875), .B2(new_n326), .ZN(new_n876));
  INV_X1    g0676(.A(new_n843), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n813), .A2(G143), .B1(new_n815), .B2(G159), .ZN(new_n878));
  INV_X1    g0678(.A(G137), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n878), .B1(new_n822), .B2(new_n879), .C1(new_n339), .C2(new_n820), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT34), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n428), .B1(new_n285), .B2(new_n800), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n798), .A2(new_n283), .B1(new_n804), .B2(new_n394), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n882), .B(new_n883), .C1(new_n839), .C2(G132), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n822), .A2(new_n834), .B1(new_n814), .B2(new_n501), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(G283), .B2(new_n819), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT99), .Z(new_n887));
  OAI221_X1 g0687(.A(new_n487), .B1(new_n804), .B2(new_n604), .C1(new_n812), .C2(new_n535), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n543), .A2(new_n798), .B1(new_n800), .B2(new_n370), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n888), .B(new_n889), .C1(new_n839), .C2(G311), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n881), .A2(new_n884), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n864), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n876), .B1(new_n877), .B2(new_n891), .C1(new_n892), .C2(new_n851), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n871), .A2(new_n893), .ZN(G384));
  INV_X1    g0694(.A(new_n606), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(G116), .A4(new_n218), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  OAI21_X1  g0699(.A(G77), .B1(new_n394), .B2(new_n283), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n900), .A2(new_n219), .B1(G50), .B2(new_n283), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n252), .A2(G13), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n774), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n779), .A2(new_n734), .A3(new_n724), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT90), .B1(new_n905), .B2(new_n718), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n670), .A2(new_n775), .A3(new_n719), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n321), .B(new_n719), .C1(new_n320), .C2(new_n311), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n319), .A2(new_n317), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n318), .B1(new_n280), .B2(G169), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n321), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n321), .A2(new_n719), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n672), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n864), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n425), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT16), .B1(new_n423), .B2(new_n399), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n392), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n717), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n476), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n432), .A2(new_n442), .A3(new_n446), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT78), .B1(new_n922), .B2(new_n463), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n469), .B2(new_n717), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n426), .A2(new_n447), .A3(new_n448), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n463), .A2(new_n469), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT100), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n463), .B2(new_n717), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n426), .A2(KEYINPUT100), .A3(new_n716), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n923), .A2(new_n927), .A3(new_n925), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n926), .A2(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n921), .B2(new_n934), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n908), .B(new_n915), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT103), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT103), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT102), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n922), .B2(new_n463), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n426), .A2(new_n447), .A3(KEYINPUT102), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT37), .B1(new_n932), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT100), .B1(new_n426), .B2(new_n716), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n463), .A2(new_n929), .A3(new_n717), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n951), .A2(new_n952), .B1(new_n463), .B2(new_n469), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n953), .A2(new_n927), .A3(new_n923), .A4(new_n925), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n930), .A2(new_n931), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n476), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n945), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT104), .B1(new_n935), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n934), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n954), .A2(new_n950), .B1(new_n476), .B2(new_n956), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n961), .C1(new_n962), .C2(new_n945), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n912), .A2(new_n672), .A3(new_n913), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n913), .B1(new_n912), .B2(new_n672), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n892), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n783), .A2(new_n966), .A3(new_n938), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n943), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n482), .A2(new_n908), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(G330), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n473), .A2(new_n717), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n964), .A2(new_n965), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n867), .B2(new_n863), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT38), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n923), .A2(new_n925), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n474), .B1(new_n978), .B2(KEYINPUT17), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n919), .B1(new_n979), .B2(new_n473), .ZN(new_n980));
  INV_X1    g0780(.A(new_n933), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n981), .A2(new_n953), .B1(KEYINPUT37), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n977), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n960), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n974), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT39), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n935), .B2(new_n958), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n320), .A2(new_n321), .A3(new_n718), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(KEYINPUT39), .A3(new_n960), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n757), .A2(new_n482), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n678), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n973), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT106), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n973), .A2(new_n996), .B1(new_n252), .B2(new_n712), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT105), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(KEYINPUT105), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n903), .B1(new_n1001), .B2(new_n1002), .ZN(G367));
  INV_X1    g0803(.A(new_n846), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n228), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n853), .B1(new_n213), .B2(new_n377), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n794), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G159), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n820), .A2(new_n1008), .B1(new_n800), .B2(new_n394), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n804), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(G68), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n487), .B1(new_n808), .B2(G137), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n813), .A2(G150), .B1(new_n815), .B2(G50), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n798), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1014), .A2(G77), .B1(G143), .B2(new_n821), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n822), .A2(new_n826), .B1(new_n798), .B2(new_n604), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G107), .B2(new_n1010), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n815), .A2(G283), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n813), .A2(G303), .B1(new_n808), .B2(G317), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n428), .B1(new_n819), .B2(G294), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT112), .B1(new_n800), .B2(new_n501), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT46), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1016), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT47), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1007), .B1(new_n1026), .B2(new_n843), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n652), .A2(new_n718), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT107), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1029), .A2(new_n654), .A3(new_n695), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n695), .B2(new_n1029), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n852), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1027), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n628), .B1(new_n627), .B2(new_n718), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT108), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n681), .A2(new_n719), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n735), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT42), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1032), .A2(KEYINPUT43), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1040), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n701), .B1(new_n1046), .B2(new_n1037), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n680), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT109), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(KEYINPUT109), .A3(new_n680), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n718), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1044), .A2(new_n1045), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT110), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1044), .A2(new_n1052), .A3(new_n1055), .A4(new_n1045), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1031), .B(KEYINPUT43), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT111), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1041), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n732), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT111), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1054), .A2(new_n1059), .A3(new_n1064), .A4(new_n1056), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n744), .B(KEYINPUT41), .Z(new_n1067));
  INV_X1    g0867(.A(new_n740), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1041), .B1(new_n1068), .B2(new_n738), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT45), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT44), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n741), .B2(new_n1041), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1062), .A2(new_n739), .A3(KEYINPUT44), .A4(new_n740), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n732), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n733), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n736), .B1(new_n731), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n789), .B(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1071), .A2(new_n732), .A3(new_n1075), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1078), .A2(new_n786), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1067), .B1(new_n1084), .B2(new_n786), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1066), .B1(new_n1085), .B2(new_n793), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1063), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1034), .B1(new_n1086), .B2(new_n1087), .ZN(G387));
  AOI211_X1 g0888(.A(G41), .B(new_n743), .C1(new_n1082), .C2(new_n786), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n786), .B2(new_n1082), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n731), .A2(new_n1033), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n813), .A2(G317), .B1(new_n815), .B2(G303), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n822), .B2(new_n833), .C1(new_n826), .C2(new_n820), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT48), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n800), .A2(new_n535), .B1(new_n804), .B2(new_n831), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT113), .Z(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT49), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT49), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n798), .A2(new_n501), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n428), .B(new_n1103), .C1(G326), .C2(new_n808), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n812), .A2(new_n285), .B1(new_n814), .B2(new_n283), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G150), .B2(new_n808), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1010), .A2(new_n378), .B1(G159), .B2(new_n821), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n800), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(G77), .B1(new_n337), .B2(new_n819), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n454), .B1(G97), .B2(new_n1014), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n877), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n846), .B1(new_n225), .B2(new_n790), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n213), .A2(new_n267), .A3(new_n746), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n336), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1117));
  OAI21_X1  g0917(.A(KEYINPUT50), .B1(new_n336), .B2(G50), .ZN(new_n1118));
  AOI21_X1  g0918(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n745), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(G107), .B2(new_n213), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n795), .B(new_n1113), .C1(new_n853), .C2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1082), .A2(new_n793), .B1(new_n1091), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1090), .A2(new_n1124), .ZN(G393));
  AND3_X1   g0925(.A1(new_n1071), .A2(new_n732), .A3(new_n1075), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n732), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n786), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1126), .A2(new_n1127), .B1(new_n1081), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1084), .A2(new_n1129), .A3(new_n744), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1062), .A2(new_n852), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1004), .A2(new_n235), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n853), .B1(new_n604), .B2(new_n213), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n794), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n813), .A2(G311), .B1(G317), .B2(new_n821), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT52), .Z(new_n1137));
  OAI22_X1  g0937(.A1(new_n800), .A2(new_n831), .B1(new_n804), .B2(new_n501), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n799), .B(new_n1138), .C1(G303), .C2(new_n819), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n487), .B1(new_n807), .B2(new_n833), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G294), .B2(new_n815), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1109), .A2(G68), .B1(new_n808), .B2(G143), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT114), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n454), .B1(new_n337), .B2(new_n815), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n804), .A2(new_n326), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n798), .A2(new_n543), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(G50), .C2(new_n819), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n813), .A2(G159), .B1(G150), .B2(new_n821), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT51), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1142), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1135), .B1(new_n1152), .B2(new_n843), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1131), .A2(new_n793), .B1(new_n1132), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1130), .A2(new_n1154), .A3(KEYINPUT115), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT115), .B1(new_n1130), .B2(new_n1154), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1155), .A2(new_n1156), .ZN(G390));
  NOR4_X1   g0957(.A1(new_n783), .A2(new_n975), .A3(new_n784), .A4(new_n864), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n754), .A2(new_n718), .A3(new_n862), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n863), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n785), .A2(new_n892), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n909), .A2(KEYINPUT116), .A3(new_n914), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT116), .B1(new_n909), .B2(new_n914), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n867), .A2(new_n863), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n975), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n785), .B2(new_n892), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1171), .B2(new_n1158), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n994), .B(new_n678), .C1(new_n483), .C2(new_n869), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n990), .B1(new_n1165), .B2(new_n1160), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1177), .A2(new_n959), .A3(new_n963), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1179), .A2(new_n989), .B1(new_n988), .B2(new_n991), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1158), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n988), .A2(new_n991), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n990), .B2(new_n976), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1158), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1177), .A2(new_n959), .A3(new_n963), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1176), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1174), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n744), .A3(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n800), .B2(new_n339), .ZN(new_n1194));
  INV_X1    g0994(.A(G125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n838), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n821), .A2(G128), .ZN(new_n1197));
  INV_X1    g0997(.A(G132), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n267), .C1(new_n1198), .C2(new_n812), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n798), .A2(new_n285), .B1(new_n804), .B2(new_n1008), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1193), .A2(new_n800), .A3(new_n339), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1196), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT54), .B(G143), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n820), .A2(new_n879), .B1(new_n814), .B2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT117), .Z(new_n1205));
  OAI22_X1  g1005(.A1(new_n283), .A2(new_n798), .B1(new_n800), .B2(new_n543), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n487), .B1(new_n814), .B2(new_n604), .C1(new_n501), .C2(new_n812), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n839), .C2(G294), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n820), .A2(new_n370), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1146), .B(new_n1209), .C1(G283), .C2(new_n821), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1202), .A2(new_n1205), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n794), .B1(new_n337), .B2(new_n874), .C1(new_n1211), .C2(new_n877), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1183), .B2(new_n872), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n793), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1192), .A2(new_n1215), .ZN(G378));
  NAND2_X1  g1016(.A1(new_n344), .A2(new_n717), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n367), .B(new_n1217), .Z(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n783), .A2(new_n966), .ZN(new_n1223));
  AOI211_X1 g1023(.A(KEYINPUT103), .B(KEYINPUT40), .C1(new_n985), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n941), .B1(new_n937), .B2(new_n938), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G330), .B(new_n968), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n993), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n968), .A2(G330), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n993), .B1(new_n943), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1222), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n968), .A2(G330), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1227), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n943), .A2(new_n993), .A3(new_n1229), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1222), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1231), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n428), .A2(G41), .ZN(new_n1239));
  INV_X1    g1039(.A(G41), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G50), .B(new_n1239), .C1(new_n264), .C2(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n812), .A2(new_n370), .B1(new_n814), .B2(new_n377), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G68), .B2(new_n1010), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1239), .C1(new_n831), .C2(new_n838), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1109), .A2(G77), .B1(G116), .B2(new_n821), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1014), .A2(G58), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n604), .C2(new_n820), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT58), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT119), .Z(new_n1251));
  OAI22_X1  g1051(.A1(new_n820), .A2(new_n1198), .B1(new_n822), .B2(new_n1195), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n813), .A2(G128), .B1(new_n815), .B2(G137), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n800), .B2(new_n1203), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1252), .B(new_n1254), .C1(G150), .C2(new_n1010), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1257));
  AOI211_X1 g1057(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT59), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1258), .B1(new_n1008), .B2(new_n798), .C1(new_n1255), .C2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1251), .B1(new_n1249), .B2(new_n1248), .C1(new_n1257), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n843), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n795), .B1(new_n285), .B2(new_n873), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n1222), .C2(new_n851), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1264), .A2(KEYINPUT120), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(KEYINPUT120), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1238), .A2(new_n793), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1191), .A2(new_n1175), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1234), .A2(new_n1236), .A3(new_n1235), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1236), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1270));
  OAI211_X1 g1070(.A(KEYINPUT57), .B(new_n1268), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n744), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1268), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1267), .B1(new_n1272), .B2(new_n1273), .ZN(G375));
  NAND2_X1  g1074(.A1(new_n1173), .A2(new_n793), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n839), .A2(G303), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n820), .A2(new_n501), .B1(new_n822), .B2(new_n535), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G97), .B2(new_n1109), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n487), .B1(new_n814), .B2(new_n370), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(G283), .B2(new_n813), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1014), .A2(G77), .B1(new_n1010), .B2(new_n378), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1276), .A2(new_n1278), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n428), .B1(new_n339), .B2(new_n814), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n1246), .B1(new_n285), .B2(new_n804), .C1(new_n1008), .C2(new_n800), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(G128), .C2(new_n839), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT122), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n821), .A2(G132), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1287), .B1(new_n812), .B2(new_n879), .C1(new_n820), .C2(new_n1203), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1282), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n843), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n794), .B1(new_n874), .B2(G68), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT121), .Z(new_n1292));
  OAI211_X1 g1092(.A(new_n1290), .B(new_n1292), .C1(new_n1165), .C2(new_n851), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1275), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1067), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1174), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1176), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT123), .ZN(G381));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1090), .A2(new_n858), .A3(new_n1301), .A4(new_n1124), .ZN(new_n1302));
  OR3_X1    g1102(.A1(G390), .A2(G378), .A3(new_n1302), .ZN(new_n1303));
  OR4_X1    g1103(.A1(G387), .A2(new_n1303), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1104(.A(G378), .ZN(new_n1305));
  INV_X1    g1105(.A(G213), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G343), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G407), .B(G213), .C1(G375), .C2(new_n1308), .ZN(G409));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1267), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1296), .B(new_n1268), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n793), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1305), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1307), .B1(new_n1311), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1297), .A2(KEYINPUT124), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1297), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1176), .A2(new_n744), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(G384), .A3(new_n1295), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1323), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1301), .B1(new_n1327), .B2(new_n1294), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1307), .A2(G2897), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1326), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1310), .B1(new_n1317), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI211_X1 g1136(.A(KEYINPUT127), .B(new_n1310), .C1(new_n1317), .C2(new_n1333), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1317), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1317), .A2(new_n1342), .A3(new_n1339), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1336), .A2(new_n1337), .A3(new_n1341), .A4(new_n1343), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(G393), .B(new_n858), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1347));
  AND2_X1   g1147(.A1(G387), .A2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(G387), .A2(new_n1347), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1346), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(G387), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(G390), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G387), .A2(new_n1347), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1352), .A2(new_n1345), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1344), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT125), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1340), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(KEYINPUT63), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1355), .A2(KEYINPUT61), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT63), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1340), .A2(new_n1357), .A3(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1338), .A2(new_n1329), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1326), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1364));
  AND3_X1   g1164(.A1(new_n1363), .A2(KEYINPUT126), .A3(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT126), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1366));
  OR3_X1    g1166(.A1(new_n1365), .A2(new_n1366), .A3(new_n1317), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1359), .A2(new_n1360), .A3(new_n1362), .A4(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1356), .A2(new_n1368), .ZN(G405));
  NAND2_X1  g1169(.A1(G375), .A2(new_n1305), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1370), .A2(new_n1311), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(new_n1339), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1370), .A2(new_n1311), .A3(new_n1338), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  XNOR2_X1  g1174(.A(new_n1374), .B(new_n1355), .ZN(G402));
endmodule


