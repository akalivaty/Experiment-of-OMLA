//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT72), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n211), .B(new_n203), .C1(new_n207), .C2(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT70), .A3(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n216), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n217), .A2(G183gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(new_n220), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n219), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n213), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n233));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT68), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n204), .B(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT23), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n205), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT23), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT25), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n241), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n239), .A2(KEYINPUT69), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT69), .B1(new_n239), .B2(new_n251), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n204), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n246), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT65), .B(G169gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(KEYINPUT23), .A3(new_n248), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n256), .A2(new_n257), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n230), .B1(new_n254), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G113gat), .ZN(new_n267));
  INV_X1    g066(.A(G113gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G120gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT73), .A3(G134gat), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G127gat), .ZN(new_n277));
  INV_X1    g076(.A(G127gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n265), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n280), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n239), .A2(new_n251), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n239), .A2(new_n251), .A3(KEYINPUT69), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n264), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n225), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n229), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n210), .A3(new_n212), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n280), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT74), .A3(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n295), .ZN(new_n296));
  OR3_X1    g095(.A1(new_n296), .A2(KEYINPUT78), .A3(KEYINPUT34), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT78), .B1(new_n296), .B2(KEYINPUT34), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(KEYINPUT34), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT77), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT74), .B1(new_n293), .B2(new_n294), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n202), .B(new_n280), .C1(new_n288), .C2(new_n292), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n293), .A2(new_n294), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT32), .B1(new_n305), .B2(new_n282), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n305), .B2(new_n282), .ZN(new_n308));
  XNOR2_X1  g107(.A(G15gat), .B(G43gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT75), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G71gat), .ZN(new_n311));
  INV_X1    g110(.A(G99gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n306), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n281), .A2(new_n283), .A3(new_n295), .ZN(new_n317));
  INV_X1    g116(.A(new_n282), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(KEYINPUT33), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n308), .A3(new_n315), .A4(new_n313), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(new_n300), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n300), .B1(new_n322), .B2(new_n323), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n301), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327));
  INV_X1    g126(.A(G64gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G92gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(G197gat), .ZN(new_n334));
  INV_X1    g133(.A(G204gat), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n335), .A2(KEYINPUT79), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(KEYINPUT79), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT79), .B(G204gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G197gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT80), .B(G211gat), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT22), .B1(new_n342), .B2(G218gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT81), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n338), .A4(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(G211gat), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n344), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n333), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n344), .A2(new_n349), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G211gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(G218gat), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n293), .A2(KEYINPUT82), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n288), .A2(new_n361), .A3(new_n292), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(KEYINPUT29), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n293), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n359), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n360), .A2(new_n362), .A3(new_n366), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n265), .A2(new_n364), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n359), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n332), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n363), .A2(new_n364), .B1(new_n293), .B2(new_n366), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n371), .B(new_n331), .C1(new_n374), .C2(new_n359), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(new_n332), .C1(new_n368), .C2(new_n372), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  XOR2_X1   g179(.A(G155gat), .B(G162gat), .Z(new_n381));
  XNOR2_X1  g180(.A(G141gat), .B(G148gat), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(KEYINPUT84), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G155gat), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT2), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n386), .C1(KEYINPUT84), .C2(new_n382), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n381), .A2(KEYINPUT83), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(KEYINPUT83), .ZN(new_n389));
  INV_X1    g188(.A(new_n386), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n294), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n387), .A2(new_n391), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n280), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n397), .B2(new_n280), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n380), .B(new_n396), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT5), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT85), .B1(new_n397), .B2(new_n280), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n397), .B2(new_n280), .ZN(new_n406));
  INV_X1    g205(.A(new_n380), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n294), .A2(KEYINPUT85), .A3(new_n392), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n397), .A2(new_n280), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT4), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n399), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n412), .A2(KEYINPUT5), .A3(new_n380), .A4(new_n396), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n404), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G57gat), .ZN(new_n417));
  INV_X1    g216(.A(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n404), .A2(new_n413), .A3(new_n422), .A4(new_n409), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  OR3_X1    g223(.A1(new_n414), .A2(new_n421), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n379), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT33), .B1(new_n317), .B2(new_n318), .ZN(new_n429));
  INV_X1    g228(.A(new_n313), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n319), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT32), .B(new_n320), .C1(new_n305), .C2(new_n282), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n323), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT77), .A3(new_n300), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n395), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n358), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G228gat), .ZN(new_n440));
  INV_X1    g239(.A(G233gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n353), .A2(new_n357), .A3(new_n437), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n353), .A2(new_n357), .A3(KEYINPUT86), .A4(new_n437), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n394), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n449), .B2(new_n392), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n358), .A2(new_n438), .B1(KEYINPUT3), .B2(new_n392), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n353), .A2(new_n357), .A3(new_n437), .A4(new_n392), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n443), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n436), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n452), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n442), .ZN(new_n456));
  INV_X1    g255(.A(new_n436), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT3), .B1(new_n445), .B2(new_n446), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n397), .B1(new_n458), .B2(new_n448), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n456), .B(new_n457), .C1(new_n459), .C2(new_n444), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(G22gat), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(new_n460), .A3(new_n463), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n326), .A2(new_n428), .A3(new_n435), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT35), .ZN(new_n469));
  INV_X1    g268(.A(new_n300), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n434), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n379), .A2(new_n426), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n322), .A2(new_n300), .A3(new_n323), .ZN(new_n474));
  AND4_X1   g273(.A1(new_n471), .A2(new_n473), .A3(new_n467), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT35), .B1(new_n427), .B2(KEYINPUT88), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n301), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n471), .B2(new_n474), .ZN(new_n480));
  INV_X1    g279(.A(new_n435), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT36), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT36), .ZN(new_n483));
  INV_X1    g282(.A(new_n467), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n427), .ZN(new_n485));
  INV_X1    g284(.A(new_n379), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n380), .B1(new_n412), .B2(new_n396), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n412), .A2(new_n396), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n490), .A3(new_n407), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n419), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT87), .B(new_n487), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n423), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n407), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n406), .A2(new_n408), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n380), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT39), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n419), .A3(new_n493), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT87), .B1(new_n501), .B2(new_n487), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n501), .A2(new_n487), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n426), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n368), .B2(new_n372), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n331), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n368), .A2(new_n372), .A3(new_n507), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n374), .B2(new_n359), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n369), .A2(new_n370), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n359), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n331), .A4(new_n508), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n506), .A2(new_n511), .A3(new_n373), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n505), .A2(new_n517), .A3(new_n467), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n482), .A2(new_n483), .A3(new_n485), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n478), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(KEYINPUT8), .A2(new_n523), .B1(new_n418), .B2(new_n330), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G99gat), .B(G106gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n529), .B1(new_n533), .B2(KEYINPUT89), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NOR2_X1   g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n530), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n528), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(new_n529), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n543), .A2(new_n540), .A3(new_n528), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT96), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n527), .B(KEYINPUT95), .Z(new_n551));
  AOI21_X1  g350(.A(KEYINPUT90), .B1(new_n542), .B2(new_n545), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555));
  AOI22_X1  g354(.A1(new_n550), .A2(new_n554), .B1(KEYINPUT97), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(KEYINPUT97), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n558), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n565), .A2(KEYINPUT98), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n559), .A2(new_n567), .A3(new_n560), .A4(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n559), .A2(new_n560), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT99), .B1(new_n570), .B2(new_n563), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT99), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n572), .B(new_n564), .C1(new_n559), .C2(new_n560), .ZN(new_n573));
  OAI22_X1  g372(.A1(new_n566), .A2(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  XOR2_X1   g374(.A(G15gat), .B(G22gat), .Z(new_n576));
  INV_X1    g375(.A(G1gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(KEYINPUT16), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT91), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n575), .B(new_n578), .C1(new_n580), .C2(new_n576), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(G8gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(G8gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT21), .ZN(new_n586));
  INV_X1    g385(.A(G57gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n328), .A2(G57gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(KEYINPUT9), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT93), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n592), .B(new_n594), .C1(G71gat), .C2(G78gat), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n588), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n593), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n585), .B1(new_n586), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n586), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G127gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(G155gat), .B(G183gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n608), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n350), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n574), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n520), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n584), .A2(new_n546), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n585), .B2(new_n553), .ZN(new_n620));
  NAND2_X1  g419(.A1(G229gat), .A2(G233gat), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(KEYINPUT18), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n584), .B(new_n546), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n621), .B(KEYINPUT13), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(KEYINPUT18), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT11), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n247), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n623), .A2(new_n634), .A3(new_n627), .A4(new_n628), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n527), .B(new_n604), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n642), .B2(KEYINPUT10), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n527), .A2(KEYINPUT10), .A3(new_n603), .A4(new_n595), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(KEYINPUT100), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n648), .B2(new_n641), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n248), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n335), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n650), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n618), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n506), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n486), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  AND2_X1   g459(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n659), .A2(G8gat), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT42), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(KEYINPUT42), .B2(new_n662), .ZN(G1325gat));
  NOR2_X1   g464(.A1(new_n324), .A2(new_n325), .ZN(new_n666));
  AOI21_X1  g465(.A(G15gat), .B1(new_n656), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n482), .A2(new_n483), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n656), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n656), .A2(new_n484), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n574), .A2(KEYINPUT102), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n570), .A2(new_n563), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n572), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n570), .A2(KEYINPUT99), .A3(new_n563), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n565), .A2(KEYINPUT98), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n568), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n676), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n520), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n678), .A2(new_n679), .B1(new_n681), .B2(new_n568), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n478), .B2(new_n519), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT101), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AND4_X1   g489(.A1(new_n482), .A2(new_n483), .A3(new_n485), .A4(new_n518), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n468), .A2(KEYINPUT35), .B1(new_n475), .B2(new_n476), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n574), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT44), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n686), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n655), .A2(new_n616), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n674), .B1(new_n699), .B2(new_n426), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(KEYINPUT103), .A3(new_n506), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(G29gat), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n693), .A2(new_n697), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n531), .A3(new_n506), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1328gat));
  OAI21_X1  g505(.A(G36gat), .B1(new_n699), .B2(new_n379), .ZN(new_n707));
  NAND2_X1  g506(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n703), .A2(new_n532), .A3(new_n486), .A4(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(new_n668), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n696), .A2(new_n713), .A3(new_n697), .ZN(new_n714));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT105), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n703), .A2(new_n715), .A3(new_n666), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI221_X1 g519(.A(new_n717), .B1(KEYINPUT105), .B2(KEYINPUT47), .C1(new_n714), .C2(new_n715), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n696), .A2(new_n467), .A3(new_n697), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n703), .A2(new_n725), .A3(new_n484), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n728), .A3(KEYINPUT48), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  OAI221_X1 g529(.A(new_n727), .B1(new_n723), .B2(new_n730), .C1(new_n724), .C2(new_n725), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(G1331gat));
  INV_X1    g531(.A(new_n654), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n638), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n618), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n426), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n587), .ZN(G1332gat));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n379), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g541(.A(new_n735), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(G71gat), .A3(new_n668), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(KEYINPUT107), .A3(new_n666), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  INV_X1    g545(.A(new_n666), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n735), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n744), .B1(new_n749), .B2(G71gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT50), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n752), .B(new_n744), .C1(new_n749), .C2(G71gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n735), .A2(new_n467), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n600), .ZN(G1335gat));
  INV_X1    g555(.A(new_n686), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n688), .A2(KEYINPUT101), .A3(new_n689), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n694), .B1(new_n693), .B2(KEYINPUT44), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n638), .A2(new_n615), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n654), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n426), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n574), .B(new_n761), .C1(new_n691), .C2(new_n692), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n520), .A2(new_n574), .A3(new_n761), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n418), .B(new_n506), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n763), .B1(new_n733), .B2(new_n775), .ZN(G1336gat));
  OAI21_X1  g575(.A(G92gat), .B1(new_n762), .B2(new_n379), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n486), .A2(new_n330), .A3(new_n654), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT110), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n777), .A2(new_n783), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n762), .B2(new_n713), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n773), .A2(new_n774), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n666), .A2(new_n312), .A3(new_n654), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT112), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(G1338gat));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n760), .A2(new_n654), .A3(new_n484), .A4(new_n761), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n795));
  INV_X1    g594(.A(G106gat), .ZN(new_n796));
  AND4_X1   g595(.A1(new_n796), .A2(new_n772), .A3(new_n654), .A4(new_n484), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AND4_X1   g597(.A1(new_n792), .A2(new_n794), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n793), .B2(G106gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n792), .B1(new_n800), .B2(new_n795), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(G1339gat));
  OR3_X1    g601(.A1(new_n620), .A2(KEYINPUT115), .A3(new_n621), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n625), .A2(new_n626), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT115), .B1(new_n620), .B2(new_n621), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n633), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n637), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n654), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  INV_X1    g609(.A(new_n648), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n643), .A2(new_n811), .A3(new_n644), .A4(new_n646), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n649), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n653), .B1(new_n649), .B2(KEYINPUT54), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n650), .A2(new_n653), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n649), .A2(KEYINPUT54), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n813), .A4(new_n653), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n809), .B1(new_n639), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n574), .A2(KEYINPUT102), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n680), .A2(new_n676), .A3(new_n682), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n819), .A2(new_n817), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n816), .A3(new_n808), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n822), .B2(new_n823), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n616), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n617), .A2(new_n829), .A3(new_n733), .A4(new_n639), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n687), .A2(new_n733), .A3(new_n639), .A4(new_n615), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT114), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n426), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n747), .A2(new_n484), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n379), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n639), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n326), .A2(new_n435), .A3(new_n467), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n826), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n675), .B2(new_n683), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n615), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n832), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n506), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT116), .B1(new_n847), .B2(new_n839), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n841), .A2(new_n848), .A3(new_n379), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n638), .A2(new_n268), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n837), .B1(new_n850), .B2(new_n851), .ZN(G1340gat));
  OAI21_X1  g651(.A(G120gat), .B1(new_n836), .B2(new_n733), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n654), .A2(new_n266), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n850), .B2(new_n854), .ZN(G1341gat));
  XNOR2_X1  g654(.A(KEYINPUT73), .B(G127gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n836), .B2(new_n616), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n850), .A2(new_n856), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n616), .ZN(G1342gat));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n849), .A2(new_n860), .A3(new_n274), .A4(new_n574), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n836), .B2(new_n687), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n841), .A2(new_n848), .A3(new_n274), .A4(new_n379), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT56), .B1(new_n863), .B2(new_n687), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT117), .ZN(G1343gat));
  AOI21_X1  g665(.A(new_n467), .B1(new_n828), .B2(new_n833), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n668), .A2(new_n426), .A3(new_n486), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(G141gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n638), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n816), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n816), .A2(new_n873), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n638), .B(new_n825), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n574), .B1(new_n876), .B2(new_n809), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n827), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n846), .B1(new_n880), .B2(new_n616), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n467), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n884), .A3(new_n868), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n639), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n886), .B2(new_n871), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n872), .C1(new_n886), .C2(new_n871), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n892), .A3(new_n654), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n826), .A2(new_n687), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n616), .B1(new_n877), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n467), .B1(new_n899), .B2(new_n831), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT57), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n654), .A3(new_n868), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n894), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  INV_X1    g706(.A(new_n885), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT59), .B(new_n892), .C1(new_n908), .C2(new_n654), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n893), .B1(new_n907), .B2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n885), .B2(new_n616), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n870), .A2(new_n384), .A3(new_n615), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n870), .B2(new_n574), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n684), .A2(new_n385), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n908), .B2(new_n915), .ZN(G1347gat));
  OAI21_X1  g715(.A(new_n426), .B1(new_n845), .B2(new_n846), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n379), .A3(new_n839), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT122), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n638), .A3(new_n258), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n506), .B1(new_n828), .B2(new_n833), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n486), .A3(new_n835), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n639), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(G1348gat));
  NOR3_X1   g723(.A1(new_n922), .A2(new_n248), .A3(new_n733), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT123), .Z(new_n926));
  AOI21_X1  g725(.A(G176gat), .B1(new_n919), .B2(new_n654), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1349gat));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n921), .A2(new_n228), .A3(new_n486), .A4(new_n840), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n616), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n918), .A2(KEYINPUT124), .A3(new_n228), .A4(new_n615), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  OAI21_X1  g733(.A(G183gat), .B1(new_n922), .B2(new_n616), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n228), .ZN(new_n940));
  NOR4_X1   g739(.A1(new_n917), .A2(new_n940), .A3(new_n379), .A4(new_n839), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT124), .B1(new_n941), .B2(new_n615), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n930), .A2(new_n929), .A3(new_n616), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n935), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT60), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n939), .A2(new_n947), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n922), .B2(new_n687), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  INV_X1    g749(.A(new_n684), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n919), .A2(new_n219), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1351gat));
  NOR2_X1   g752(.A1(new_n506), .A2(new_n379), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n713), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n905), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n639), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n867), .A2(new_n956), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n334), .A3(new_n638), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n335), .A3(new_n654), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  AOI211_X1 g762(.A(new_n733), .B(new_n955), .C1(new_n897), .C2(new_n904), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n335), .ZN(G1353gat));
  AOI211_X1 g764(.A(new_n616), .B(new_n955), .C1(new_n897), .C2(new_n904), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT63), .B1(new_n966), .B2(new_n350), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n968), .B(G211gat), .C1(new_n957), .C2(new_n616), .ZN(new_n969));
  INV_X1    g768(.A(new_n342), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n970), .A3(new_n615), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n967), .A2(new_n969), .A3(new_n972), .ZN(G1354gat));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n333), .A3(new_n687), .ZN(new_n974));
  AOI21_X1  g773(.A(G218gat), .B1(new_n959), .B2(new_n951), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT127), .Z(new_n976));
  NOR2_X1   g775(.A1(new_n974), .A2(new_n976), .ZN(G1355gat));
endmodule


