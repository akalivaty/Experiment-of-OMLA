//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT66), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n464), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n473), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OR2_X1    g058(.A1(new_n462), .A2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n469), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n473), .A2(new_n488), .A3(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n478), .B2(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  OR2_X1    g071(.A1(KEYINPUT67), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT67), .A2(G651), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(KEYINPUT6), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n503), .A3(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  AND3_X1   g083(.A1(new_n508), .A2(KEYINPUT69), .A3(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT69), .B1(new_n508), .B2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n505), .A2(new_n506), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n508), .A2(KEYINPUT69), .A3(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n518), .A2(new_n519), .B1(KEYINPUT5), .B2(new_n506), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n497), .A2(new_n498), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(G51), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n499), .A2(new_n504), .A3(G543), .A4(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(KEYINPUT71), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT71), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n531));
  AND3_X1   g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT73), .B(G89), .Z(new_n534));
  NAND4_X1  g109(.A1(new_n520), .A2(new_n499), .A3(new_n504), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n523), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n520), .A2(G90), .A3(new_n499), .A4(new_n504), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n499), .A2(new_n504), .A3(G52), .A4(G543), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n523), .B1(new_n547), .B2(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(G81), .A2(new_n512), .B1(new_n514), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT76), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT77), .Z(G188));
  NAND4_X1  g137(.A1(new_n499), .A2(new_n504), .A3(G53), .A4(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G651), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n568), .B1(new_n505), .B2(new_n511), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n520), .A2(KEYINPUT78), .A3(new_n499), .A4(new_n504), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(G91), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n564), .A2(new_n567), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(G168), .ZN(G286));
  OR2_X1    g148(.A1(new_n516), .A2(new_n524), .ZN(G303));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n566), .B1(new_n511), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(G49), .B2(new_n514), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n569), .A2(G87), .A3(new_n570), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n569), .A2(G86), .A3(new_n570), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n511), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n522), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n499), .A2(new_n504), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n587), .A2(G48), .A3(G543), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n582), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n511), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT80), .B(new_n591), .C1(new_n511), .C2(new_n592), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n595), .A2(new_n596), .A3(new_n522), .ZN(new_n597));
  AOI22_X1  g172(.A1(G85), .A2(new_n512), .B1(new_n514), .B2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  NAND3_X1  g174(.A1(new_n569), .A2(G92), .A3(new_n570), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n569), .A2(KEYINPUT10), .A3(G92), .A4(new_n570), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n499), .A2(new_n504), .A3(G54), .A4(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(G66), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n604), .B(new_n605), .C1(new_n608), .C2(new_n566), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n566), .B1(new_n606), .B2(new_n607), .ZN(new_n610));
  INV_X1    g185(.A(new_n605), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT81), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n602), .A2(new_n603), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n613), .A2(KEYINPUT82), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(KEYINPUT82), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(G301), .B(new_n616), .S(new_n617), .Z(G284));
  MUX2_X1   g193(.A(G301), .B(new_n616), .S(new_n617), .Z(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n617), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n617), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(new_n616), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  OAI21_X1  g200(.A(new_n624), .B1(new_n614), .B2(new_n615), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n471), .A2(new_n484), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n478), .A2(G123), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n473), .A2(G135), .ZN(new_n638));
  NOR3_X1   g213(.A1(new_n469), .A2(KEYINPUT85), .A3(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT85), .B1(new_n469), .B2(G111), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(G2104), .A3(new_n641), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT86), .B(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n634), .A2(new_n635), .A3(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n677), .A2(new_n680), .A3(new_n684), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(KEYINPUT99), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n696), .A2(G32), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n471), .A2(G105), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT97), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n473), .A2(G141), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n478), .A2(G129), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n697), .B1(new_n707), .B2(G29), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G11), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT30), .B(G28), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(new_n696), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n711), .B(new_n713), .C1(new_n643), .C2(new_n696), .ZN(new_n714));
  INV_X1    g289(.A(G2084), .ZN(new_n715));
  AND2_X1   g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NOR2_X1   g291(.A1(KEYINPUT24), .A2(G34), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n696), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT95), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n475), .B2(new_n696), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n714), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n696), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n473), .A2(G140), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n478), .A2(G128), .ZN(new_n725));
  OR2_X1    g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(new_n696), .ZN(new_n729));
  INV_X1    g304(.A(G2067), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n708), .A2(new_n709), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n710), .A2(new_n721), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n696), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n696), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT98), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT98), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n736), .A2(G2078), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(G2078), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G20), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT23), .ZN(new_n743));
  INV_X1    g318(.A(G299), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n741), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n720), .A2(new_n715), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n696), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n696), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G2090), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n741), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n555), .B2(new_n741), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT91), .B(G1341), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT92), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n752), .A2(G2090), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n749), .A2(new_n753), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n740), .A2(new_n747), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n696), .A2(G33), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT25), .Z(new_n765));
  INV_X1    g340(.A(G139), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n485), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT93), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n484), .A2(G127), .ZN(new_n769));
  AND2_X1   g344(.A1(G115), .A2(G2104), .ZN(new_n770));
  OAI21_X1  g345(.A(G2105), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n763), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(G171), .A2(new_n741), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G5), .B2(new_n741), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n775), .A2(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n772), .B(KEYINPUT94), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n762), .B1(new_n782), .B2(new_n696), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n781), .B1(new_n783), .B2(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n741), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n741), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(G1966), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n755), .A2(new_n757), .B1(G1966), .B2(new_n786), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n780), .A2(new_n784), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n761), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G4), .A2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT90), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n616), .B2(new_n741), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n696), .A2(G25), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n473), .A2(G131), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n478), .A2(G119), .ZN(new_n797));
  OR2_X1    g372(.A1(G95), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(new_n696), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  AND2_X1   g379(.A1(new_n741), .A2(G24), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G290), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1986), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n741), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n741), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1971), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n741), .A2(G23), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G288), .B2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT33), .B(G1976), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n816), .A2(new_n818), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n741), .A2(G6), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n582), .A2(new_n589), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n741), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT32), .B(G1981), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n821), .A2(new_n826), .A3(KEYINPUT34), .A4(new_n827), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n811), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT89), .B(KEYINPUT36), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n790), .B(new_n794), .C1(new_n832), .C2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(KEYINPUT89), .A3(KEYINPUT36), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n695), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n790), .A2(new_n794), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n832), .A2(new_n834), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT99), .A4(new_n836), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n838), .A2(new_n841), .ZN(G311));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n840), .A3(new_n836), .ZN(G150));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n523), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT100), .B(G93), .Z(new_n848));
  NAND3_X1  g423(.A1(new_n587), .A2(new_n520), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n499), .A2(new_n504), .A3(G55), .A4(G543), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n849), .A2(KEYINPUT101), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT101), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT102), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(new_n847), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n554), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n853), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n555), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n623), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n845), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n844), .B1(new_n845), .B2(new_n863), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n853), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n800), .B(KEYINPUT106), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n478), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n469), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(G142), .B2(new_n473), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(new_n632), .Z(new_n879));
  NAND3_X1  g454(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n706), .B(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(new_n495), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n495), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n782), .A2(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n782), .A2(KEYINPUT105), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n882), .A2(KEYINPUT105), .A3(new_n782), .A4(new_n883), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n475), .B(new_n482), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n643), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n887), .A2(new_n879), .A3(new_n893), .A4(new_n888), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(new_n879), .A3(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT107), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n891), .B1(new_n898), .B2(new_n889), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n903));
  AND2_X1   g478(.A1(G290), .A2(G288), .ZN(new_n904));
  NOR2_X1   g479(.A1(G290), .A2(G288), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G166), .B1(new_n582), .B2(new_n589), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G288), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n597), .A3(new_n598), .ZN(new_n910));
  NAND2_X1  g485(.A1(G290), .A2(G288), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT111), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n582), .A2(G166), .A3(new_n589), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n906), .A2(new_n908), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n904), .A2(new_n905), .ZN(new_n915));
  INV_X1    g490(.A(new_n913), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n915), .B(KEYINPUT111), .C1(new_n916), .C2(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n626), .B(new_n860), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n602), .A2(new_n603), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n609), .A2(new_n612), .ZN(new_n923));
  AND4_X1   g498(.A1(KEYINPUT108), .A2(new_n922), .A3(G299), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT108), .B1(new_n613), .B2(G299), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(G299), .A3(new_n923), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n613), .A2(KEYINPUT108), .A3(G299), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n613), .A2(G299), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n920), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n613), .A2(G299), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n929), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT110), .B1(new_n937), .B2(KEYINPUT41), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n933), .B1(new_n924), .B2(new_n925), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n936), .A2(new_n941), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n938), .A2(new_n942), .B1(new_n932), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n935), .B1(new_n920), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT112), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n935), .B(new_n947), .C1(new_n920), .C2(new_n944), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n919), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n919), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n858), .ZN(G331));
  XNOR2_X1  g528(.A(G301), .B(G168), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n857), .A2(new_n859), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n857), .B2(new_n859), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n938), .A2(new_n942), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n932), .A2(new_n943), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n954), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n860), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n857), .A2(new_n954), .A3(new_n859), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n936), .B1(new_n926), .B2(new_n931), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n917), .B(new_n914), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT113), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n918), .B1(new_n934), .B2(new_n957), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n968), .B(new_n969), .C1(new_n944), .C2(new_n957), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n934), .A2(new_n957), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n943), .B1(new_n925), .B2(new_n924), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n943), .B(KEYINPUT114), .C1(new_n925), .C2(new_n924), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n964), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n972), .B(new_n977), .C1(KEYINPUT41), .C2(new_n965), .ZN(new_n978));
  AOI21_X1  g553(.A(G37), .B1(new_n978), .B2(new_n918), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n972), .B1(new_n944), .B2(new_n957), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n918), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT43), .B1(new_n971), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT44), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n971), .A2(new_n986), .A3(new_n979), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n971), .B2(new_n982), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  NAND2_X1  g565(.A1(new_n728), .A2(new_n730), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n880), .A2(G2067), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT116), .Z(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n706), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n495), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G40), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n475), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n995), .A2(new_n997), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n996), .A3(new_n706), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n801), .A2(new_n803), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n801), .A2(new_n803), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1005), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n490), .B2(new_n494), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1003), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n823), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n512), .A2(G86), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n588), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(KEYINPUT118), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1021), .A2(KEYINPUT118), .B1(new_n522), .B2(new_n585), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1017), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1024), .B1(new_n823), .B2(new_n1018), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1029), .A2(KEYINPUT119), .A3(KEYINPUT49), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT119), .B1(new_n1029), .B2(KEYINPUT49), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1017), .B1(G1976), .B2(new_n909), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(new_n1033), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1971), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1015), .A2(KEYINPUT45), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1000), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1003), .B1(new_n1015), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1015), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT117), .B(G2090), .Z(new_n1049));
  NAND4_X1  g624(.A1(new_n1046), .A2(new_n1003), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(G166), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1051), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1051), .B2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1032), .A2(new_n1039), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT126), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1029), .A2(KEYINPUT119), .A3(KEYINPUT49), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1038), .B1(new_n1066), .B2(new_n1028), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT126), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1059), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(G301), .B(KEYINPUT54), .Z(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1001), .A2(new_n1003), .A3(new_n1041), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(G2078), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1046), .A2(new_n1003), .A3(new_n1048), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(G1961), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1072), .A2(G2078), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1001), .A2(new_n1003), .A3(new_n1041), .A4(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT125), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1071), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n999), .A2(new_n1000), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1003), .B1(new_n1015), .B2(KEYINPUT45), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1083), .A2(new_n1072), .A3(G2078), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1076), .A2(new_n1084), .A3(new_n1071), .ZN(new_n1085));
  INV_X1    g660(.A(G1966), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1046), .A2(new_n1003), .A3(new_n1048), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT121), .B(G2084), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1087), .B(G168), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1092), .A2(KEYINPUT51), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1075), .A2(new_n1089), .ZN(new_n1094));
  AOI21_X1  g669(.A(G168), .B1(new_n1094), .B2(new_n1087), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1080), .A2(new_n1085), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1075), .A2(G1348), .B1(G2067), .B2(new_n1016), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n616), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1016), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1088), .A2(new_n1101), .B1(new_n730), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n623), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(G299), .B(KEYINPUT57), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1088), .A2(new_n746), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1001), .A2(new_n1003), .A3(new_n1041), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1112));
  OR3_X1    g687(.A1(new_n1111), .A2(new_n1112), .A3(KEYINPUT61), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1111), .B2(KEYINPUT61), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n554), .A2(KEYINPUT124), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1001), .A2(new_n996), .A3(new_n1003), .A4(new_n1041), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1016), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  AND4_X1   g696(.A1(new_n1106), .A2(new_n1113), .A3(new_n1114), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1107), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1124), .B2(new_n1123), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1098), .A2(new_n623), .A3(KEYINPUT122), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1103), .B2(new_n616), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1123), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1126), .A2(new_n1130), .B1(new_n1107), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1097), .B1(new_n1122), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1093), .A2(new_n1096), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1135), .A2(G171), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1070), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1017), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1029), .B2(KEYINPUT49), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n909), .A2(new_n1034), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1019), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT120), .B(new_n1019), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1141), .A3(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1054), .B(G286), .C1(new_n1094), .C2(new_n1087), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1032), .A2(new_n1039), .A3(new_n1059), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1067), .A2(KEYINPUT63), .A3(new_n1059), .A4(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1067), .A2(new_n1057), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1149), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1014), .B1(new_n1140), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1005), .A2(new_n996), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT46), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n995), .A2(new_n1005), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n991), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1005), .ZN(new_n1166));
  NOR4_X1   g741(.A1(new_n1001), .A2(G1986), .A3(G290), .A4(new_n1004), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT48), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1012), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT127), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1158), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(G227), .A2(new_n460), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n662), .A2(new_n693), .A3(new_n1174), .ZN(new_n1175));
  OAI211_X1 g749(.A(new_n901), .B(new_n1175), .C1(new_n987), .C2(new_n988), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


