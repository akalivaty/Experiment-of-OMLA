//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n219), .A2(new_n220), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  INV_X1    g0033(.A(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n225), .B1(new_n206), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n253), .B2(G20), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(new_n255), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT75), .ZN(new_n261));
  INV_X1    g0061(.A(G58), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n264), .B2(new_n201), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G159), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G33), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(G20), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT74), .B1(new_n275), .B2(KEYINPUT7), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT74), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n273), .B1(new_n281), .B2(G33), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n277), .B(new_n278), .C1(new_n282), .C2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n275), .A2(KEYINPUT7), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n276), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n268), .B1(new_n285), .B2(G68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT16), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n278), .B1(new_n288), .B2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n257), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n226), .A2(KEYINPUT7), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n268), .B1(new_n294), .B2(G68), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n258), .B1(new_n295), .B2(KEYINPUT16), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n261), .B1(new_n287), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT17), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G223), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n234), .B2(new_n300), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n271), .A2(new_n302), .A3(new_n274), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G41), .A2(G45), .ZN(new_n308));
  INV_X1    g0108(.A(G274), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n308), .A2(G1), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n308), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n306), .B1(new_n253), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n312), .B2(G232), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G190), .B2(new_n314), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n298), .A2(new_n299), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT76), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n298), .A2(new_n319), .A3(new_n317), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n260), .B(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n323), .B(new_n268), .C1(new_n285), .C2(G68), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n317), .B(new_n322), .C1(new_n324), .C2(new_n296), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n318), .B1(new_n327), .B2(new_n299), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n314), .A2(G179), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n314), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n296), .B1(new_n286), .B2(KEYINPUT16), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n261), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n333), .B(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT77), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n288), .A2(new_n300), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n234), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n306), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n310), .B1(new_n312), .B2(G238), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n330), .A2(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n343), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n344), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n349), .B(new_n351), .C1(new_n352), .C2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n254), .A2(G68), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n263), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n257), .A2(G20), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n258), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT11), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n366), .B1(new_n259), .B2(G68), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n366), .B2(new_n365), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n357), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n346), .A2(G200), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n369), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n356), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n288), .A2(G223), .A3(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G222), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n379), .B1(new_n363), .B2(new_n288), .C1(new_n339), .C2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(KEYINPUT68), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(KEYINPUT68), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n306), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n310), .B1(new_n312), .B2(G226), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G200), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(G190), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n254), .A2(G50), .ZN(new_n391));
  INV_X1    g0191(.A(new_n258), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n255), .A2(new_n362), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n391), .B(new_n396), .C1(G50), .C2(new_n259), .ZN(new_n397));
  XOR2_X1   g0197(.A(new_n397), .B(KEYINPUT9), .Z(new_n398));
  NAND4_X1  g0198(.A1(new_n390), .A2(KEYINPUT69), .A3(KEYINPUT10), .A4(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n387), .B2(new_n389), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT69), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n402), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n386), .A2(G179), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n388), .A2(G169), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n397), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n288), .A2(G238), .A3(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n288), .A2(G232), .A3(new_n300), .ZN(new_n411));
  INV_X1    g0211(.A(G107), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n288), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n306), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n310), .B1(new_n312), .B2(G244), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G169), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n352), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n259), .A2(G77), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G77), .B2(new_n254), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n255), .A2(G20), .A3(G33), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT15), .B(G87), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n361), .B1(G20), .B2(G77), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n392), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n416), .A2(new_n315), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G190), .B2(new_n416), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n427), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n409), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n399), .A2(new_n406), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(KEYINPUT70), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(KEYINPUT70), .ZN(new_n437));
  AOI211_X1 g0237(.A(new_n336), .B(new_n378), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n328), .A2(new_n335), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT77), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n282), .A2(G244), .A3(new_n300), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT4), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n300), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n306), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n253), .A2(G45), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT78), .B1(new_n454), .B2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT78), .ZN(new_n456));
  INV_X1    g0256(.A(G41), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT5), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n455), .B(new_n458), .C1(KEYINPUT5), .C2(new_n457), .ZN(new_n459));
  NOR4_X1   g0259(.A1(new_n453), .A2(new_n459), .A3(new_n309), .A4(new_n306), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n453), .A2(new_n459), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n306), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(G257), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n452), .B2(new_n463), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n330), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n464), .A2(G179), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n294), .A2(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n412), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  XOR2_X1   g0272(.A(G97), .B(G107), .Z(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(KEYINPUT6), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n392), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n254), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n210), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n258), .B1(new_n253), .B2(G33), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n254), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(new_n210), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n468), .A2(new_n470), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n482), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n464), .B2(G200), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n488));
  INV_X1    g0288(.A(new_n460), .ZN(new_n489));
  INV_X1    g0289(.A(new_n306), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(new_n490), .C1(new_n453), .C2(new_n459), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n446), .B2(new_n450), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n466), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n487), .B1(new_n496), .B2(new_n374), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n490), .B1(new_n453), .B2(G274), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n209), .B2(new_n453), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n282), .A2(G244), .A3(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n282), .A2(new_n502), .A3(G244), .A4(G1698), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n257), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n282), .A2(G238), .A3(new_n300), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n501), .A2(new_n503), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n499), .B1(new_n508), .B2(new_n306), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n352), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n480), .A2(new_n423), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n338), .B2(G20), .ZN(new_n513));
  XOR2_X1   g0313(.A(new_n513), .B(KEYINPUT82), .Z(new_n514));
  NAND3_X1  g0314(.A1(new_n282), .A2(new_n226), .A3(G68), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n226), .B1(new_n338), .B2(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n208), .A2(new_n210), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(G107), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n519), .A2(new_n392), .B1(new_n254), .B2(new_n424), .ZN(new_n520));
  OAI221_X1 g0320(.A(new_n510), .B1(G169), .B2(new_n509), .C1(new_n511), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n509), .A2(G190), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n480), .A2(new_n208), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n524), .C1(new_n315), .C2(new_n509), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n485), .A2(new_n497), .A3(new_n521), .A4(new_n525), .ZN(new_n526));
  MUX2_X1   g0326(.A(new_n254), .B(new_n480), .S(G116), .Z(new_n527));
  NAND2_X1  g0327(.A1(new_n257), .A2(G97), .ZN(new_n528));
  AOI21_X1  g0328(.A(G20), .B1(new_n528), .B2(new_n449), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n226), .A2(new_n504), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n258), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g0331(.A(new_n531), .B(KEYINPUT20), .Z(new_n532));
  AND2_X1   g0332(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G264), .A2(G1698), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n211), .B2(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n282), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G303), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n288), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n306), .ZN(new_n539));
  OAI211_X1 g0339(.A(G270), .B(new_n490), .C1(new_n453), .C2(new_n459), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n489), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n533), .B1(new_n542), .B2(new_n315), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT83), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n533), .B(new_n545), .C1(new_n542), .C2(new_n315), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(G190), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(G169), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n352), .B2(new_n541), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n527), .A2(new_n532), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n460), .B1(new_n538), .B2(new_n306), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n330), .B1(new_n553), .B2(new_n540), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n552), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n551), .A2(new_n552), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n462), .A2(G264), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G257), .A2(G1698), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n209), .B2(G1698), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n282), .A2(new_n559), .B1(G33), .B2(G294), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n489), .C1(new_n490), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n315), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G190), .B2(new_n561), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  AOI22_X1  g0364(.A1(KEYINPUT85), .A2(new_n564), .B1(new_n412), .B2(G20), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(KEYINPUT85), .B2(new_n564), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n565), .B(KEYINPUT86), .C1(KEYINPUT85), .C2(new_n564), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n226), .A2(KEYINPUT23), .A3(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n226), .B2(new_n505), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n282), .A2(new_n226), .A3(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  XNOR2_X1  g0374(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n288), .A2(new_n575), .A3(new_n226), .A4(G87), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n392), .B1(new_n577), .B2(KEYINPUT24), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(KEYINPUT24), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n480), .A2(new_n412), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n477), .B2(new_n412), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n254), .A2(KEYINPUT25), .A3(G107), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n563), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n557), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n560), .A2(new_n490), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(G179), .A3(new_n489), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n561), .A2(G169), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n579), .A2(new_n584), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n548), .A2(new_n556), .A3(new_n585), .A4(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n443), .A2(new_n526), .A3(new_n594), .ZN(G372));
  OAI21_X1  g0395(.A(new_n371), .B1(new_n376), .B2(new_n429), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n328), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n333), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n334), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n333), .B(KEYINPUT87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT18), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT88), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n399), .A2(new_n406), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n399), .B2(new_n406), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n409), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n555), .A2(new_n550), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n541), .A2(new_n352), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(KEYINPUT21), .B2(new_n554), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n612), .B2(new_n533), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n589), .A2(new_n590), .B1(new_n579), .B2(new_n584), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n585), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n521), .B1(new_n526), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(G169), .B1(new_n488), .B2(new_n495), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n617), .A2(new_n469), .A3(new_n482), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n521), .A4(new_n525), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n521), .A2(new_n525), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT26), .B1(new_n621), .B2(new_n485), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n609), .B1(new_n443), .B2(new_n624), .ZN(G369));
  AND2_X1   g0425(.A1(new_n226), .A2(G13), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n253), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G213), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G343), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n592), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n585), .A2(new_n593), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT90), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n585), .A2(new_n593), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n632), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n635), .B(new_n637), .C1(new_n593), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n552), .A2(new_n632), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n548), .A2(new_n556), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n613), .A2(new_n552), .A3(new_n632), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n641), .B2(new_n642), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n639), .B(G330), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT91), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n642), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n644), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT91), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(G330), .A4(new_n639), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n556), .A2(new_n632), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n635), .B2(new_n637), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n593), .A2(new_n632), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n221), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n517), .A2(G107), .A3(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n228), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT92), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT30), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n611), .A2(new_n509), .A3(new_n588), .A4(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n465), .A2(new_n467), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n670), .A3(new_n674), .A4(KEYINPUT30), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(KEYINPUT30), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n496), .B2(new_n672), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n561), .A2(new_n541), .A3(new_n352), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n678), .A2(new_n509), .A3(new_n494), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT31), .B1(new_n680), .B2(new_n632), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT93), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n526), .A2(new_n594), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n638), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n632), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n669), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n638), .B1(new_n616), .B2(new_n623), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n621), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .A3(new_n618), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n619), .B1(new_n621), .B2(new_n485), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(KEYINPUT94), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(KEYINPUT94), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT29), .B(new_n638), .C1(new_n697), .C2(new_n616), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n688), .B1(new_n691), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n668), .B1(new_n699), .B2(G1), .ZN(G364));
  NAND2_X1  g0500(.A1(new_n626), .A2(G45), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n664), .A2(G1), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n651), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n669), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n651), .A2(G330), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(G13), .A2(G33), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n374), .A2(G20), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G179), .A2(G200), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G159), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT32), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n315), .A2(G179), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n712), .A2(new_n352), .A3(G200), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n721), .A2(G107), .B1(G77), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n352), .A2(new_n315), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n226), .A2(new_n374), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n718), .B(new_n723), .C1(new_n202), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n719), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G87), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n352), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n262), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n226), .B1(new_n714), .B2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n210), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n713), .A2(new_n724), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n288), .B1(new_n737), .B2(new_n263), .ZN(new_n738));
  OR3_X1    g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n730), .A2(G303), .B1(new_n726), .B2(G326), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  INV_X1    g0541(.A(new_n722), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT33), .B(G317), .Z(new_n743));
  OAI221_X1 g0543(.A(new_n740), .B1(new_n741), .B2(new_n742), .C1(new_n737), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n715), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G329), .A2(new_n745), .B1(new_n721), .B2(G283), .ZN(new_n746));
  INV_X1    g0546(.A(new_n733), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n288), .B1(new_n747), .B2(G322), .ZN(new_n748));
  INV_X1    g0548(.A(G294), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n746), .B(new_n748), .C1(new_n749), .C2(new_n735), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n728), .A2(new_n739), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n330), .A2(KEYINPUT95), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n330), .A2(KEYINPUT95), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n226), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n225), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n710), .ZN(new_n756));
  INV_X1    g0556(.A(new_n288), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n662), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n504), .B2(new_n662), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n229), .A2(G45), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n247), .B2(G45), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n282), .A2(new_n662), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n759), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n751), .A2(new_n755), .B1(new_n756), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n702), .B1(new_n711), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n707), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT96), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G396));
  NOR2_X1   g0569(.A1(new_n755), .A2(new_n708), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n702), .B1(new_n770), .B2(new_n363), .ZN(new_n771));
  INV_X1    g0571(.A(new_n755), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n720), .A2(new_n208), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n288), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n774), .B1(new_n412), .B2(new_n729), .C1(new_n741), .C2(new_n715), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n742), .A2(new_n504), .B1(new_n749), .B2(new_n733), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n727), .A2(new_n537), .B1(new_n737), .B2(new_n777), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n775), .A2(new_n736), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n737), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n780), .A2(G150), .B1(new_n747), .B2(G143), .ZN(new_n781));
  INV_X1    g0581(.A(G137), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n781), .B1(new_n782), .B2(new_n727), .C1(new_n716), .C2(new_n742), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n784));
  XNOR2_X1  g0584(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n282), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n721), .A2(G68), .ZN(new_n787));
  INV_X1    g0587(.A(G132), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n787), .B1(new_n202), .B2(new_n729), .C1(new_n788), .C2(new_n715), .ZN(new_n789));
  INV_X1    g0589(.A(new_n735), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n786), .B(new_n789), .C1(G58), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n779), .B1(new_n785), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n432), .B1(new_n427), .B2(new_n638), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(new_n429), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n429), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n638), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n771), .B1(new_n772), .B2(new_n792), .C1(new_n799), .C2(new_n709), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n689), .B(new_n799), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n703), .B1(new_n801), .B2(new_n688), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(new_n688), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G384));
  OAI211_X1 g0605(.A(G116), .B(new_n227), .C1(new_n474), .C2(KEYINPUT35), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(KEYINPUT35), .B2(new_n474), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT36), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n264), .A2(new_n228), .A3(new_n363), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT98), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n809), .A2(new_n810), .B1(new_n202), .B2(G68), .ZN(new_n812));
  AOI211_X1 g0612(.A(G13), .B(new_n253), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT38), .ZN(new_n815));
  OR2_X1    g0615(.A1(KEYINPUT100), .A2(KEYINPUT16), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n286), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n286), .A2(new_n816), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n258), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n630), .B1(new_n819), .B2(new_n260), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n439), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n325), .B(new_n319), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  INV_X1    g0624(.A(new_n630), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n332), .B2(new_n261), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n333), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n333), .A2(new_n826), .A3(new_n827), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT101), .B1(new_n327), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n819), .A2(new_n260), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n331), .B2(new_n825), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n823), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n829), .A2(new_n831), .B1(new_n834), .B2(KEYINPUT37), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n815), .B1(new_n822), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(KEYINPUT38), .A3(new_n821), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n638), .B(new_n799), .C1(new_n616), .C2(new_n623), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n797), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n369), .A2(new_n638), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n371), .A2(new_n377), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n370), .B(new_n632), .C1(new_n357), .C2(new_n376), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n840), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  AOI211_X1 g0649(.A(KEYINPUT99), .B(new_n849), .C1(new_n841), .C2(new_n797), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n839), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n600), .A2(new_n602), .A3(new_n630), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT102), .B1(new_n298), .B2(new_n317), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT102), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n325), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n826), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n827), .B1(new_n858), .B2(new_n599), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT103), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n824), .B1(new_n823), .B2(new_n828), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n327), .A2(new_n830), .A3(KEYINPUT101), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT103), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n826), .B1(new_n603), .B2(new_n328), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n815), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT104), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT104), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(new_n815), .C1(new_n865), .C2(new_n866), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n868), .A2(new_n869), .A3(new_n838), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n371), .A2(new_n632), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n853), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n438), .A2(new_n698), .A3(new_n442), .A4(new_n691), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n609), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n847), .A2(new_n799), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n686), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n680), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n632), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n681), .B1(new_n684), .B2(new_n638), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT40), .B1(new_n839), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n868), .A2(new_n838), .A3(new_n871), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n889), .B(new_n880), .C1(new_n884), .C2(new_n885), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n443), .B1(new_n885), .B2(new_n884), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n669), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n879), .A2(new_n894), .B1(new_n253), .B2(new_n626), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n879), .A2(new_n894), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n814), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT106), .Z(G367));
  AND2_X1   g0698(.A1(new_n485), .A2(new_n497), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n658), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n468), .A2(new_n470), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n486), .A2(new_n632), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n899), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n485), .B1(new_n905), .B2(new_n593), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n638), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n901), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n524), .A2(new_n638), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n521), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n692), .B2(new_n910), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n909), .A2(KEYINPUT43), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n655), .A2(new_n905), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n663), .B(KEYINPUT41), .Z(new_n922));
  NAND2_X1  g0722(.A1(new_n698), .A2(new_n691), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n683), .A2(new_n687), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G330), .ZN(new_n925));
  INV_X1    g0725(.A(new_n647), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n639), .B1(new_n651), .B2(G330), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n657), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n639), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n706), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n656), .A3(new_n647), .ZN(new_n931));
  AND4_X1   g0731(.A1(new_n923), .A2(new_n925), .A3(new_n928), .A4(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n905), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT44), .B1(new_n660), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT44), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n905), .C1(new_n658), .C2(new_n659), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT45), .B1(new_n660), .B2(new_n933), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT45), .ZN(new_n938));
  NOR4_X1   g0738(.A1(new_n658), .A2(new_n905), .A3(new_n938), .A4(new_n659), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n934), .B(new_n936), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(new_n654), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n940), .A2(KEYINPUT107), .A3(new_n654), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT107), .B1(new_n940), .B2(new_n654), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n932), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n922), .B1(new_n944), .B2(new_n699), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n701), .A2(G1), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n921), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n912), .A2(new_n710), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n710), .B(new_n755), .C1(new_n662), .C2(new_n424), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n239), .A2(new_n762), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n702), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n742), .A2(new_n202), .B1(new_n363), .B2(new_n720), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n757), .B(new_n952), .C1(G137), .C2(new_n745), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n780), .A2(G159), .B1(new_n747), .B2(G150), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n730), .A2(G58), .B1(new_n726), .B2(G143), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n790), .A2(G68), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n729), .A2(new_n504), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT46), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n737), .A2(new_n749), .B1(new_n733), .B2(new_n537), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n959), .A2(new_n282), .A3(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n745), .A2(G317), .B1(new_n726), .B2(G311), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(new_n210), .C2(new_n720), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n742), .A2(new_n777), .B1(new_n735), .B2(new_n412), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT108), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n957), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT47), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n755), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n948), .B(new_n951), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n947), .A2(new_n970), .ZN(G387));
  NOR2_X1   g0771(.A1(new_n932), .A2(new_n664), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n928), .A2(new_n931), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n699), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G150), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n715), .A2(new_n975), .B1(new_n733), .B2(new_n202), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G77), .B2(new_n730), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n721), .A2(G97), .B1(new_n726), .B2(G159), .ZN(new_n978));
  INV_X1    g0778(.A(new_n255), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n780), .A2(new_n979), .B1(new_n722), .B2(G68), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n735), .A2(new_n423), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n786), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n978), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n730), .A2(G294), .B1(new_n790), .B2(G283), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n726), .A2(G322), .B1(new_n722), .B2(G303), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n985), .B1(new_n741), .B2(new_n737), .C1(new_n986), .C2(new_n733), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT48), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n988), .B2(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT49), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G326), .A2(new_n745), .B1(new_n721), .B2(G116), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n786), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n990), .A2(KEYINPUT49), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n983), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n755), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n236), .A2(G45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n979), .A2(new_n202), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g0802(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n665), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n762), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n288), .A2(new_n221), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(G107), .B2(new_n221), .C1(new_n665), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT109), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n756), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(KEYINPUT109), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n999), .B(new_n703), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT111), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n929), .A2(new_n710), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n973), .A2(new_n946), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n974), .A2(new_n1014), .ZN(G393));
  XNOR2_X1  g0815(.A(new_n655), .B(new_n940), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n944), .B(new_n663), .C1(new_n1016), .C2(new_n932), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n905), .A2(new_n710), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n244), .A2(new_n763), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n756), .B1(new_n210), .B2(new_n221), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n703), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n727), .A2(new_n975), .B1(new_n733), .B2(new_n716), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n737), .A2(new_n202), .B1(new_n729), .B2(new_n263), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G143), .B2(new_n745), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n790), .A2(G77), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n773), .B(new_n786), .C1(new_n979), .C2(new_n722), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n745), .A2(G322), .B1(new_n730), .B2(G283), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n757), .C1(new_n412), .C2(new_n720), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  OAI22_X1  g0831(.A1(new_n727), .A2(new_n986), .B1(new_n733), .B2(new_n741), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT52), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n780), .A2(G303), .B1(G294), .B2(new_n722), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n504), .C2(new_n735), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1028), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1021), .B1(new_n1036), .B2(new_n755), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1016), .A2(new_n946), .B1(new_n1018), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1017), .A2(new_n1038), .ZN(G390));
  NAND2_X1  g0839(.A1(new_n842), .A2(new_n847), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n371), .B2(new_n632), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n872), .A2(new_n873), .A3(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n638), .B(new_n795), .C1(new_n697), .C2(new_n616), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n797), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n875), .B1(new_n1044), .B2(new_n847), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n888), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n884), .A2(new_n885), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(G330), .A3(new_n799), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n849), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n688), .A2(new_n799), .A3(new_n847), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1042), .A2(new_n1046), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n438), .A2(new_n1048), .A3(G330), .A4(new_n442), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n877), .A2(new_n1055), .A3(new_n609), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n847), .B1(new_n688), .B2(new_n799), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n842), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1049), .A2(new_n849), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1059), .A2(new_n1052), .A3(new_n797), .A4(new_n1043), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1056), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1054), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1051), .A2(new_n1053), .A3(new_n1061), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n663), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n872), .A2(new_n708), .A3(new_n873), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n742), .A2(new_n1067), .B1(new_n782), .B2(new_n737), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1068), .A2(KEYINPUT113), .B1(new_n716), .B2(new_n735), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(KEYINPUT113), .B2(new_n1068), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT114), .Z(new_n1071));
  INV_X1    g0871(.A(G128), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n727), .A2(new_n1072), .B1(new_n720), .B2(new_n202), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n757), .B1(new_n747), .B2(G132), .ZN(new_n1074));
  OR3_X1    g0874(.A1(new_n729), .A2(KEYINPUT53), .A3(new_n975), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT53), .B1(new_n729), .B2(new_n975), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(G125), .C2(new_n745), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1026), .B1(new_n504), .B2(new_n733), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT115), .Z(new_n1080));
  OAI22_X1  g0880(.A1(new_n727), .A2(new_n777), .B1(new_n715), .B2(new_n749), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n722), .A2(G97), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n787), .A2(new_n757), .A3(new_n731), .A4(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(G107), .C2(new_n780), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1071), .A2(new_n1078), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n772), .B1(new_n1085), .B2(KEYINPUT116), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n702), .B(new_n1088), .C1(new_n255), .C2(new_n770), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n946), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1054), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1065), .A2(new_n1093), .ZN(G378));
  NAND2_X1  g0894(.A1(new_n871), .A2(new_n838), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n859), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n829), .A2(KEYINPUT103), .A3(new_n831), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT103), .B1(new_n829), .B2(new_n831), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n601), .A2(KEYINPUT18), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n599), .A2(new_n334), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n328), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n857), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n870), .B1(new_n1104), .B2(new_n815), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n890), .B1(new_n1095), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n839), .A2(new_n886), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n889), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(G330), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n397), .A2(new_n630), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n409), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n608), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n606), .A2(new_n607), .A3(new_n409), .A4(new_n1110), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1109), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1106), .A2(new_n1121), .A3(G330), .A4(new_n1108), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n876), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n874), .A2(new_n875), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n853), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1123), .A2(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT57), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1042), .A2(new_n1046), .A3(new_n1052), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1050), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1056), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n663), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1056), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1064), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1121), .B1(new_n891), .B2(G330), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1124), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n876), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT57), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1136), .A2(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1072), .A2(new_n733), .B1(new_n729), .B2(new_n1067), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT119), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n726), .A2(G125), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n788), .B2(new_n737), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n742), .A2(new_n782), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1148), .B(new_n1152), .C1(new_n975), .C2(new_n735), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(G33), .A2(G41), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT117), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n745), .B2(G124), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1154), .B(new_n1157), .C1(new_n716), .C2(new_n720), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT58), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n721), .A2(G58), .B1(new_n730), .B2(G77), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n747), .A2(G107), .B1(new_n726), .B2(G116), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n956), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n282), .A2(G41), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n742), .A2(new_n423), .B1(new_n715), .B2(new_n777), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G97), .B2(new_n780), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1158), .A2(new_n1159), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1156), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1164), .A2(G50), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1167), .B2(new_n1160), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT118), .Z(new_n1172));
  OAI21_X1  g0972(.A(new_n755), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n702), .B1(new_n770), .B2(new_n202), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n1121), .C2(new_n709), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1144), .B2(new_n946), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1146), .A2(new_n1177), .ZN(G375));
  NAND2_X1  g0978(.A1(new_n849), .A2(new_n708), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT121), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n747), .A2(G137), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n716), .B2(new_n729), .C1(new_n737), .C2(new_n1067), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n720), .A2(new_n262), .B1(new_n715), .B2(new_n1072), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n727), .A2(new_n788), .B1(new_n742), .B2(new_n975), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n282), .B1(new_n202), .B2(new_n735), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n715), .A2(new_n537), .B1(new_n729), .B2(new_n210), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT122), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n727), .A2(new_n749), .B1(new_n733), .B2(new_n777), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n742), .A2(new_n412), .B1(new_n504), .B2(new_n737), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n757), .B1(new_n720), .B2(new_n363), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n981), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1186), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n772), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n702), .B(new_n1194), .C1(new_n263), .C2(new_n770), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1134), .A2(new_n946), .B1(new_n1180), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n922), .B(KEYINPUT120), .Z(new_n1198));
  AND2_X1   g0998(.A1(new_n1062), .A2(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1056), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1197), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G381));
  AOI21_X1  g1003(.A(new_n664), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1092), .B1(new_n1064), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1146), .A2(new_n1205), .A3(new_n1177), .ZN(new_n1206));
  INV_X1    g1006(.A(G384), .ZN(new_n1207));
  INV_X1    g1007(.A(G390), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n974), .A2(new_n768), .A3(new_n1014), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1202), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  OR3_X1    g1011(.A1(new_n1206), .A2(G387), .A3(new_n1211), .ZN(G407));
  NAND2_X1  g1012(.A1(new_n631), .A2(G213), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1206), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(G407), .A2(new_n1214), .A3(G213), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(G407), .A2(KEYINPUT123), .A3(G213), .A4(new_n1214), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(G409));
  AOI21_X1  g1019(.A(new_n768), .B1(new_n974), .B2(new_n1014), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT126), .B1(new_n1210), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1220), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1209), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G390), .B1(new_n947), .B2(new_n970), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n947), .A2(new_n970), .A3(G390), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(KEYINPUT127), .B2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1226), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1222), .A2(new_n1209), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1227), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G378), .B(new_n1177), .C1(new_n1136), .C2(new_n1145), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1138), .A2(new_n1144), .A3(new_n1198), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1175), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1142), .A2(KEYINPUT124), .A3(new_n1143), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1091), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1205), .B1(new_n1238), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1236), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1062), .A2(new_n663), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT60), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1200), .A2(new_n1248), .A3(new_n1056), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1207), .B1(new_n1250), .B2(new_n1197), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1247), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1061), .A2(new_n664), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(G384), .A3(new_n1196), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1244), .A2(new_n1245), .A3(new_n1213), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1213), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1236), .B2(new_n1243), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1260), .A2(G2897), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1251), .A2(new_n1255), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1251), .B2(new_n1255), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1258), .B(new_n1259), .C1(new_n1261), .C2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1260), .B(new_n1256), .C1(new_n1236), .C2(new_n1243), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n1245), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1235), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1265), .B1(new_n1261), .B2(KEYINPUT125), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1244), .A2(new_n1213), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1259), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1267), .B2(KEYINPUT63), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1271), .B2(new_n1256), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1269), .A2(new_n1279), .ZN(G405));
  NAND2_X1  g1080(.A1(new_n1235), .A2(new_n1257), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1256), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(G375), .B(new_n1205), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1283), .B(new_n1284), .ZN(G402));
endmodule


