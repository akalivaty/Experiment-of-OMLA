

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U323 ( .A(n392), .B(n391), .ZN(n537) );
  XNOR2_X1 U324 ( .A(n415), .B(KEYINPUT54), .ZN(n416) );
  XNOR2_X1 U325 ( .A(n301), .B(n300), .ZN(n308) );
  XOR2_X1 U326 ( .A(n363), .B(n307), .Z(n291) );
  XNOR2_X1 U327 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n464) );
  XNOR2_X1 U328 ( .A(n465), .B(n464), .ZN(n469) );
  XNOR2_X1 U329 ( .A(n404), .B(n403), .ZN(n405) );
  INV_X1 U330 ( .A(KEYINPUT10), .ZN(n294) );
  XNOR2_X1 U331 ( .A(n453), .B(n405), .ZN(n406) );
  XNOR2_X1 U332 ( .A(n293), .B(n292), .ZN(n339) );
  XNOR2_X1 U333 ( .A(n339), .B(n294), .ZN(n296) );
  XNOR2_X1 U334 ( .A(n390), .B(KEYINPUT48), .ZN(n391) );
  XNOR2_X1 U335 ( .A(n417), .B(n416), .ZN(n440) );
  XNOR2_X1 U336 ( .A(n441), .B(KEYINPUT55), .ZN(n442) );
  XNOR2_X1 U337 ( .A(n443), .B(n442), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n308), .B(n291), .ZN(n562) );
  XNOR2_X1 U339 ( .A(n414), .B(n413), .ZN(n527) );
  XNOR2_X1 U340 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U341 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U342 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(G99GAT), .B(G106GAT), .Z(n293) );
  XNOR2_X1 U345 ( .A(G85GAT), .B(KEYINPUT71), .ZN(n292) );
  XOR2_X1 U346 ( .A(G162GAT), .B(G50GAT), .Z(n320) );
  XNOR2_X1 U347 ( .A(n320), .B(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n301) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(G36GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n297), .B(G190GAT), .ZN(n404) );
  XOR2_X1 U351 ( .A(n404), .B(G92GAT), .Z(n299) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT68), .B(G43GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(G29GAT), .B(n304), .Z(n363) );
  XOR2_X1 U358 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n306) );
  XNOR2_X1 U359 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  INV_X1 U361 ( .A(n562), .ZN(n493) );
  XOR2_X1 U362 ( .A(KEYINPUT89), .B(KEYINPUT2), .Z(n310) );
  XNOR2_X1 U363 ( .A(KEYINPUT88), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U365 ( .A(KEYINPUT3), .B(n311), .Z(n433) );
  XOR2_X1 U366 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n313) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n314), .B(KEYINPUT22), .Z(n319) );
  XOR2_X1 U370 ( .A(G197GAT), .B(KEYINPUT87), .Z(n316) );
  XNOR2_X1 U371 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n394) );
  XNOR2_X1 U373 ( .A(G148GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n317), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U375 ( .A(n394), .B(n338), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U377 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n322) );
  XOR2_X1 U378 ( .A(G155GAT), .B(G22GAT), .Z(n352) );
  XNOR2_X1 U379 ( .A(n320), .B(n352), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U381 ( .A(n324), .B(n323), .Z(n326) );
  XNOR2_X1 U382 ( .A(G218GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n433), .B(n327), .ZN(n475) );
  XOR2_X1 U385 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n329) );
  XNOR2_X1 U386 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U388 ( .A(KEYINPUT72), .B(G120GAT), .Z(n331) );
  NAND2_X1 U389 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(n333), .B(n332), .Z(n337) );
  XNOR2_X1 U392 ( .A(G57GAT), .B(G71GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n334), .B(KEYINPUT13), .ZN(n355) );
  XNOR2_X1 U394 ( .A(G92GAT), .B(G64GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n335), .B(G176GAT), .ZN(n393) );
  XNOR2_X1 U396 ( .A(n355), .B(n393), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n381) );
  XOR2_X1 U400 ( .A(KEYINPUT36), .B(n562), .Z(n590) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n343) );
  XNOR2_X1 U402 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT78), .B(G64GAT), .Z(n345) );
  XNOR2_X1 U405 ( .A(G78GAT), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U407 ( .A(n346), .B(KEYINPUT12), .Z(n348) );
  XOR2_X1 U408 ( .A(G183GAT), .B(G8GAT), .Z(n409) );
  XNOR2_X1 U409 ( .A(G127GAT), .B(n409), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n360) );
  XNOR2_X1 U412 ( .A(G1GAT), .B(G15GAT), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n351), .B(KEYINPUT69), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n352), .B(n362), .ZN(n354) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n492) );
  NOR2_X1 U421 ( .A1(n590), .A2(n492), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n361), .B(KEYINPUT45), .ZN(n378) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U424 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U426 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n367) );
  XNOR2_X1 U427 ( .A(G113GAT), .B(G8GAT), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n377) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XOR2_X1 U431 ( .A(G197GAT), .B(G169GAT), .Z(n371) );
  XNOR2_X1 U432 ( .A(G141GAT), .B(G22GAT), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U434 ( .A(G36GAT), .B(G50GAT), .Z(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n566) );
  NAND2_X1 U438 ( .A1(n378), .A2(n566), .ZN(n379) );
  NOR2_X1 U439 ( .A1(n381), .A2(n379), .ZN(n389) );
  XOR2_X1 U440 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n387) );
  INV_X1 U441 ( .A(KEYINPUT65), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(KEYINPUT41), .B(n382), .ZN(n571) );
  NOR2_X1 U444 ( .A1(n566), .A2(n571), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(KEYINPUT46), .ZN(n384) );
  NOR2_X1 U446 ( .A1(n384), .A2(n562), .ZN(n385) );
  XOR2_X1 U447 ( .A(n492), .B(KEYINPUT111), .Z(n575) );
  AND2_X1 U448 ( .A1(n385), .A2(n575), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n388) );
  NOR2_X1 U450 ( .A1(n389), .A2(n388), .ZN(n392) );
  XOR2_X1 U451 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n390) );
  INV_X1 U452 ( .A(n409), .ZN(n408) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n407) );
  INV_X1 U454 ( .A(KEYINPUT83), .ZN(n402) );
  XNOR2_X1 U455 ( .A(KEYINPUT18), .B(G169GAT), .ZN(n400) );
  INV_X1 U456 ( .A(KEYINPUT17), .ZN(n395) );
  NAND2_X1 U457 ( .A1(KEYINPUT19), .A2(n395), .ZN(n398) );
  INV_X1 U458 ( .A(KEYINPUT19), .ZN(n396) );
  NAND2_X1 U459 ( .A1(n396), .A2(KEYINPUT17), .ZN(n397) );
  NAND2_X1 U460 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n453) );
  XOR2_X1 U463 ( .A(KEYINPUT93), .B(G204GAT), .Z(n403) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n410) );
  OR2_X1 U465 ( .A1(n408), .A2(n410), .ZN(n412) );
  NAND2_X1 U466 ( .A1(n408), .A2(n410), .ZN(n411) );
  NAND2_X1 U467 ( .A1(n412), .A2(n411), .ZN(n414) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  NOR2_X1 U469 ( .A1(n537), .A2(n527), .ZN(n417) );
  INV_X1 U470 ( .A(KEYINPUT119), .ZN(n415) );
  XOR2_X1 U471 ( .A(G57GAT), .B(G148GAT), .Z(n419) );
  XNOR2_X1 U472 ( .A(G85GAT), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U474 ( .A(G29GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n437) );
  XOR2_X1 U476 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n423) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U479 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n425) );
  XNOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n435) );
  XOR2_X1 U483 ( .A(G127GAT), .B(G113GAT), .Z(n429) );
  XNOR2_X1 U484 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U486 ( .A(n430), .B(KEYINPUT0), .Z(n432) );
  XNOR2_X1 U487 ( .A(G120GAT), .B(G134GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n454) );
  XNOR2_X1 U489 ( .A(n433), .B(n454), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n439) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n506) );
  INV_X1 U494 ( .A(n506), .ZN(n524) );
  NAND2_X1 U495 ( .A1(n440), .A2(n524), .ZN(n578) );
  NOR2_X1 U496 ( .A1(n475), .A2(n578), .ZN(n443) );
  INV_X1 U497 ( .A(KEYINPUT120), .ZN(n441) );
  XOR2_X1 U498 ( .A(G15GAT), .B(G99GAT), .Z(n445) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(G71GAT), .B(n446), .Z(n448) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n450) );
  XNOR2_X1 U505 ( .A(G183GAT), .B(G176GAT), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U507 ( .A(n452), .B(n451), .Z(n456) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n530) );
  INV_X1 U510 ( .A(n530), .ZN(n539) );
  NAND2_X1 U511 ( .A1(n457), .A2(n539), .ZN(n574) );
  NOR2_X1 U512 ( .A1(n493), .A2(n574), .ZN(n461) );
  XNOR2_X1 U513 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n459) );
  XNOR2_X1 U514 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n458) );
  NOR2_X1 U515 ( .A1(n381), .A2(n566), .ZN(n497) );
  NOR2_X1 U516 ( .A1(n530), .A2(n527), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT96), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n475), .A2(n463), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n475), .A2(n530), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT95), .B(n466), .Z(n467) );
  XNOR2_X1 U521 ( .A(KEYINPUT26), .B(n467), .ZN(n579) );
  XNOR2_X1 U522 ( .A(n527), .B(KEYINPUT27), .ZN(n473) );
  NOR2_X1 U523 ( .A1(n579), .A2(n473), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT98), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n471), .A2(n506), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT99), .ZN(n479) );
  NOR2_X1 U528 ( .A1(n524), .A2(n473), .ZN(n474) );
  XOR2_X1 U529 ( .A(KEYINPUT94), .B(n474), .Z(n538) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n476) );
  XNOR2_X1 U531 ( .A(n476), .B(n475), .ZN(n509) );
  NOR2_X1 U532 ( .A1(n538), .A2(n509), .ZN(n477) );
  NAND2_X1 U533 ( .A1(n477), .A2(n530), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n496) );
  NAND2_X1 U535 ( .A1(n496), .A2(n492), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n590), .A2(n480), .ZN(n482) );
  XNOR2_X1 U537 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n482), .B(n481), .ZN(n523) );
  NAND2_X1 U539 ( .A1(n497), .A2(n523), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT38), .B(n483), .Z(n510) );
  NAND2_X1 U541 ( .A1(n510), .A2(n539), .ZN(n487) );
  XOR2_X1 U542 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n485) );
  INV_X1 U543 ( .A(G43GAT), .ZN(n484) );
  INV_X1 U544 ( .A(n527), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n510), .A2(n488), .ZN(n491) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(G36GAT), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1329GAT) );
  INV_X1 U549 ( .A(n492), .ZN(n586) );
  NAND2_X1 U550 ( .A1(n493), .A2(n586), .ZN(n494) );
  XOR2_X1 U551 ( .A(KEYINPUT16), .B(n494), .Z(n495) );
  AND2_X1 U552 ( .A1(n496), .A2(n495), .ZN(n512) );
  NAND2_X1 U553 ( .A1(n497), .A2(n512), .ZN(n503) );
  NOR2_X1 U554 ( .A1(n524), .A2(n503), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT34), .B(n498), .Z(n499) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NOR2_X1 U557 ( .A1(n527), .A2(n503), .ZN(n500) );
  XOR2_X1 U558 ( .A(G8GAT), .B(n500), .Z(G1325GAT) );
  NOR2_X1 U559 ( .A1(n530), .A2(n503), .ZN(n502) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  INV_X1 U562 ( .A(n509), .ZN(n540) );
  NOR2_X1 U563 ( .A1(n540), .A2(n503), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT100), .B(n504), .Z(n505) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  XOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .Z(n508) );
  NAND2_X1 U567 ( .A1(n506), .A2(n510), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  NAND2_X1 U569 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U570 ( .A(n511), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U571 ( .A(n566), .ZN(n580) );
  NOR2_X1 U572 ( .A1(n580), .A2(n571), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n522), .A2(n512), .ZN(n518) );
  NOR2_X1 U574 ( .A1(n524), .A2(n518), .ZN(n513) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n527), .A2(n518), .ZN(n515) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n530), .A2(n518), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n540), .A2(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n524), .A2(n533), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n533), .ZN(n528) );
  XOR2_X1 U591 ( .A(KEYINPUT108), .B(n528), .Z(n529) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n533), .ZN(n532) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U596 ( .A1(n540), .A2(n533), .ZN(n535) );
  XNOR2_X1 U597 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  OR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U602 ( .A1(n551), .A2(n541), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n548), .A2(n580), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  INV_X1 U606 ( .A(n571), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n548), .A2(n555), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  INV_X1 U609 ( .A(n548), .ZN(n545) );
  NOR2_X1 U610 ( .A1(n575), .A2(n545), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U614 ( .A1(n548), .A2(n562), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT115), .Z(n554) );
  NOR2_X1 U617 ( .A1(n579), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT114), .B(n552), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n580), .A2(n563), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XNOR2_X1 U621 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n559) );
  XOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .Z(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n563), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT117), .Z(n561) );
  NAND2_X1 U627 ( .A1(n563), .A2(n586), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT118), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n565), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n574), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n571), .A2(n574), .ZN(n572) );
  XOR2_X1 U639 ( .A(n573), .B(n572), .Z(G1349GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1350GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n588) );
  NAND2_X1 U645 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n588), .A2(n381), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n588), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(G218GAT), .B(n593), .Z(G1355GAT) );
endmodule

