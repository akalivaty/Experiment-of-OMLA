

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X2 U325 ( .A(n409), .B(n425), .Z(n489) );
  NOR2_X1 U326 ( .A1(n584), .A2(n482), .ZN(n483) );
  XNOR2_X1 U327 ( .A(n457), .B(KEYINPUT96), .ZN(n458) );
  XOR2_X1 U328 ( .A(KEYINPUT38), .B(n485), .Z(n496) );
  XOR2_X1 U329 ( .A(n402), .B(n401), .Z(n293) );
  XOR2_X1 U330 ( .A(G64GAT), .B(G92GAT), .Z(n294) );
  XNOR2_X1 U331 ( .A(n319), .B(KEYINPUT10), .ZN(n320) );
  XNOR2_X1 U332 ( .A(n321), .B(n320), .ZN(n324) );
  INV_X1 U333 ( .A(KEYINPUT97), .ZN(n469) );
  OR2_X1 U334 ( .A1(n468), .A2(n467), .ZN(n470) );
  XNOR2_X1 U335 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U336 ( .A(n470), .B(n469), .ZN(n481) );
  XNOR2_X1 U337 ( .A(n331), .B(n330), .ZN(n388) );
  INV_X1 U338 ( .A(G190GAT), .ZN(n450) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U340 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT82), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(n297), .ZN(n444) );
  XOR2_X1 U345 ( .A(KEYINPUT65), .B(KEYINPUT83), .Z(n299) );
  XNOR2_X1 U346 ( .A(G15GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n300), .B(G99GAT), .Z(n302) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n370) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(n370), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(n444), .B(n303), .Z(n316) );
  XOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT87), .Z(n305) );
  XNOR2_X1 U354 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U356 ( .A(G183GAT), .B(n306), .Z(n308) );
  NAND2_X1 U357 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n309), .B(KEYINPUT85), .Z(n314) );
  XOR2_X1 U360 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n311) );
  XNOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(G169GAT), .B(n312), .Z(n405) );
  XNOR2_X1 U364 ( .A(n405), .B(KEYINPUT88), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U366 ( .A(n316), .B(n315), .Z(n520) );
  INV_X1 U367 ( .A(n520), .ZN(n531) );
  XOR2_X1 U368 ( .A(G36GAT), .B(G190GAT), .Z(n398) );
  XOR2_X1 U369 ( .A(G50GAT), .B(G162GAT), .Z(n414) );
  XOR2_X1 U370 ( .A(G29GAT), .B(G43GAT), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n362) );
  XNOR2_X1 U373 ( .A(n414), .B(n362), .ZN(n321) );
  AND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n322), .B(KEYINPUT75), .ZN(n373) );
  XOR2_X1 U377 ( .A(n373), .B(KEYINPUT11), .Z(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U379 ( .A(n398), .B(n325), .Z(n331) );
  XOR2_X1 U380 ( .A(KEYINPUT9), .B(KEYINPUT78), .Z(n327) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(G92GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n329) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(G218GAT), .ZN(n328) );
  XOR2_X1 U384 ( .A(KEYINPUT36), .B(n388), .Z(n584) );
  XOR2_X1 U385 ( .A(G211GAT), .B(G71GAT), .Z(n333) );
  XNOR2_X1 U386 ( .A(G22GAT), .B(G127GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n348) );
  XOR2_X1 U388 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n335) );
  XNOR2_X1 U389 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .Z(n401) );
  XOR2_X1 U392 ( .A(n401), .B(G78GAT), .Z(n337) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n354) );
  XNOR2_X1 U394 ( .A(n354), .B(G155GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U396 ( .A(n339), .B(n338), .Z(n341) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U399 ( .A(n342), .B(KEYINPUT14), .Z(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n344) );
  XNOR2_X1 U401 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n369) );
  XNOR2_X1 U403 ( .A(n369), .B(KEYINPUT15), .ZN(n345) );
  XOR2_X1 U404 ( .A(n346), .B(n345), .Z(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n551) );
  INV_X1 U406 ( .A(n551), .ZN(n563) );
  NOR2_X1 U407 ( .A1(n584), .A2(n563), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n349), .B(KEYINPUT45), .ZN(n386) );
  XOR2_X1 U409 ( .A(G8GAT), .B(G113GAT), .Z(n351) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(G197GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n366) );
  XOR2_X1 U412 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n353) );
  XNOR2_X1 U413 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U415 ( .A(G36GAT), .B(G50GAT), .Z(n356) );
  XOR2_X1 U416 ( .A(G141GAT), .B(G22GAT), .Z(n415) );
  XNOR2_X1 U417 ( .A(n415), .B(n354), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U419 ( .A(n358), .B(n357), .Z(n360) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U422 ( .A(n361), .B(KEYINPUT69), .Z(n364) );
  XNOR2_X1 U423 ( .A(n362), .B(KEYINPUT70), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n499) );
  INV_X1 U426 ( .A(n499), .ZN(n570) );
  XOR2_X1 U427 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n368) );
  XNOR2_X1 U428 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n383) );
  XOR2_X1 U430 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n372) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U433 ( .A(n373), .B(KEYINPUT73), .Z(n375) );
  NAND2_X1 U434 ( .A1(G230GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U436 ( .A(n377), .B(n376), .Z(n381) );
  XNOR2_X1 U437 ( .A(G106GAT), .B(G78GAT), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n378), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U439 ( .A(G176GAT), .B(G204GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n294), .B(n379), .ZN(n397) );
  XNOR2_X1 U441 ( .A(n422), .B(n397), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n575) );
  INV_X1 U444 ( .A(n575), .ZN(n384) );
  NOR2_X1 U445 ( .A1(n570), .A2(n384), .ZN(n385) );
  AND2_X1 U446 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n387), .B(KEYINPUT113), .ZN(n395) );
  XNOR2_X1 U448 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n389), .B(n575), .ZN(n558) );
  NAND2_X1 U450 ( .A1(n570), .A2(n558), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n390), .B(KEYINPUT46), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n391), .A2(n563), .ZN(n392) );
  NOR2_X1 U453 ( .A1(n388), .A2(n392), .ZN(n393) );
  XNOR2_X1 U454 ( .A(KEYINPUT47), .B(n393), .ZN(n394) );
  NAND2_X1 U455 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n396), .B(KEYINPUT48), .ZN(n528) );
  XOR2_X1 U457 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U460 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n293), .B(n403), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U463 ( .A(KEYINPUT89), .B(G218GAT), .Z(n407) );
  XNOR2_X1 U464 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U466 ( .A(G197GAT), .B(n408), .ZN(n425) );
  INV_X1 U467 ( .A(n489), .ZN(n517) );
  NAND2_X1 U468 ( .A1(n528), .A2(n517), .ZN(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n567) );
  XOR2_X1 U471 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT22), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U474 ( .A(G204GAT), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U481 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n424), .B(KEYINPUT3), .ZN(n436) );
  XOR2_X1 U483 ( .A(n425), .B(n436), .Z(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n461) );
  XOR2_X1 U485 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n443) );
  XOR2_X1 U488 ( .A(G162GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(G120GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U491 ( .A(G57GAT), .B(KEYINPUT1), .Z(n433) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n441) );
  XOR2_X1 U495 ( .A(G85GAT), .B(n436), .Z(n438) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U498 ( .A(G29GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n514) );
  NOR2_X1 U502 ( .A1(n461), .A2(n514), .ZN(n446) );
  AND2_X1 U503 ( .A1(n567), .A2(n446), .ZN(n447) );
  XOR2_X1 U504 ( .A(n447), .B(KEYINPUT55), .Z(n448) );
  XNOR2_X1 U505 ( .A(n448), .B(KEYINPUT121), .ZN(n449) );
  NOR2_X2 U506 ( .A1(n531), .A2(n449), .ZN(n564) );
  NAND2_X1 U507 ( .A1(n564), .A2(n388), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n474) );
  OR2_X1 U510 ( .A1(n563), .A2(n388), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n454), .B(KEYINPUT16), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT81), .ZN(n471) );
  INV_X1 U513 ( .A(n514), .ZN(n566) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(n489), .ZN(n463) );
  NOR2_X1 U515 ( .A1(n566), .A2(n463), .ZN(n529) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT28), .ZN(n456) );
  XOR2_X1 U517 ( .A(n456), .B(KEYINPUT66), .Z(n495) );
  NAND2_X1 U518 ( .A1(n529), .A2(n495), .ZN(n457) );
  NOR2_X1 U519 ( .A1(n458), .A2(n520), .ZN(n468) );
  NOR2_X1 U520 ( .A1(n531), .A2(n489), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n461), .A2(n459), .ZN(n460) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n460), .Z(n465) );
  NAND2_X1 U523 ( .A1(n461), .A2(n531), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U525 ( .A1(n569), .A2(n463), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n514), .A2(n466), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n471), .A2(n481), .ZN(n500) );
  NAND2_X1 U529 ( .A1(n570), .A2(n575), .ZN(n484) );
  NOR2_X1 U530 ( .A1(n500), .A2(n484), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT98), .ZN(n479) );
  NAND2_X1 U532 ( .A1(n514), .A2(n479), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n479), .A2(n517), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U538 ( .A1(n479), .A2(n520), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  INV_X1 U540 ( .A(n495), .ZN(n534) );
  NAND2_X1 U541 ( .A1(n479), .A2(n534), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n563), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n483), .ZN(n513) );
  NOR2_X1 U545 ( .A1(n513), .A2(n484), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n496), .A2(n566), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT100), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(n488), .ZN(G1328GAT) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n491) );
  NOR2_X1 U551 ( .A1(n496), .A2(n489), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1329GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n493) );
  NOR2_X1 U554 ( .A1(n531), .A2(n496), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U556 ( .A(G43GAT), .B(n494), .Z(G1330GAT) );
  NOR2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n502) );
  NAND2_X1 U561 ( .A1(n499), .A2(n558), .ZN(n512) );
  NOR2_X1 U562 ( .A1(n500), .A2(n512), .ZN(n507) );
  NAND2_X1 U563 ( .A1(n507), .A2(n514), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  XOR2_X1 U566 ( .A(G64GAT), .B(KEYINPUT105), .Z(n505) );
  NAND2_X1 U567 ( .A1(n507), .A2(n517), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n520), .A2(n507), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U572 ( .A1(n507), .A2(n534), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT106), .Z(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n516) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n514), .A2(n524), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  XOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U581 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n522) );
  NAND2_X1 U584 ( .A1(n524), .A2(n520), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n526) );
  NAND2_X1 U588 ( .A1(n524), .A2(n534), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  NAND2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n530), .B(KEYINPUT114), .ZN(n545) );
  NOR2_X1 U593 ( .A1(n531), .A2(n545), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n532), .B(KEYINPUT115), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n570), .A2(n542), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U599 ( .A1(n542), .A2(n558), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U603 ( .A1(n542), .A2(n551), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U607 ( .A1(n542), .A2(n388), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n547) );
  NOR2_X1 U610 ( .A1(n545), .A2(n569), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n570), .A2(n554), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U614 ( .A1(n554), .A2(n558), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT119), .Z(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n388), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n564), .A2(n570), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT122), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  NAND2_X1 U626 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  INV_X1 U630 ( .A(n563), .ZN(n580) );
  NAND2_X1 U631 ( .A1(n564), .A2(n580), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .Z(n572) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  INV_X1 U640 ( .A(n581), .ZN(n583) );
  NOR2_X1 U641 ( .A1(n583), .A2(n575), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

