//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  XOR2_X1   g000(.A(G113), .B(G122), .Z(new_n187));
  XOR2_X1   g001(.A(KEYINPUT85), .B(G104), .Z(new_n188));
  XOR2_X1   g002(.A(new_n187), .B(new_n188), .Z(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G143), .A4(G214), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT83), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT64), .A2(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT64), .A2(G143), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n200), .A2(new_n190), .A3(new_n191), .A4(G214), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT18), .A2(G131), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n194), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT72), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(G146), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n205), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n194), .B2(new_n202), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT18), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n217), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n194), .A2(new_n216), .A3(new_n202), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n211), .A2(KEYINPUT16), .A3(new_n212), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT16), .ZN(new_n226));
  INV_X1    g040(.A(G125), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G140), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n228), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n221), .B2(new_n220), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n189), .B(new_n219), .C1(new_n224), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT19), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n206), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n211), .A2(KEYINPUT19), .A3(new_n212), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n207), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n222), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n232), .B(new_n240), .C1(new_n241), .C2(new_n217), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n219), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n189), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(G475), .A2(G902), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT86), .B1(new_n236), .B2(new_n245), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(KEYINPUT20), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n246), .A2(KEYINPUT86), .A3(new_n251), .A4(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n199), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(new_n255), .C1(G128), .C2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT64), .B(G143), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n256), .A2(G128), .ZN(new_n261));
  OAI21_X1  g075(.A(G134), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g077(.A1(KEYINPUT68), .A2(G116), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT68), .A2(G116), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(G122), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  INV_X1    g081(.A(G122), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G116), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n264), .A2(KEYINPUT14), .A3(G122), .A4(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n269), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(G107), .C1(new_n272), .C2(KEYINPUT14), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT9), .B(G234), .ZN(new_n275));
  INV_X1    g089(.A(G217), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(G953), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n261), .B1(new_n260), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n254), .A2(KEYINPUT89), .A3(new_n278), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT89), .B1(new_n254), .B2(new_n278), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n283), .A2(G134), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n272), .A2(G107), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n270), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n257), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n274), .B(new_n277), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n277), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(G134), .B2(new_n283), .ZN(new_n290));
  INV_X1    g104(.A(new_n274), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G478), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(KEYINPUT15), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n219), .B1(new_n224), .B2(new_n235), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n244), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n233), .B1(KEYINPUT17), .B2(new_n217), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n301), .A2(new_n223), .B1(new_n215), .B2(new_n218), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT87), .B1(new_n302), .B2(new_n189), .ZN(new_n303));
  INV_X1    g117(.A(new_n236), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n297), .B(new_n300), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G475), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n253), .A2(new_n296), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT82), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n207), .B1(new_n197), .B2(new_n198), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n207), .A2(G143), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(KEYINPUT0), .A2(G128), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n256), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT64), .A2(G143), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(G146), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n256), .A2(G146), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(new_n316), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n227), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n312), .A2(new_n314), .B1(G128), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n323), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n323), .A2(new_n333), .A3(new_n325), .A4(new_n330), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n329), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n327), .B1(new_n335), .B2(new_n227), .ZN(new_n336));
  INV_X1    g150(.A(G224), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G953), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(new_n340), .B2(G107), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n267), .A3(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(G107), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G101), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n349), .A3(new_n346), .A4(G101), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n341), .A2(new_n343), .A3(new_n351), .A4(new_n344), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n345), .B2(G101), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n348), .A2(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT67), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n264), .A2(KEYINPUT69), .A3(G119), .A4(new_n265), .ZN(new_n356));
  AND2_X1   g170(.A1(KEYINPUT68), .A2(G116), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT68), .A2(G116), .ZN(new_n358));
  INV_X1    g172(.A(G119), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(G116), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT69), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n355), .B(new_n356), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT2), .B(G113), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n264), .A2(G119), .A3(new_n265), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n362), .A3(new_n361), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(new_n355), .A3(new_n365), .A4(new_n356), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n354), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n344), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n340), .A2(G107), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n352), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n356), .B1(new_n360), .B2(new_n363), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n366), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n380));
  OAI21_X1  g194(.A(G113), .B1(new_n361), .B2(KEYINPUT5), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n377), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G122), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n372), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n372), .B2(new_n382), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT81), .B(KEYINPUT6), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(new_n382), .ZN(new_n387));
  INV_X1    g201(.A(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n339), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n338), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n336), .A2(new_n395), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n394), .B(new_n327), .C1(new_n335), .C2(new_n227), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n372), .A2(new_n382), .A3(new_n383), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n383), .B(KEYINPUT8), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n379), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n381), .B1(new_n378), .B2(KEYINPUT5), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n376), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n401), .B1(new_n382), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n399), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n297), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n311), .B1(new_n392), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n339), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n390), .B1(new_n389), .B2(new_n399), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n385), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n405), .A2(new_n396), .A3(new_n397), .ZN(new_n414));
  AOI21_X1  g228(.A(G902), .B1(new_n414), .B2(new_n399), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n415), .A3(new_n310), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(G234), .A2(G237), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G952), .A3(new_n191), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT90), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT21), .B(G898), .Z(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(G902), .A3(G953), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n307), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n432));
  AOI221_X4 g246(.A(new_n329), .B1(new_n352), .B2(new_n375), .C1(new_n332), .C2(new_n334), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n332), .A2(new_n334), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n259), .B1(new_n312), .B2(KEYINPUT1), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n324), .B1(new_n199), .B2(G146), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n323), .A2(new_n325), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT1), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n258), .B2(new_n207), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT76), .B(new_n439), .C1(new_n441), .C2(new_n259), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n433), .B1(new_n377), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT11), .B1(new_n255), .B2(G137), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G134), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT65), .B1(new_n447), .B2(G134), .ZN(new_n450));
  OR3_X1    g264(.A1(new_n447), .A2(KEYINPUT65), .A3(G134), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G131), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n449), .A2(new_n216), .A3(new_n451), .A4(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n431), .B(new_n432), .C1(new_n444), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n443), .A2(new_n377), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n335), .A2(new_n376), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(KEYINPUT77), .A3(new_n430), .A4(new_n455), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT10), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n437), .A2(new_n316), .B1(new_n315), .B2(new_n318), .ZN(new_n465));
  INV_X1    g279(.A(new_n329), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n333), .B1(new_n437), .B2(new_n330), .ZN(new_n467));
  INV_X1    g281(.A(new_n334), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n376), .A2(new_n463), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n354), .A2(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n464), .A2(new_n471), .A3(new_n456), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n191), .A2(G227), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT79), .B1(new_n457), .B2(new_n461), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n429), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n457), .A2(new_n461), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT79), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(KEYINPUT80), .A3(new_n477), .A4(new_n462), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n469), .A2(new_n470), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n348), .A2(new_n350), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n353), .A2(new_n352), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n465), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT10), .B1(new_n443), .B2(new_n377), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n455), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT78), .B(new_n455), .C1(new_n489), .C2(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n472), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n475), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n484), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n297), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n457), .A2(new_n472), .A3(new_n461), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n495), .A2(new_n477), .B1(new_n501), .B2(new_n475), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G469), .ZN(new_n503));
  NAND2_X1  g317(.A1(G469), .A2(G902), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G221), .ZN(new_n506));
  INV_X1    g320(.A(new_n275), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n297), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n428), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n371), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n255), .A2(G137), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n447), .A2(G134), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n454), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n434), .B2(new_n466), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n313), .B1(new_n258), .B2(new_n207), .ZN(new_n517));
  INV_X1    g331(.A(new_n318), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n326), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n454), .B2(new_n453), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT30), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n455), .A2(new_n465), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n335), .C2(new_n515), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n511), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n516), .A2(new_n520), .A3(new_n371), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n190), .A2(new_n191), .A3(G210), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n527), .B(KEYINPUT27), .Z(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT26), .B(G101), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NOR4_X1   g344(.A1(new_n525), .A2(KEYINPUT31), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n530), .ZN(new_n532));
  INV_X1    g346(.A(new_n515), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n469), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n511), .B1(new_n534), .B2(new_n522), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT28), .B1(new_n535), .B2(new_n526), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n522), .A3(new_n511), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT28), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT70), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n521), .A2(new_n524), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n371), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n537), .A3(new_n532), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT31), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n541), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G472), .A2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(KEYINPUT32), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n551), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n536), .A2(new_n532), .A3(new_n539), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n525), .A2(new_n526), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n532), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n561), .B(new_n297), .C1(new_n559), .C2(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G472), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n550), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n551), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n554), .A2(new_n557), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n276), .B1(G234), .B2(new_n297), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n232), .A2(new_n208), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n359), .B2(G128), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  INV_X1    g385(.A(G110), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n359), .A2(G128), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n259), .A2(G119), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G110), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT74), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n575), .A2(new_n583), .A3(new_n576), .A4(new_n580), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n568), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n570), .A2(new_n573), .A3(new_n571), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n587), .A2(new_n572), .B1(new_n578), .B2(new_n579), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n234), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n585), .B2(new_n589), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n297), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT25), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n594), .A2(KEYINPUT25), .A3(new_n596), .A4(new_n297), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n567), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n594), .A2(new_n596), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n566), .A2(G902), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n510), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n351), .ZN(G3));
  INV_X1    g422(.A(new_n555), .ZN(new_n609));
  INV_X1    g423(.A(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n550), .B2(new_n297), .ZN(new_n611));
  INV_X1    g425(.A(new_n605), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n505), .A3(new_n509), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT91), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n392), .A2(new_n408), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT91), .B1(new_n413), .B2(new_n415), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n309), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n615), .B1(new_n392), .B2(new_n408), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n308), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n426), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n250), .A2(new_n252), .B1(new_n305), .B2(G475), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n288), .A2(new_n292), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n292), .A2(KEYINPUT92), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n288), .B(new_n292), .C1(KEYINPUT92), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(G478), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n294), .A2(new_n297), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n293), .B2(new_n294), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n622), .A2(new_n424), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n614), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n340), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  INV_X1    g452(.A(new_n620), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT91), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n308), .B1(new_n619), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n425), .B(new_n423), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n293), .B(new_n295), .Z(new_n643));
  XOR2_X1   g457(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n644));
  NAND3_X1  g458(.A1(new_n246), .A2(new_n247), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n247), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n236), .B2(new_n245), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n251), .A2(KEYINPUT94), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n643), .A2(new_n306), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n638), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n650), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n621), .A2(KEYINPUT95), .A3(new_n423), .A4(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n614), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT35), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  OR2_X1    g470(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n657));
  OR3_X1    g471(.A1(new_n585), .A2(new_n589), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n657), .B1(new_n585), .B2(new_n589), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n603), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n658), .A2(KEYINPUT96), .A3(new_n659), .A4(new_n603), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n601), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n609), .A2(new_n611), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n428), .A2(new_n666), .A3(new_n505), .A4(new_n509), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT97), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n667), .B(new_n669), .ZN(G12));
  AND2_X1   g484(.A1(new_n505), .A2(new_n509), .ZN(new_n671));
  INV_X1    g485(.A(new_n665), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n418), .A2(new_n673), .A3(G902), .A4(G953), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT98), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n420), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n650), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n621), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n671), .A2(new_n565), .A3(new_n672), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  OAI21_X1  g496(.A(new_n371), .B1(new_n516), .B2(new_n520), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n532), .B1(new_n537), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n297), .B1(new_n542), .B2(new_n684), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n555), .A2(new_n556), .B1(G472), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n554), .A3(new_n564), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n554), .A3(new_n689), .A4(new_n564), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n672), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n676), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n671), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n417), .B(new_n698), .Z(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n253), .A2(new_n306), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n643), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n700), .A2(new_n426), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n693), .A2(new_n696), .A3(new_n697), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n199), .B(KEYINPUT101), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G45));
  AND2_X1   g520(.A1(new_n565), .A2(new_n672), .ZN(new_n707));
  INV_X1    g521(.A(new_n631), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n701), .A2(new_n708), .A3(new_n676), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n671), .A3(new_n621), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  INV_X1    g526(.A(new_n633), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n498), .A2(new_n499), .A3(new_n297), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n499), .B1(new_n498), .B2(new_n297), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n508), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(new_n716), .A3(new_n565), .A4(new_n605), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND2_X1  g533(.A1(new_n498), .A2(new_n297), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n509), .A3(new_n500), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n606), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n651), .A2(new_n653), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NOR3_X1   g540(.A1(new_n701), .A2(new_n643), .A3(new_n424), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n565), .A2(new_n727), .A3(new_n672), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n509), .A2(new_n721), .A3(new_n500), .A4(new_n621), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(new_n551), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n543), .B1(new_n560), .B2(new_n532), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n531), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n536), .A2(new_n539), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n536), .A2(KEYINPUT102), .A3(new_n539), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n530), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n732), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n611), .A2(new_n612), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n642), .A2(new_n702), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n716), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND2_X1  g558(.A1(new_n550), .A2(new_n297), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(G472), .ZN(new_n746));
  INV_X1    g560(.A(new_n740), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n672), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n740), .B1(new_n745), .B2(G472), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n672), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n729), .A3(new_n710), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n502), .B2(G469), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n495), .A2(new_n477), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n501), .A2(new_n475), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n756), .A2(new_n758), .A3(new_n759), .A4(G469), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n500), .A2(new_n761), .A3(new_n504), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n509), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT105), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n765), .A3(new_n509), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n409), .A2(new_n416), .A3(new_n425), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n409), .A2(new_n416), .A3(KEYINPUT106), .A4(new_n425), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n555), .A2(new_n556), .B1(G472), .B2(new_n562), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n612), .B(new_n709), .C1(new_n773), .C2(new_n552), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n764), .A2(new_n766), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT42), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n771), .B1(new_n763), .B2(KEYINPUT105), .ZN(new_n777));
  INV_X1    g591(.A(new_n606), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n766), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  INV_X1    g596(.A(new_n766), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n765), .B1(new_n762), .B2(new_n509), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n771), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(KEYINPUT107), .A3(new_n778), .A4(new_n678), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n777), .A2(new_n778), .A3(new_n678), .A4(new_n766), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT108), .B(G134), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G36));
  NOR3_X1   g606(.A1(new_n701), .A2(KEYINPUT43), .A3(new_n631), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT43), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n622), .B2(new_n708), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n746), .A2(new_n555), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n672), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n771), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n758), .A2(new_n759), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n499), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n805), .A2(KEYINPUT109), .B1(KEYINPUT45), .B2(new_n502), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(KEYINPUT109), .B2(new_n805), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n504), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n714), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n504), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n508), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n694), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n802), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n447), .ZN(G39));
  NOR4_X1   g630(.A1(new_n565), .A2(new_n605), .A3(new_n771), .A4(new_n709), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(KEYINPUT47), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n812), .B2(new_n508), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n210), .ZN(G42));
  NOR2_X1   g637(.A1(new_n722), .A2(new_n771), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n793), .A2(new_n420), .A3(new_n795), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n773), .A2(new_n552), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n605), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT48), .Z(new_n829));
  NAND2_X1  g643(.A1(new_n191), .A2(G952), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n825), .A2(new_n741), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n729), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n612), .A2(new_n420), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n692), .A2(new_n824), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n631), .B1(new_n253), .B2(new_n306), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n832), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n826), .A2(new_n753), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n622), .A2(new_n631), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n831), .A2(new_n426), .A3(new_n700), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n722), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n841), .A2(new_n844), .A3(new_n722), .ZN(new_n845));
  OAI221_X1 g659(.A(new_n839), .B1(new_n834), .B2(new_n840), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n714), .A2(new_n715), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n819), .B(new_n821), .C1(new_n509), .C2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n831), .A2(new_n772), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n838), .B1(new_n851), .B2(KEYINPUT51), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(KEYINPUT51), .B2(new_n851), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n751), .B1(new_n750), .B2(new_n672), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n611), .A2(new_n740), .A3(new_n665), .A4(KEYINPUT103), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n710), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n509), .A3(new_n621), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n565), .A2(new_n505), .A3(new_n509), .A4(new_n672), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n857), .A2(new_n858), .B1(new_n859), .B2(new_n679), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT114), .B1(new_n754), .B2(new_n681), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n676), .B(KEYINPUT115), .Z(new_n865));
  NAND4_X1  g679(.A1(new_n621), .A2(new_n643), .A3(new_n701), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n763), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n691), .A2(new_n867), .A3(new_n665), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n711), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n854), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n869), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n860), .A2(new_n861), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n754), .A2(new_n681), .A3(KEYINPUT114), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n874), .A3(KEYINPUT116), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n868), .A2(new_n711), .A3(new_n681), .A4(new_n754), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n870), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n296), .A2(new_n306), .A3(new_n649), .A4(new_n676), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n769), .A2(new_n880), .A3(new_n770), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n769), .A2(new_n880), .A3(KEYINPUT112), .A4(new_n770), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n707), .A3(new_n886), .A4(new_n671), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT113), .B1(new_n859), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n667), .B1(new_n510), .B2(new_n606), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n253), .A2(new_n643), .A3(new_n306), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n417), .A3(new_n427), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n835), .A2(KEYINPUT111), .A3(new_n417), .A4(new_n427), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n417), .A2(new_n427), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT111), .B1(new_n896), .B2(new_n835), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n614), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n777), .A2(new_n710), .A3(new_n753), .A4(new_n766), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n890), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n717), .A2(new_n725), .A3(new_n730), .A4(new_n743), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n790), .A3(new_n781), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n879), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n860), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n871), .A2(new_n907), .B1(new_n876), .B2(new_n877), .ZN(new_n908));
  XOR2_X1   g722(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n909));
  NOR3_X1   g723(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT54), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n904), .B2(new_n908), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n871), .A2(new_n874), .A3(KEYINPUT116), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT116), .B1(new_n871), .B2(new_n874), .ZN(new_n915));
  INV_X1    g729(.A(new_n878), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n890), .A2(new_n900), .A3(new_n901), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n789), .B2(new_n786), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n717), .A2(new_n743), .ZN(new_n920));
  AOI22_X1  g734(.A1(new_n723), .A2(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n776), .A2(new_n920), .A3(new_n921), .A4(new_n780), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT118), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n903), .A2(new_n924), .A3(new_n776), .A4(new_n780), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n919), .A2(KEYINPUT53), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n912), .B(new_n913), .C1(new_n917), .C2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n853), .A2(new_n911), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(G952), .B2(G953), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n612), .A2(new_n508), .A3(new_n426), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n622), .A3(new_n708), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n699), .B(new_n931), .C1(new_n848), .C2(KEYINPUT49), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(KEYINPUT49), .B2(new_n848), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n929), .B1(new_n691), .B2(new_n933), .ZN(G75));
  AND3_X1   g748(.A1(new_n902), .A2(KEYINPUT53), .A3(new_n790), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n922), .B(new_n924), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n879), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n297), .B1(new_n937), .B2(new_n913), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(KEYINPUT119), .A3(G210), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n411), .A2(new_n412), .A3(new_n410), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n392), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT119), .B1(new_n938), .B2(G210), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n191), .A2(G952), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n938), .B2(G210), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n943), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n946), .A2(new_n950), .ZN(G51));
  AOI211_X1 g765(.A(new_n297), .B(new_n807), .C1(new_n937), .C2(new_n913), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n504), .B(KEYINPUT57), .Z(new_n953));
  INV_X1    g767(.A(new_n927), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n912), .B1(new_n937), .B2(new_n913), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n498), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT120), .B1(new_n957), .B2(new_n947), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT120), .ZN(new_n959));
  INV_X1    g773(.A(new_n498), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n913), .B1(new_n917), .B2(new_n926), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT54), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n927), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(new_n953), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n959), .B(new_n948), .C1(new_n964), .C2(new_n952), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n958), .A2(new_n965), .ZN(G54));
  NAND3_X1  g780(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .ZN(new_n967));
  INV_X1    g781(.A(new_n246), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n947), .ZN(G60));
  XNOR2_X1  g785(.A(new_n629), .B(KEYINPUT59), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n911), .B2(new_n927), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n625), .A2(new_n627), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n948), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n625), .B2(new_n627), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n963), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  NAND4_X1  g796(.A1(new_n961), .A2(new_n658), .A3(new_n659), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n961), .A2(new_n982), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n948), .B(new_n983), .C1(new_n984), .C2(new_n602), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n985), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT61), .B1(new_n985), .B2(KEYINPUT122), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(G66));
  AOI21_X1  g802(.A(new_n191), .B1(new_n421), .B2(G224), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n903), .A2(new_n900), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n191), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n386), .B(new_n391), .C1(G898), .C2(new_n191), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n991), .B(new_n992), .Z(G69));
  NAND2_X1  g807(.A1(new_n827), .A2(new_n605), .ZN(new_n994));
  INV_X1    g808(.A(new_n621), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n994), .A2(new_n995), .A3(new_n702), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n814), .B1(new_n802), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n822), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n874), .A2(new_n711), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n999), .A2(new_n781), .A3(new_n790), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n191), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(G900), .B2(new_n191), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n545), .B(KEYINPUT123), .Z(new_n1004));
  NAND2_X1  g818(.A1(new_n238), .A2(new_n239), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G227), .A2(G900), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(G953), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n892), .A2(new_n835), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n695), .A2(new_n606), .A3(new_n771), .A4(new_n1010), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n815), .A2(new_n822), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1000), .A2(new_n704), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT124), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT124), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1012), .A2(new_n1014), .A3(new_n1018), .A4(new_n1015), .ZN(new_n1019));
  AOI21_X1  g833(.A(G953), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1007), .B(new_n1009), .C1(new_n1020), .C2(new_n1006), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1006), .ZN(new_n1022));
  OAI211_X1 g836(.A(G953), .B(new_n1008), .C1(new_n1003), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(G72));
  XNOR2_X1  g838(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n610), .A2(new_n297), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(new_n1001), .B2(new_n990), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n560), .B(KEYINPUT126), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1029), .A2(new_n532), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n947), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n906), .A2(new_n910), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n560), .A2(new_n532), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1027), .B1(new_n1033), .B2(new_n542), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1031), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1029), .A2(new_n532), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1017), .A2(new_n903), .A3(new_n900), .A4(new_n1019), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1036), .B1(new_n1037), .B2(new_n1027), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1035), .A2(new_n1038), .ZN(G57));
endmodule


