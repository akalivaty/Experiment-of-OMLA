

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n678), .B(KEYINPUT27), .ZN(n679) );
  XNOR2_X1 U552 ( .A(n680), .B(n679), .ZN(n682) );
  INV_X1 U553 ( .A(KEYINPUT28), .ZN(n683) );
  INV_X1 U554 ( .A(G168), .ZN(n712) );
  XNOR2_X1 U555 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n717) );
  NOR2_X1 U556 ( .A1(G2084), .A2(n726), .ZN(n676) );
  XNOR2_X1 U557 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U558 ( .A1(n674), .A2(G1384), .ZN(n774) );
  XNOR2_X1 U559 ( .A(n531), .B(KEYINPUT64), .ZN(n873) );
  NOR2_X1 U560 ( .A1(G651), .A2(n610), .ZN(n635) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n628) );
  NAND2_X1 U562 ( .A1(G89), .A2(n628), .ZN(n515) );
  XNOR2_X1 U563 ( .A(n515), .B(KEYINPUT72), .ZN(n516) );
  XNOR2_X1 U564 ( .A(n516), .B(KEYINPUT4), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n610) );
  INV_X1 U566 ( .A(G651), .ZN(n520) );
  NOR2_X1 U567 ( .A1(n610), .A2(n520), .ZN(n626) );
  NAND2_X1 U568 ( .A1(G76), .A2(n626), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U570 ( .A(n519), .B(KEYINPUT5), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n521), .Z(n629) );
  NAND2_X1 U573 ( .A1(G63), .A2(n629), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G51), .A2(n635), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(n527), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U579 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U580 ( .A(KEYINPUT85), .ZN(n530) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X2 U582 ( .A(KEYINPUT17), .B(n528), .Z(n876) );
  NAND2_X1 U583 ( .A1(G138), .A2(n876), .ZN(n529) );
  XOR2_X1 U584 ( .A(n530), .B(n529), .Z(n540) );
  INV_X1 U585 ( .A(KEYINPUT84), .ZN(n535) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U587 ( .A1(G114), .A2(n872), .ZN(n533) );
  INV_X1 U588 ( .A(G2105), .ZN(n536) );
  NOR2_X1 U589 ( .A1(n536), .A2(G2104), .ZN(n531) );
  NAND2_X1 U590 ( .A1(G126), .A2(n873), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n535), .B(n534), .ZN(n538) );
  AND2_X1 U593 ( .A1(n536), .A2(G2104), .ZN(n878) );
  NAND2_X1 U594 ( .A1(n878), .A2(G102), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n674) );
  BUF_X1 U597 ( .A(n674), .Z(G164) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  NAND2_X1 U600 ( .A1(G64), .A2(n629), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G52), .A2(n635), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G90), .A2(n628), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G77), .A2(n626), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  NOR2_X1 U607 ( .A1(n547), .A2(n546), .ZN(G171) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G7), .A2(G661), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n548), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U611 ( .A(G223), .ZN(n818) );
  NAND2_X1 U612 ( .A1(n818), .A2(G567), .ZN(n549) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(n549), .Z(G234) );
  NAND2_X1 U614 ( .A1(G81), .A2(n628), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT69), .B(n550), .Z(n551) );
  XNOR2_X1 U616 ( .A(n551), .B(KEYINPUT12), .ZN(n553) );
  NAND2_X1 U617 ( .A1(G68), .A2(n626), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(KEYINPUT13), .B(n554), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G56), .A2(n629), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n555), .Z(n558) );
  NAND2_X1 U622 ( .A1(n635), .A2(G43), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT70), .B(n556), .Z(n557) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n967) );
  INV_X1 U626 ( .A(G860), .ZN(n604) );
  OR2_X1 U627 ( .A1(n967), .A2(n604), .ZN(G153) );
  INV_X1 U628 ( .A(G171), .ZN(G301) );
  NAND2_X1 U629 ( .A1(G868), .A2(G301), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G66), .A2(n629), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G92), .A2(n628), .ZN(n562) );
  NAND2_X1 U632 ( .A1(G79), .A2(n626), .ZN(n561) );
  NAND2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U634 ( .A1(G54), .A2(n635), .ZN(n563) );
  XNOR2_X1 U635 ( .A(KEYINPUT71), .B(n563), .ZN(n564) );
  NOR2_X1 U636 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U638 ( .A(n568), .B(KEYINPUT15), .ZN(n970) );
  OR2_X1 U639 ( .A1(n970), .A2(G868), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(G284) );
  NAND2_X1 U641 ( .A1(G91), .A2(n628), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n571), .B(KEYINPUT66), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G78), .A2(n626), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G65), .A2(n629), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G53), .A2(n635), .ZN(n574) );
  XNOR2_X1 U647 ( .A(KEYINPUT67), .B(n574), .ZN(n575) );
  NOR2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G299) );
  INV_X1 U650 ( .A(G868), .ZN(n649) );
  NOR2_X1 U651 ( .A1(G286), .A2(n649), .ZN(n580) );
  NOR2_X1 U652 ( .A1(G868), .A2(G299), .ZN(n579) );
  NOR2_X1 U653 ( .A1(n580), .A2(n579), .ZN(G297) );
  NAND2_X1 U654 ( .A1(n604), .A2(G559), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n581), .A2(n970), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n582), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U657 ( .A1(G868), .A2(n967), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G868), .A2(n970), .ZN(n583) );
  NOR2_X1 U659 ( .A1(G559), .A2(n583), .ZN(n584) );
  NOR2_X1 U660 ( .A1(n585), .A2(n584), .ZN(G282) );
  XNOR2_X1 U661 ( .A(G2100), .B(KEYINPUT75), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G99), .A2(n878), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G111), .A2(n872), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT74), .B(n588), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n873), .A2(G123), .ZN(n589) );
  XOR2_X1 U667 ( .A(KEYINPUT18), .B(n589), .Z(n590) );
  XNOR2_X1 U668 ( .A(n590), .B(KEYINPUT73), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G135), .A2(n876), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n921) );
  XNOR2_X1 U672 ( .A(n921), .B(G2096), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(G156) );
  NAND2_X1 U674 ( .A1(G93), .A2(n628), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G80), .A2(n626), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U677 ( .A1(G67), .A2(n629), .ZN(n600) );
  NAND2_X1 U678 ( .A1(G55), .A2(n635), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  OR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n648) );
  XNOR2_X1 U681 ( .A(n648), .B(KEYINPUT76), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G559), .A2(n970), .ZN(n603) );
  XOR2_X1 U683 ( .A(n967), .B(n603), .Z(n646) );
  NAND2_X1 U684 ( .A1(n646), .A2(n604), .ZN(n605) );
  XNOR2_X1 U685 ( .A(n606), .B(n605), .ZN(G145) );
  NAND2_X1 U686 ( .A1(G49), .A2(n635), .ZN(n608) );
  NAND2_X1 U687 ( .A1(G74), .A2(G651), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n629), .A2(n609), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n610), .A2(G87), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(G288) );
  NAND2_X1 U692 ( .A1(G88), .A2(n628), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G75), .A2(n626), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G62), .A2(n629), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G50), .A2(n635), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(G166) );
  NAND2_X1 U699 ( .A1(G60), .A2(n629), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G47), .A2(n635), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G85), .A2(n628), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G72), .A2(n626), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n625), .B(KEYINPUT65), .ZN(G290) );
  NAND2_X1 U707 ( .A1(G73), .A2(n626), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n627), .Z(n634) );
  NAND2_X1 U709 ( .A1(G86), .A2(n628), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G61), .A2(n629), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U712 ( .A(KEYINPUT77), .B(n632), .Z(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n635), .A2(G48), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(G305) );
  XOR2_X1 U716 ( .A(KEYINPUT78), .B(KEYINPUT19), .Z(n639) );
  XNOR2_X1 U717 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U719 ( .A(G166), .B(n640), .ZN(n642) );
  INV_X1 U720 ( .A(G299), .ZN(n686) );
  XNOR2_X1 U721 ( .A(G290), .B(n686), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n648), .B(n643), .ZN(n644) );
  XNOR2_X1 U724 ( .A(G288), .B(n644), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(G305), .ZN(n889) );
  XNOR2_X1 U726 ( .A(n646), .B(n889), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n647), .A2(G868), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(G295) );
  NAND2_X1 U730 ( .A1(G2078), .A2(G2084), .ZN(n652) );
  XOR2_X1 U731 ( .A(KEYINPUT20), .B(n652), .Z(n653) );
  NAND2_X1 U732 ( .A1(G2090), .A2(n653), .ZN(n654) );
  XNOR2_X1 U733 ( .A(KEYINPUT21), .B(n654), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n655), .A2(G2072), .ZN(G158) );
  XOR2_X1 U735 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  XNOR2_X1 U736 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U737 ( .A1(G219), .A2(G220), .ZN(n656) );
  XNOR2_X1 U738 ( .A(KEYINPUT22), .B(n656), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n657), .A2(G96), .ZN(n658) );
  NOR2_X1 U740 ( .A1(n658), .A2(G218), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n659), .B(KEYINPUT81), .ZN(n910) );
  NAND2_X1 U742 ( .A1(n910), .A2(G2106), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G120), .A2(G108), .ZN(n660) );
  NOR2_X1 U744 ( .A1(G237), .A2(n660), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n661), .A2(G69), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(KEYINPUT82), .ZN(n909) );
  NAND2_X1 U747 ( .A1(G567), .A2(n909), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n664), .A2(n663), .ZN(n822) );
  NAND2_X1 U749 ( .A1(G661), .A2(G483), .ZN(n665) );
  XOR2_X1 U750 ( .A(KEYINPUT83), .B(n665), .Z(n666) );
  NOR2_X1 U751 ( .A1(n822), .A2(n666), .ZN(n821) );
  NAND2_X1 U752 ( .A1(n821), .A2(G36), .ZN(G176) );
  NAND2_X1 U753 ( .A1(n872), .A2(G113), .ZN(n669) );
  NAND2_X1 U754 ( .A1(G101), .A2(n878), .ZN(n667) );
  XOR2_X1 U755 ( .A(KEYINPUT23), .B(n667), .Z(n668) );
  NAND2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G137), .A2(n876), .ZN(n671) );
  NAND2_X1 U758 ( .A1(G125), .A2(n873), .ZN(n670) );
  NAND2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U760 ( .A1(n673), .A2(n672), .ZN(G160) );
  INV_X1 U761 ( .A(G166), .ZN(G303) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n775) );
  INV_X1 U763 ( .A(n775), .ZN(n675) );
  NAND2_X2 U764 ( .A1(n675), .A2(n774), .ZN(n726) );
  XOR2_X1 U765 ( .A(KEYINPUT92), .B(n676), .Z(n709) );
  INV_X1 U766 ( .A(n709), .ZN(n677) );
  NAND2_X1 U767 ( .A1(n677), .A2(G8), .ZN(n724) );
  NAND2_X1 U768 ( .A1(G8), .A2(n726), .ZN(n758) );
  NOR2_X1 U769 ( .A1(G1966), .A2(n758), .ZN(n722) );
  INV_X1 U770 ( .A(n726), .ZN(n692) );
  NAND2_X1 U771 ( .A1(G2072), .A2(n692), .ZN(n680) );
  INV_X1 U772 ( .A(KEYINPUT93), .ZN(n678) );
  INV_X1 U773 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U774 ( .A1(n692), .A2(n998), .ZN(n681) );
  NOR2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n685) );
  NOR2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n684) );
  XNOR2_X1 U777 ( .A(n684), .B(n683), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n701) );
  INV_X1 U779 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U780 ( .A1(n726), .A2(n942), .ZN(n687) );
  XOR2_X1 U781 ( .A(n687), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U782 ( .A1(n726), .A2(G1341), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n967), .A2(n690), .ZN(n691) );
  OR2_X1 U785 ( .A1(n970), .A2(n691), .ZN(n699) );
  NAND2_X1 U786 ( .A1(n970), .A2(n691), .ZN(n697) );
  AND2_X1 U787 ( .A1(n692), .A2(G2067), .ZN(n693) );
  XOR2_X1 U788 ( .A(n693), .B(KEYINPUT94), .Z(n695) );
  NAND2_X1 U789 ( .A1(n726), .A2(G1348), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U795 ( .A(KEYINPUT29), .B(n704), .Z(n708) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NOR2_X1 U797 ( .A1(n726), .A2(n943), .ZN(n706) );
  AND2_X1 U798 ( .A1(n726), .A2(G1961), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n714) );
  NAND2_X1 U800 ( .A1(G171), .A2(n714), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n720) );
  NAND2_X1 U802 ( .A1(G8), .A2(n709), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n722), .A2(n710), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n711), .B(KEYINPUT30), .ZN(n713) );
  AND2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U806 ( .A1(G171), .A2(n714), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n725) );
  INV_X1 U809 ( .A(n725), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U811 ( .A1(n724), .A2(n723), .ZN(n750) );
  NAND2_X1 U812 ( .A1(G1976), .A2(G288), .ZN(n972) );
  AND2_X1 U813 ( .A1(n750), .A2(n972), .ZN(n736) );
  NAND2_X1 U814 ( .A1(n725), .A2(G286), .ZN(n734) );
  INV_X1 U815 ( .A(G8), .ZN(n732) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n758), .ZN(n728) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n726), .ZN(n727) );
  NOR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n729), .A2(G303), .ZN(n730) );
  XNOR2_X1 U820 ( .A(n730), .B(KEYINPUT96), .ZN(n731) );
  OR2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  AND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U823 ( .A(n735), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n736), .A2(n749), .ZN(n741) );
  INV_X1 U825 ( .A(n972), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n743) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n737) );
  NOR2_X1 U828 ( .A1(n743), .A2(n737), .ZN(n976) );
  OR2_X1 U829 ( .A1(n738), .A2(n976), .ZN(n739) );
  OR2_X1 U830 ( .A1(n758), .A2(n739), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U832 ( .A1(KEYINPUT33), .A2(n742), .ZN(n748) );
  XOR2_X1 U833 ( .A(G1981), .B(G305), .Z(n964) );
  INV_X1 U834 ( .A(n964), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n743), .A2(KEYINPUT33), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n758), .A2(n744), .ZN(n745) );
  NOR2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n762) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n753) );
  NOR2_X1 U840 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U841 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n754), .A2(n758), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n755), .B(KEYINPUT91), .ZN(n756) );
  XNOR2_X1 U846 ( .A(n756), .B(KEYINPUT24), .ZN(n757) );
  OR2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n778) );
  NAND2_X1 U850 ( .A1(G104), .A2(n878), .ZN(n764) );
  NAND2_X1 U851 ( .A1(G140), .A2(n876), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n766) );
  XOR2_X1 U853 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n765) );
  XNOR2_X1 U854 ( .A(n766), .B(n765), .ZN(n771) );
  NAND2_X1 U855 ( .A1(G116), .A2(n872), .ZN(n768) );
  NAND2_X1 U856 ( .A1(G128), .A2(n873), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U858 ( .A(KEYINPUT35), .B(n769), .Z(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(n772), .B(KEYINPUT36), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(KEYINPUT88), .ZN(n887) );
  XNOR2_X1 U862 ( .A(KEYINPUT37), .B(G2067), .ZN(n810) );
  NOR2_X1 U863 ( .A1(n887), .A2(n810), .ZN(n917) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U865 ( .A(n776), .B(KEYINPUT86), .ZN(n813) );
  NAND2_X1 U866 ( .A1(n917), .A2(n813), .ZN(n777) );
  XNOR2_X1 U867 ( .A(n777), .B(KEYINPUT89), .ZN(n807) );
  NOR2_X1 U868 ( .A1(n778), .A2(n807), .ZN(n797) );
  INV_X1 U869 ( .A(n813), .ZN(n779) );
  XOR2_X1 U870 ( .A(G1986), .B(G290), .Z(n969) );
  OR2_X1 U871 ( .A1(n779), .A2(n969), .ZN(n795) );
  NAND2_X1 U872 ( .A1(G95), .A2(n878), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G131), .A2(n876), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G107), .A2(n872), .ZN(n783) );
  NAND2_X1 U876 ( .A1(G119), .A2(n873), .ZN(n782) );
  NAND2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n784) );
  OR2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n856) );
  XNOR2_X1 U879 ( .A(KEYINPUT90), .B(G1991), .ZN(n951) );
  NAND2_X1 U880 ( .A1(n856), .A2(n951), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G117), .A2(n872), .ZN(n787) );
  NAND2_X1 U882 ( .A1(G141), .A2(n876), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n878), .A2(G105), .ZN(n788) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G129), .A2(n873), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n855) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n855), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n916) );
  NAND2_X1 U891 ( .A1(n813), .A2(n916), .ZN(n799) );
  AND2_X1 U892 ( .A1(n795), .A2(n799), .ZN(n796) );
  AND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U894 ( .A(n798), .B(KEYINPUT97), .ZN(n816) );
  INV_X1 U895 ( .A(n799), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n856), .A2(n951), .ZN(n920) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n920), .A2(n800), .ZN(n801) );
  NOR2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n855), .A2(G1996), .ZN(n803) );
  XNOR2_X1 U901 ( .A(n803), .B(KEYINPUT98), .ZN(n914) );
  NOR2_X1 U902 ( .A1(n804), .A2(n914), .ZN(n805) );
  XOR2_X1 U903 ( .A(n805), .B(KEYINPUT39), .Z(n806) );
  XNOR2_X1 U904 ( .A(KEYINPUT99), .B(n806), .ZN(n809) );
  INV_X1 U905 ( .A(n807), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n810), .A2(n887), .ZN(n811) );
  XNOR2_X1 U908 ( .A(n811), .B(KEYINPUT100), .ZN(n936) );
  NAND2_X1 U909 ( .A1(n812), .A2(n936), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U912 ( .A(n817), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U915 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(G188) );
  INV_X1 U918 ( .A(n822), .ZN(G319) );
  XNOR2_X1 U919 ( .A(G2067), .B(G2078), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(G2678), .ZN(n833) );
  XOR2_X1 U921 ( .A(KEYINPUT42), .B(KEYINPUT103), .Z(n825) );
  XNOR2_X1 U922 ( .A(KEYINPUT104), .B(G2100), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U924 ( .A(G2096), .B(G2090), .Z(n827) );
  XNOR2_X1 U925 ( .A(G2072), .B(G2084), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U927 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U928 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(G227) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(G2474), .Z(n838) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n846) );
  XOR2_X1 U937 ( .A(G1976), .B(G1981), .Z(n840) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1971), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT108), .B(G1956), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1961), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U945 ( .A1(G112), .A2(n872), .ZN(n848) );
  NAND2_X1 U946 ( .A1(G136), .A2(n876), .ZN(n847) );
  NAND2_X1 U947 ( .A1(n848), .A2(n847), .ZN(n854) );
  NAND2_X1 U948 ( .A1(n873), .A2(G124), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n849), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G100), .A2(n878), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n850), .B(KEYINPUT110), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(G162) );
  XNOR2_X1 U954 ( .A(n921), .B(n855), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n858), .B(KEYINPUT46), .Z(n860) );
  XNOR2_X1 U957 ( .A(G160), .B(KEYINPUT48), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n861), .B(G162), .Z(n871) );
  NAND2_X1 U960 ( .A1(G103), .A2(n878), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G139), .A2(n876), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT112), .B(n864), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G115), .A2(n872), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G127), .A2(n873), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n867), .Z(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n927) );
  XNOR2_X1 U969 ( .A(G164), .B(n927), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n885) );
  NAND2_X1 U971 ( .A1(G118), .A2(n872), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G130), .A2(n873), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n883) );
  NAND2_X1 U974 ( .A1(n876), .A2(G142), .ZN(n877) );
  XOR2_X1 U975 ( .A(KEYINPUT111), .B(n877), .Z(n880) );
  NAND2_X1 U976 ( .A1(n878), .A2(G106), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U978 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(n885), .B(n884), .Z(n886) );
  XOR2_X1 U981 ( .A(n887), .B(n886), .Z(n888) );
  NOR2_X1 U982 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U983 ( .A(n967), .B(n889), .ZN(n891) );
  XNOR2_X1 U984 ( .A(G171), .B(n970), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n892), .B(G286), .ZN(n893) );
  NOR2_X1 U987 ( .A1(G37), .A2(n893), .ZN(G397) );
  XOR2_X1 U988 ( .A(G2454), .B(G2435), .Z(n895) );
  XNOR2_X1 U989 ( .A(G2438), .B(G2427), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n902) );
  XOR2_X1 U991 ( .A(KEYINPUT101), .B(G2446), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2443), .B(G2430), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n898), .B(G2451), .Z(n900) );
  XNOR2_X1 U995 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  NAND2_X1 U998 ( .A1(n903), .A2(G14), .ZN(n912) );
  NAND2_X1 U999 ( .A1(G319), .A2(n912), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(G225) );
  XNOR2_X1 U1005 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  XOR2_X1 U1006 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U1008 ( .A(G120), .ZN(G236) );
  INV_X1 U1009 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(KEYINPUT102), .ZN(G325) );
  INV_X1 U1012 ( .A(G325), .ZN(G261) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  INV_X1 U1014 ( .A(n912), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n915), .Z(n926) );
  XNOR2_X1 U1018 ( .A(G160), .B(G2084), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT115), .B(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n934) );
  XNOR2_X1 U1025 ( .A(G164), .B(G2078), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(G2072), .B(n927), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(n928), .B(KEYINPUT116), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT117), .ZN(n932) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n932), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(G29), .ZN(n1021) );
  XOR2_X1 U1035 ( .A(G2090), .B(G35), .Z(n941) );
  XOR2_X1 U1036 ( .A(G34), .B(KEYINPUT54), .Z(n939) );
  XNOR2_X1 U1037 ( .A(n939), .B(G2084), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n959) );
  XNOR2_X1 U1039 ( .A(G32), .B(n942), .ZN(n950) );
  XOR2_X1 U1040 ( .A(n943), .B(G27), .Z(n948) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(KEYINPUT119), .B(n946), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n955) );
  XOR2_X1 U1047 ( .A(G25), .B(n951), .Z(n952) );
  NAND2_X1 U1048 ( .A1(n952), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(KEYINPUT118), .B(n953), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT120), .B(n957), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(KEYINPUT121), .B(n960), .Z(n961) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n962), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(G11), .ZN(n1019) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n986) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT57), .ZN(n984) );
  XOR2_X1 U1062 ( .A(G1341), .B(n967), .Z(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n982) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n970), .ZN(n980) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G299), .B(G1956), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n1017) );
  INV_X1 U1076 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1077 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1013) );
  XOR2_X1 U1078 ( .A(G1971), .B(G22), .Z(n989) );
  XOR2_X1 U1079 ( .A(G23), .B(KEYINPUT124), .Z(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(G1976), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1082 ( .A(KEYINPUT125), .B(G1986), .Z(n990) );
  XNOR2_X1 U1083 ( .A(G24), .B(n990), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(KEYINPUT126), .B(n993), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n994), .B(KEYINPUT58), .ZN(n1011) );
  XNOR2_X1 U1087 ( .A(G1961), .B(G5), .ZN(n1009) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT122), .B(n997), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n998), .B(G20), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT59), .B(G1348), .Z(n1001) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1004), .Z(n1006) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(KEYINPUT123), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

