//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT65), .Z(new_n461));
  AND2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT66), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(KEYINPUT67), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n467), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n464), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  INV_X1    g057(.A(new_n479), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n483), .A2(G136), .B1(G124), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G100), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n486), .A2(new_n464), .A3(KEYINPUT68), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT68), .B1(new_n486), .B2(new_n464), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT69), .Z(G162));
  OAI211_X1 g066(.A(KEYINPUT4), .B(G138), .C1(new_n469), .C2(new_n470), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n478), .B2(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n497), .B2(new_n464), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n467), .A2(new_n471), .A3(G138), .A4(new_n464), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G50), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n507), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(new_n503), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n504), .A2(new_n505), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n506), .B(KEYINPUT70), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n526), .B1(G51), .B2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n515), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n513), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G651), .B1(G90), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n527), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n527), .A2(G43), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n530), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(G81), .B2(new_n533), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G860), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT71), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n530), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(G91), .B2(new_n533), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n506), .A2(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n506), .A2(new_n559), .A3(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(new_n527), .A2(G51), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n563), .A2(new_n525), .A3(new_n523), .ZN(G286));
  OR2_X1    g139(.A1(new_n514), .A2(new_n517), .ZN(G303));
  NAND2_X1  g140(.A1(new_n533), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n506), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n513), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n519), .A2(new_n515), .A3(KEYINPUT72), .A4(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n510), .B2(new_n509), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G48), .B2(new_n506), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n530), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G85), .B2(new_n533), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n535), .B2(new_n584), .ZN(G290));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(G301), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n527), .A2(KEYINPUT73), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n527), .A2(KEYINPUT73), .ZN(new_n589));
  OAI21_X1  g164(.A(G54), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n513), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n530), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n591), .A2(new_n594), .B1(new_n597), .B2(G651), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(new_n586), .ZN(G284));
  AOI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(new_n586), .ZN(G321));
  MUX2_X1   g176(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n599), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(new_n544), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n586), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n604), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n586), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT11), .Z(G282));
  INV_X1    g185(.A(new_n609), .ZN(G323));
  AND2_X1   g186(.A1(new_n467), .A2(new_n471), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n476), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT13), .B(G2100), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n484), .A2(G123), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  AND2_X1   g195(.A1(G111), .A2(G2105), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G99), .B2(new_n464), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n619), .B1(new_n620), .B2(new_n479), .C1(new_n475), .C2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G2096), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n617), .A2(new_n618), .A3(new_n625), .ZN(G156));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2427), .ZN(new_n630));
  INV_X1    g205(.A(G2430), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT75), .Z(new_n644));
  NOR2_X1   g219(.A1(G2072), .A2(G2078), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n444), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(KEYINPUT17), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n649), .C1(new_n644), .C2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n644), .A3(new_n648), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n648), .B(new_n643), .C1(new_n444), .C2(new_n645), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n624), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(G227));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT76), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n661), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n664), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n662), .A2(new_n664), .A3(new_n668), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT78), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  INV_X1    g258(.A(G288), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT81), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT33), .B(G1976), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT32), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(G16), .A2(G22), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G166), .B2(G16), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1971), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n697));
  MUX2_X1   g272(.A(G24), .B(G290), .S(G16), .Z(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G1986), .ZN(new_n699));
  INV_X1    g274(.A(G25), .ZN(new_n700));
  OAI21_X1  g275(.A(KEYINPUT79), .B1(new_n700), .B2(G29), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n700), .A2(KEYINPUT79), .A3(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n483), .A2(G131), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n484), .A2(G119), .ZN(new_n704));
  MUX2_X1   g279(.A(G95), .B(G107), .S(G2105), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G2104), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n701), .B(new_n702), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT80), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n698), .A2(G1986), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n699), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n696), .A2(new_n697), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT36), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n623), .A2(new_n709), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT88), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT31), .B(G11), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT30), .B(G28), .Z(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(G168), .A2(new_n682), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n682), .B2(G21), .ZN(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n719), .B(new_n722), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  NOR2_X1   g302(.A1(G171), .A2(new_n682), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G5), .B2(new_n682), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(new_n725), .C2(new_n724), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n682), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT23), .Z(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT89), .B(G1956), .Z(new_n734));
  AOI22_X1  g309(.A1(new_n729), .A2(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(G4), .A2(G16), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n599), .B2(G16), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT82), .B(G1348), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT83), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n730), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G35), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G162), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT29), .ZN(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n709), .A2(G32), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n483), .A2(G141), .B1(G129), .B2(new_n484), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G105), .B2(new_n476), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT87), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT87), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n748), .B1(new_n759), .B2(new_n709), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G27), .A2(G29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G164), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(new_n443), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n709), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G160), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n709), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n762), .A2(new_n765), .A3(new_n772), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n760), .A2(new_n761), .B1(new_n771), .B2(new_n770), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n606), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1341), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n709), .A2(G26), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT28), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n483), .A2(G140), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT84), .ZN(new_n781));
  MUX2_X1   g356(.A(G104), .B(G116), .S(G2105), .Z(new_n782));
  AOI22_X1  g357(.A1(G128), .A2(new_n484), .B1(new_n782), .B2(G2104), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n779), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT85), .B(G2067), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n773), .A2(new_n774), .A3(new_n777), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n709), .A2(G33), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n612), .A2(G127), .ZN(new_n790));
  INV_X1    g365(.A(G115), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n475), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n464), .B1(new_n792), .B2(KEYINPUT86), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(KEYINPUT86), .B2(new_n792), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n476), .A2(G103), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT25), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n796), .A2(new_n797), .B1(G139), .B2(new_n483), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(new_n709), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(new_n442), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n742), .A2(new_n747), .A3(new_n788), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n717), .A2(new_n802), .ZN(G150));
  INV_X1    g378(.A(G150), .ZN(G311));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  INV_X1    g380(.A(G67), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n530), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n503), .B1(new_n807), .B2(KEYINPUT90), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(KEYINPUT90), .B2(new_n807), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT91), .B(G93), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n527), .A2(G55), .B1(new_n533), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT37), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n812), .B(new_n544), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT38), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n598), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n604), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n545), .B1(new_n821), .B2(KEYINPUT39), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n815), .B1(new_n822), .B2(new_n823), .ZN(G145));
  NAND2_X1  g399(.A1(new_n483), .A2(G142), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  MUX2_X1   g402(.A(G106), .B(G118), .S(G2105), .Z(new_n828));
  AOI22_X1  g403(.A1(G130), .A2(new_n484), .B1(new_n828), .B2(G2104), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n707), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n615), .ZN(new_n832));
  OAI21_X1  g407(.A(G126), .B1(new_n469), .B2(new_n470), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n464), .B1(new_n833), .B2(new_n495), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT4), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n499), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n494), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n758), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n832), .B(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n799), .B(new_n784), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(G162), .B(new_n769), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n623), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(G37), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g423(.A(new_n608), .B(new_n816), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n599), .A2(G299), .ZN(new_n850));
  INV_X1    g425(.A(G299), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT94), .B1(new_n818), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n599), .A2(new_n853), .A3(G299), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n850), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G290), .B(G288), .ZN(new_n857));
  XNOR2_X1  g432(.A(G166), .B(G305), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT42), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n855), .A2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n856), .B(new_n860), .C1(new_n865), .C2(new_n849), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n856), .B1(new_n865), .B2(new_n849), .ZN(new_n870));
  INV_X1    g445(.A(new_n860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G868), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(KEYINPUT96), .A3(G868), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n812), .A2(new_n586), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G295));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G331));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n881));
  INV_X1    g456(.A(new_n864), .ZN(new_n882));
  XNOR2_X1  g457(.A(G286), .B(G301), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n816), .B(new_n883), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n885), .A3(new_n862), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT98), .ZN(new_n887));
  INV_X1    g462(.A(new_n855), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n882), .A2(new_n885), .A3(new_n890), .A4(new_n862), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n859), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  INV_X1    g469(.A(new_n859), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n887), .A2(new_n895), .A3(new_n889), .A4(new_n891), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT97), .B(KEYINPUT43), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n893), .A2(new_n894), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n886), .A2(new_n889), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n859), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n894), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n881), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n897), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n893), .A2(new_n894), .A3(new_n896), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n897), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT44), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n903), .A2(new_n907), .ZN(G397));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G164), .B2(G1384), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n472), .A2(new_n473), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G2105), .ZN(new_n912));
  INV_X1    g487(.A(new_n481), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(G40), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(G1996), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT46), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n784), .B(G2067), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n919), .B2(new_n758), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT127), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n708), .A2(new_n711), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n919), .B1(G1996), .B2(new_n758), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(G1996), .B2(new_n758), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n927), .B2(new_n915), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n784), .A2(G2067), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n928), .A2(KEYINPUT125), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT125), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n915), .A3(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n707), .B(new_n711), .Z(new_n933));
  OAI21_X1  g508(.A(new_n915), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(G290), .A2(G1986), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n916), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n937), .A2(KEYINPUT48), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(KEYINPUT48), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n924), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT102), .B(G8), .Z(new_n942));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(G164), .B2(G1384), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n838), .A2(KEYINPUT50), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n474), .A2(new_n948), .A3(new_n481), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT108), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n951), .B(new_n914), .C1(new_n944), .C2(new_n946), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n746), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n836), .B2(new_n837), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n910), .A2(new_n955), .A3(new_n949), .ZN(new_n956));
  INV_X1    g531(.A(G1971), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n942), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT100), .B(KEYINPUT55), .Z(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(G303), .A2(G8), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(G166), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT109), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n968));
  INV_X1    g543(.A(new_n958), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n970));
  AOI211_X1 g545(.A(new_n943), .B(G1384), .C1(new_n836), .C2(new_n837), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n949), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n951), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n914), .B1(new_n944), .B2(new_n946), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n969), .B1(new_n976), .B2(new_n746), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n968), .B(new_n965), .C1(new_n977), .C2(new_n942), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n967), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n965), .B(KEYINPUT101), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n746), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n963), .B1(new_n981), .B2(new_n958), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  INV_X1    g560(.A(G1981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n574), .A2(new_n986), .A3(new_n578), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n506), .A2(G48), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n519), .A2(new_n515), .A3(G86), .ZN(new_n989));
  INV_X1    g564(.A(new_n576), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n515), .B2(G61), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n988), .B(new_n989), .C1(new_n991), .C2(new_n503), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n993), .A3(G1981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n992), .B2(G1981), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n996), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n994), .A4(new_n987), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n942), .B1(new_n949), .B2(new_n954), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(new_n999), .A3(KEYINPUT105), .A4(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n684), .A2(G1976), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(KEYINPUT103), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(KEYINPUT103), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1000), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  NAND3_X1  g587(.A1(G288), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1005), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1005), .A2(KEYINPUT110), .A3(new_n1014), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n984), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n771), .A2(new_n974), .B1(new_n956), .B2(new_n725), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1020), .A2(G286), .A3(new_n942), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n979), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1003), .A2(new_n1004), .B1(new_n1025), .B2(new_n1009), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n746), .A2(new_n974), .B1(new_n956), .B2(new_n957), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n965), .B1(new_n1028), .B2(new_n963), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n983), .A2(new_n1021), .A3(KEYINPUT63), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1024), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(G1976), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT107), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1005), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n987), .B(KEYINPUT106), .Z(new_n1039));
  OAI21_X1  g614(.A(new_n1000), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n984), .A2(new_n1026), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1033), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1042), .ZN(new_n1047));
  INV_X1    g622(.A(new_n942), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G286), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1020), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n1020), .B2(new_n942), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  AOI211_X1 g627(.A(G2084), .B(new_n914), .C1(new_n944), .C2(new_n946), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n914), .B1(KEYINPUT45), .B2(new_n954), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1966), .B1(new_n1054), .B2(new_n910), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1052), .B(new_n1048), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1049), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1051), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n956), .A2(new_n725), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n947), .A2(new_n771), .A3(new_n949), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n963), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1049), .B(KEYINPUT119), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT121), .B(new_n1050), .C1(new_n1059), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1052), .B1(new_n1069), .B2(new_n1048), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1065), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1050), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1067), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT123), .B(G1961), .Z(new_n1075));
  NAND4_X1  g650(.A1(new_n910), .A2(new_n955), .A3(new_n443), .A4(new_n949), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n972), .A2(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI21_X1  g654(.A(G301), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n979), .A2(new_n1019), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1058), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n942), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n1052), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1063), .B1(new_n1020), .B2(new_n963), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1084), .A2(new_n1051), .B1(new_n1085), .B2(KEYINPUT51), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT121), .B1(new_n1086), .B2(new_n1050), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1071), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1074), .A2(new_n1081), .A3(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1092));
  AOI211_X1 g667(.A(new_n1077), .B(G2078), .C1(new_n954), .C2(KEYINPUT45), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1093), .A2(new_n910), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n972), .A2(new_n1075), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1098));
  AND4_X1   g673(.A1(G301), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1092), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1078), .B2(new_n1096), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1078), .A2(new_n1079), .A3(G301), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT54), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n974), .A2(G1956), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT114), .B1(new_n558), .B2(new_n560), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n558), .A2(KEYINPUT114), .A3(new_n560), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n556), .A3(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT115), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n556), .A2(new_n1109), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT115), .B(new_n1111), .C1(new_n1113), .C2(new_n1107), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1106), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1054), .A2(new_n910), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1105), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n974), .B2(G1956), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1120), .A2(KEYINPUT116), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(KEYINPUT116), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n1106), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1121), .A2(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G2067), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n949), .A2(new_n954), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n972), .A2(new_n739), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n818), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1119), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1116), .B1(new_n1105), .B2(new_n1118), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1119), .B1(new_n1132), .B2(KEYINPUT61), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1105), .A2(new_n1116), .A3(new_n1134), .A4(new_n1118), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n818), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n818), .B1(new_n1129), .B2(KEYINPUT60), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(KEYINPUT60), .B2(new_n1129), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT58), .B(G1341), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n956), .A2(G1996), .B1(new_n1128), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n606), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1143), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n606), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1133), .A2(new_n1137), .A3(new_n1139), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1104), .B1(new_n1131), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n979), .A2(new_n1019), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1091), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1044), .A2(new_n1047), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n916), .B1(new_n1155), .B2(new_n936), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT99), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n934), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n941), .B1(new_n1154), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g734(.A(new_n462), .ZN(new_n1161));
  NOR3_X1   g735(.A1(G227), .A2(G401), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n680), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1163), .B1(new_n845), .B2(new_n846), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n1164), .A2(new_n906), .A3(new_n905), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


