//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(new_n188), .A3(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n190), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(G137), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n195), .B2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(new_n196), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .A3(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n211), .A2(new_n212), .A3(new_n217), .A4(G128), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n215), .B2(new_n218), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n207), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT64), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n222), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n224), .A2(new_n227), .B1(new_n213), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n201), .A2(new_n203), .A3(new_n196), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n205), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n221), .A2(KEYINPUT30), .A3(new_n234), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n225), .A2(G128), .B1(new_n217), .B2(new_n212), .ZN(new_n236));
  INV_X1    g050(.A(new_n218), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n206), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n229), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n226), .B1(new_n225), .B2(new_n222), .ZN(new_n241));
  AND4_X1   g055(.A1(new_n226), .A2(new_n211), .A3(new_n212), .A4(new_n222), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(new_n232), .B2(new_n205), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n239), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n194), .B(new_n235), .C1(new_n247), .C2(KEYINPUT30), .ZN(new_n248));
  INV_X1    g062(.A(new_n194), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n221), .A2(new_n249), .A3(new_n234), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n250), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT31), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n233), .B1(new_n230), .B2(KEYINPUT65), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n243), .A2(new_n244), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n194), .B1(new_n260), .B2(new_n239), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n221), .A2(KEYINPUT28), .A3(new_n249), .A4(new_n234), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n255), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT31), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n248), .A2(new_n268), .A3(new_n250), .A4(new_n255), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n257), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n257), .A2(new_n272), .A3(new_n267), .A4(new_n269), .ZN(new_n273));
  NOR2_X1   g087(.A1(G472), .A2(G902), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n271), .A2(KEYINPUT32), .A3(new_n273), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n248), .A2(new_n250), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n266), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n282), .A3(new_n266), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n263), .A2(new_n264), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n261), .A4(new_n255), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n261), .A2(new_n263), .A3(new_n264), .A4(new_n255), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n287), .B2(KEYINPUT69), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n281), .A2(new_n283), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n221), .A2(new_n234), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n194), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n284), .A2(KEYINPUT29), .A3(new_n255), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT71), .B1(new_n296), .B2(G472), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n298));
  INV_X1    g112(.A(G472), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n298), .B(new_n299), .C1(new_n289), .C2(new_n295), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n277), .B(new_n278), .C1(new_n297), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G140), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n305), .A3(new_n210), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT76), .A2(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(KEYINPUT76), .A3(G125), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n306), .B1(new_n310), .B2(new_n210), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT86), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n306), .C1(new_n310), .C2(new_n210), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT18), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n204), .ZN(new_n320));
  INV_X1    g134(.A(new_n318), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT18), .B(G131), .C1(new_n321), .C2(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G131), .B1(new_n321), .B2(new_n316), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n204), .A3(new_n318), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n329), .A3(new_n327), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT16), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n305), .B2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n334), .A3(new_n304), .A4(G125), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n210), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n332), .A3(G146), .A4(new_n335), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n328), .A2(new_n330), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G113), .B(G122), .ZN(new_n340));
  INV_X1    g154(.A(G104), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n325), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n325), .B2(new_n339), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n293), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G475), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n347));
  NOR2_X1   g161(.A1(G475), .A2(G902), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT19), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n303), .A2(new_n305), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n310), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n338), .B1(new_n351), .B2(G146), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n326), .A2(new_n329), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT87), .B(new_n338), .C1(new_n351), .C2(G146), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n342), .B1(new_n357), .B2(new_n325), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n347), .B(new_n348), .C1(new_n358), .C2(new_n343), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n325), .A2(new_n339), .A3(new_n342), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n352), .A2(new_n353), .B1(new_n326), .B2(new_n329), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n362), .A2(new_n356), .B1(new_n315), .B2(new_n324), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(new_n342), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n347), .B1(new_n364), .B2(new_n348), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n346), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(G953), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G122), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G116), .ZN(new_n372));
  INV_X1    g186(.A(G116), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(G107), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n208), .A2(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n214), .A2(G143), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n195), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n214), .B2(G143), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(KEYINPUT88), .A3(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n378), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT89), .A4(new_n378), .ZN(new_n389));
  INV_X1    g203(.A(new_n377), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n380), .B1(new_n392), .B2(G134), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n375), .A2(new_n394), .A3(G107), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n372), .B(new_n374), .C1(KEYINPUT14), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n379), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n195), .B1(new_n377), .B2(new_n378), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n395), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n370), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n386), .A2(new_n387), .B1(KEYINPUT13), .B2(new_n390), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n195), .B1(new_n403), .B2(new_n389), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n400), .B(new_n369), .C1(new_n404), .C2(new_n380), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n293), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n366), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(G234), .A2(G237), .ZN(new_n412));
  INV_X1    g226(.A(G953), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(G952), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT21), .B(G898), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(G902), .A3(G953), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n396), .A3(G104), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT3), .B1(new_n341), .B2(G107), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n341), .A2(G107), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(G101), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(G101), .ZN(new_n432));
  INV_X1    g246(.A(G101), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n194), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n437));
  NOR2_X1   g251(.A1(new_n373), .A2(G119), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n189), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n193), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n439), .A2(new_n441), .B1(new_n192), .B2(new_n193), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n396), .A2(G104), .ZN(new_n443));
  OAI21_X1  g257(.A(G101), .B1(new_n428), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n434), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n436), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(G110), .A2(G122), .ZN(new_n448));
  NAND2_X1  g262(.A1(G110), .A2(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n436), .A2(new_n454), .A3(new_n446), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT6), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n230), .A2(G125), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n215), .A2(new_n218), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n302), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n413), .A2(G224), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT83), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n462), .B(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n447), .A2(new_n467), .A3(new_n455), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n458), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n439), .A2(new_n441), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n434), .A2(new_n444), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n192), .A2(new_n193), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n454), .A2(KEYINPUT8), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n451), .A2(new_n477), .A3(new_n453), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n193), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n439), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n473), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n471), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n474), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n445), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n442), .A2(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT85), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n462), .A2(KEYINPUT7), .A3(new_n465), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n459), .B(new_n461), .C1(new_n493), .C2(new_n464), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n487), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n457), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n293), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n424), .B1(new_n470), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(new_n469), .A3(new_n293), .A4(new_n423), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G214), .B1(G237), .B2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n218), .A2(KEYINPUT79), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n225), .A2(new_n505), .A3(new_n217), .A4(G128), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n215), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n445), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT10), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n473), .A2(new_n509), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n219), .B2(new_n220), .ZN(new_n512));
  INV_X1    g326(.A(new_n233), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n230), .A2(new_n435), .A3(new_n431), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n510), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G110), .B(G140), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n413), .A2(G227), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n516), .B(new_n517), .Z(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT80), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n233), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n515), .A2(KEYINPUT80), .A3(new_n518), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n238), .A2(new_n473), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n508), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT12), .B1(new_n527), .B2(new_n233), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n529), .B(new_n513), .C1(new_n508), .C2(new_n526), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n515), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n525), .A2(G469), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n515), .B(new_n518), .C1(new_n528), .C2(new_n530), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n518), .B1(new_n523), .B2(new_n515), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n535), .B(new_n293), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n535), .A2(new_n293), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n422), .A2(new_n503), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n368), .B1(G234), .B2(new_n293), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n548));
  INV_X1    g362(.A(G119), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G128), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT23), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT73), .B1(new_n214), .B2(G119), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(G128), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT23), .B(new_n550), .C1(new_n554), .C2(KEYINPUT73), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT74), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n555), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(KEYINPUT75), .A3(G110), .A4(new_n556), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n337), .A2(new_n338), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT72), .ZN(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n559), .A2(new_n563), .A3(new_n564), .A4(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n560), .A2(G110), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n306), .B(new_n338), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n413), .A2(G221), .A3(G234), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n572), .A3(new_n576), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n293), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n547), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n578), .A2(new_n293), .A3(new_n579), .A4(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n578), .A2(new_n579), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n546), .A2(G902), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n583), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n301), .A2(new_n545), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n402), .B2(new_n405), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(G478), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n407), .A2(KEYINPUT91), .A3(new_n408), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n402), .A2(KEYINPUT33), .A3(new_n405), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT33), .B1(new_n402), .B2(new_n405), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n408), .A2(G902), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n595), .A2(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n348), .B1(new_n358), .B2(new_n343), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT20), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n603), .A2(new_n359), .B1(G475), .B2(new_n345), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n592), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n598), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n402), .A2(KEYINPUT33), .A3(new_n405), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n600), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT91), .B1(new_n407), .B2(new_n408), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n594), .A2(new_n593), .A3(G478), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n366), .A3(KEYINPUT92), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n502), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n498), .B2(new_n500), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n421), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT93), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n420), .B(new_n614), .C1(new_n498), .C2(new_n500), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT93), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n605), .A4(new_n612), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n271), .A2(new_n293), .A3(new_n273), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n589), .A2(new_n542), .A3(new_n543), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n275), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT90), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(new_n624), .A3(new_n627), .A4(new_n275), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n621), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  XOR2_X1   g445(.A(new_n420), .B(KEYINPUT94), .Z(new_n632));
  AND2_X1   g446(.A1(new_n615), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n633), .A2(new_n410), .A3(new_n604), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n626), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n623), .A2(new_n275), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n583), .A2(new_n586), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n573), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n588), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n640), .A2(KEYINPUT95), .A3(new_n643), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n639), .A2(new_n545), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  NOR2_X1   g465(.A1(new_n503), .A2(new_n544), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n604), .A2(new_n410), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n419), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n414), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n301), .A2(new_n652), .A3(new_n648), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  INV_X1    g474(.A(new_n544), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT96), .B(KEYINPUT39), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n656), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n501), .B(KEYINPUT38), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n366), .A2(new_n410), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n644), .A2(new_n667), .A3(new_n614), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n266), .B1(new_n248), .B2(new_n250), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n291), .A2(new_n250), .A3(new_n266), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n293), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n277), .A2(new_n278), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n669), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n208), .ZN(G45));
  NOR3_X1   g492(.A1(new_n601), .A2(new_n604), .A3(new_n657), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n301), .A2(new_n652), .A3(new_n648), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n684), .A2(new_n511), .B1(new_n508), .B2(new_n509), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n513), .B1(new_n685), .B2(new_n514), .ZN(new_n686));
  INV_X1    g500(.A(new_n515), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n532), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(G902), .B1(new_n688), .B2(new_n536), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n535), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n543), .A3(new_n539), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n621), .A2(new_n589), .A3(new_n301), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT97), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G15));
  NAND4_X1  g511(.A1(new_n301), .A2(new_n634), .A3(new_n589), .A4(new_n693), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT98), .B(G116), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G18));
  NOR3_X1   g514(.A1(new_n422), .A2(new_n692), .A3(new_n503), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n297), .A2(new_n300), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n277), .A2(new_n278), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n648), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT99), .B(G119), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G21));
  AND4_X1   g520(.A1(new_n410), .A2(new_n615), .A3(new_n366), .A4(new_n632), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n284), .A2(new_n291), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n257), .B(new_n269), .C1(new_n708), .C2(new_n255), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n622), .A2(G472), .B1(new_n274), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n710), .A3(new_n589), .A4(new_n693), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  AND2_X1   g526(.A1(new_n710), .A2(new_n644), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n692), .A2(new_n503), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n679), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  INV_X1    g530(.A(new_n543), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n540), .B1(new_n689), .B2(new_n535), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n531), .A2(new_n719), .A3(new_n532), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n719), .B1(new_n531), .B2(new_n532), .ZN(new_n721));
  OAI211_X1 g535(.A(G469), .B(new_n525), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n717), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n679), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n301), .A2(new_n589), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n589), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n277), .A2(new_n278), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n288), .A2(new_n286), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n282), .B1(new_n279), .B2(new_n266), .ZN(new_n732));
  AOI211_X1 g546(.A(KEYINPUT70), .B(new_n255), .C1(new_n248), .C2(new_n250), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n294), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n298), .B1(new_n735), .B2(new_n299), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n296), .A2(KEYINPUT71), .A3(G472), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n729), .B1(new_n730), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n725), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  AND3_X1   g556(.A1(new_n658), .A2(new_n723), .A3(new_n724), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n301), .A2(new_n589), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n195), .ZN(G36));
  OAI211_X1 g559(.A(KEYINPUT45), .B(new_n525), .C1(new_n720), .C2(new_n721), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n525), .A2(new_n533), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n746), .B(G469), .C1(new_n747), .C2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n541), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT101), .B1(new_n749), .B2(new_n539), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(KEYINPUT101), .A3(new_n539), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n748), .A2(new_n541), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n751), .B(new_n752), .C1(KEYINPUT46), .C2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n717), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n663), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n601), .A2(new_n366), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT43), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n638), .A3(new_n644), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n762), .B2(new_n761), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n756), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n717), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n679), .A2(new_n729), .A3(new_n724), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n301), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  NAND2_X1  g588(.A1(new_n691), .A2(new_n539), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT102), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT49), .Z(new_n777));
  NAND3_X1  g591(.A1(new_n759), .A2(new_n502), .A3(new_n543), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n666), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n589), .A3(new_n675), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n760), .A2(new_n415), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n710), .A2(new_n589), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n666), .A2(new_n502), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n693), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT50), .Z(new_n785));
  NOR3_X1   g599(.A1(new_n692), .A2(new_n414), .A3(new_n758), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n713), .A2(new_n760), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n675), .A2(new_n589), .A3(new_n786), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n611), .A2(new_n366), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n776), .A2(new_n717), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n768), .B2(new_n769), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n781), .A2(new_n782), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n724), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n796), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n804), .B1(new_n803), .B2(new_n805), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT104), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n545), .A2(new_n648), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n739), .A2(new_n545), .B1(new_n809), .B2(new_n639), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n704), .A2(new_n711), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n739), .B(new_n693), .C1(new_n621), .C2(new_n634), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n653), .B1(new_n604), .B2(new_n601), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n633), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n626), .A2(new_n628), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n744), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n725), .A2(new_n644), .A3(new_n710), .ZN(new_n818));
  INV_X1    g632(.A(new_n648), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n730), .B2(new_n738), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT103), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n411), .A2(new_n656), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n758), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n724), .A2(KEYINPUT103), .A3(new_n411), .A4(new_n656), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(new_n661), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n818), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT42), .B1(new_n739), .B2(new_n725), .ZN(new_n827));
  AND4_X1   g641(.A1(KEYINPUT42), .A2(new_n301), .A3(new_n589), .A4(new_n725), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n817), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n808), .B1(new_n816), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n694), .A2(new_n698), .A3(new_n815), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n590), .A2(new_n704), .A3(new_n649), .A4(new_n711), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n744), .B1(new_n728), .B2(new_n740), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(KEYINPUT104), .A3(new_n834), .A4(new_n826), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n503), .A2(new_n667), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n644), .A2(new_n657), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n674), .A2(new_n836), .A3(new_n723), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n659), .A2(new_n680), .A3(new_n715), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n830), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT54), .ZN(new_n845));
  XOR2_X1   g659(.A(KEYINPUT106), .B(KEYINPUT54), .Z(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n816), .A2(new_n829), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n841), .A2(new_n848), .A3(KEYINPUT53), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n842), .A2(KEYINPUT105), .A3(new_n843), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT105), .B1(new_n842), .B2(new_n843), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n847), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n801), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n856));
  OAI211_X1 g670(.A(KEYINPUT51), .B(new_n795), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n800), .A2(new_n714), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(G952), .A3(new_n413), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n789), .A2(new_n605), .A3(new_n612), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT111), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT111), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT48), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n739), .A2(new_n760), .A3(new_n786), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n863), .A2(KEYINPUT48), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n857), .A2(new_n861), .A3(new_n862), .A4(new_n867), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n806), .A2(new_n807), .A3(new_n853), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n780), .B1(new_n869), .B2(new_n870), .ZN(G75));
  OAI21_X1  g685(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(G210), .A3(G902), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n458), .A2(new_n468), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n466), .ZN(new_n879));
  INV_X1    g693(.A(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n877), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n413), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  NAND2_X1  g699(.A1(new_n872), .A2(new_n846), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(KEYINPUT114), .A3(new_n852), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n872), .A2(new_n888), .A3(new_n846), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n540), .B(KEYINPUT57), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n538), .B2(new_n537), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n872), .A2(G902), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(new_n748), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n884), .B1(new_n892), .B2(new_n894), .ZN(G54));
  NAND2_X1  g709(.A1(KEYINPUT58), .A2(G475), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n872), .A2(G902), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n364), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR3_X1    g714(.A1(new_n898), .A2(KEYINPUT116), .A3(new_n899), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT116), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n884), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(G60));
  XOR2_X1   g717(.A(new_n599), .B(KEYINPUT117), .Z(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n887), .A2(new_n889), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n884), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(KEYINPUT119), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT119), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n904), .B1(new_n853), .B2(new_n907), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n872), .A2(new_n642), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n910), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n587), .B1(new_n872), .B2(new_n917), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n921), .B(new_n922), .Z(G66));
  INV_X1    g737(.A(G224), .ZN(new_n924));
  OAI21_X1  g738(.A(G953), .B1(new_n417), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n833), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n878), .B1(G898), .B2(new_n413), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT121), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  NAND2_X1  g743(.A1(new_n654), .A2(G953), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT124), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n773), .A2(new_n765), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n659), .A2(new_n680), .A3(new_n715), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n739), .A2(new_n836), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n757), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n933), .A2(new_n834), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n932), .B1(new_n938), .B2(new_n413), .ZN(new_n939));
  MUX2_X1   g753(.A(new_n247), .B(new_n290), .S(KEYINPUT30), .Z(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(new_n351), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n677), .B1(new_n944), .B2(KEYINPUT62), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n935), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n944), .A3(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n944), .B2(KEYINPUT62), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n664), .A2(new_n758), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n739), .A2(new_n813), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n933), .A2(new_n948), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n952), .B2(new_n413), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n943), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT123), .B1(new_n939), .B2(new_n942), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n413), .B1(G227), .B2(G900), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n954), .B(new_n958), .ZN(G72));
  XNOR2_X1  g773(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n299), .A2(new_n293), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n938), .B2(new_n816), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n279), .A2(new_n255), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n962), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n734), .B2(new_n256), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT127), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n844), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n952), .B2(new_n816), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n884), .B1(new_n972), .B2(new_n670), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n967), .A2(new_n971), .A3(new_n973), .ZN(G57));
endmodule


