//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G141gat), .B(G148gat), .Z(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT2), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n204), .A2(new_n207), .B1(new_n208), .B2(KEYINPUT74), .ZN(new_n209));
  INV_X1    g008(.A(new_n208), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n210), .A2(new_n204), .A3(new_n211), .A4(new_n207), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT75), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n218));
  INV_X1    g017(.A(G113gat), .ZN(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT1), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n219), .B2(new_n220), .ZN(new_n222));
  INV_X1    g021(.A(G127gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G134gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(G134gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n222), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT68), .B(G120gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G113gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n223), .A2(G134gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n231), .A2(new_n221), .A3(new_n224), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n218), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n217), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n214), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n238), .B(KEYINPUT76), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(new_n234), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n203), .B1(new_n237), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT39), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n215), .A2(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n239), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n202), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT0), .ZN(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G85gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  OAI211_X1 g055(.A(new_n247), .B(new_n203), .C1(new_n237), .C2(new_n245), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT40), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT81), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n252), .A2(KEYINPUT40), .A3(new_n256), .A4(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT83), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n257), .A2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT40), .A4(new_n252), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n249), .B2(new_n203), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT77), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n269), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n203), .B1(new_n217), .B2(new_n236), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT4), .B1(new_n235), .B2(new_n238), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n243), .B2(KEYINPUT4), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n243), .A2(new_n244), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n240), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n277), .A2(new_n272), .A3(new_n267), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT82), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n270), .A2(new_n271), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n274), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n272), .A3(new_n267), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n256), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G8gat), .B(G36gat), .Z(new_n288));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G211gat), .B(G218gat), .Z(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n292), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n309), .A2(KEYINPUT27), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n304), .B1(new_n310), .B2(KEYINPUT64), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n306), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n316), .A2(KEYINPUT26), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n317), .A2(KEYINPUT26), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n317), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT24), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n316), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n304), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT24), .A3(new_n319), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n330), .B(KEYINPUT25), .Z(new_n331));
  NAND2_X1  g130(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G226gat), .ZN(new_n335));
  INV_X1    g134(.A(G233gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(G226gat), .A3(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n339), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n300), .B(new_n337), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n299), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n290), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n342), .A2(new_n290), .A3(new_n344), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(KEYINPUT30), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n290), .A3(new_n344), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n348), .A2(KEYINPUT73), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT73), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT40), .B1(new_n263), .B2(new_n252), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(KEYINPUT81), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n266), .A2(new_n287), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n299), .B1(new_n218), .B2(KEYINPUT29), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(new_n299), .B2(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n215), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n298), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n362), .A2(new_n291), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n333), .B1(new_n362), .B2(new_n291), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n242), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n357), .A2(new_n356), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G22gat), .ZN(new_n369));
  XOR2_X1   g168(.A(G78gat), .B(G106gat), .Z(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT31), .B(G50gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT79), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n368), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n282), .A2(new_n256), .A3(new_n284), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n287), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT84), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n286), .B(new_n385), .C1(new_n275), .C2(new_n278), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n287), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n342), .A2(new_n344), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT37), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n290), .A2(new_n391), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n390), .A2(new_n391), .B1(new_n345), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n346), .B1(new_n393), .B2(KEYINPUT38), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n343), .B2(new_n300), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n300), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT85), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n345), .B2(new_n392), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n355), .B(new_n379), .C1(new_n389), .C2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n379), .B(KEYINPUT80), .ZN(new_n403));
  INV_X1    g202(.A(new_n352), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n286), .B1(new_n275), .B2(new_n278), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n380), .A3(new_n381), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n386), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT34), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n323), .A2(new_n331), .A3(new_n234), .ZN(new_n412));
  INV_X1    g211(.A(new_n322), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n305), .B2(new_n312), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n330), .B(KEYINPUT25), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n235), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n416), .A3(new_n409), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT32), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT69), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n421));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n417), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n412), .A2(new_n416), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n409), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n417), .B(KEYINPUT32), .C1(new_n425), .C2(new_n424), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n427), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n411), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n429), .ZN(new_n437));
  INV_X1    g236(.A(new_n411), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n432), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(KEYINPUT36), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT36), .B1(new_n435), .B2(new_n439), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n403), .A2(new_n408), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444));
  INV_X1    g243(.A(new_n379), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n433), .A2(new_n411), .A3(new_n434), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n438), .B1(new_n437), .B2(new_n432), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n389), .A2(new_n444), .A3(new_n448), .A4(new_n404), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n446), .A2(new_n447), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n379), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT35), .B1(new_n408), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n402), .A2(new_n443), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(G1gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT16), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n455), .A2(G1gat), .ZN(new_n459));
  OAI21_X1  g258(.A(G8gat), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n457), .ZN(new_n461));
  INV_X1    g260(.A(G8gat), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n462), .C1(G1gat), .C2(new_n455), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT15), .ZN(new_n465));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(KEYINPUT87), .ZN(new_n467));
  INV_X1    g266(.A(G43gat), .ZN(new_n468));
  INV_X1    g267(.A(G50gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g270(.A1(G43gat), .A2(G50gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n475));
  INV_X1    g274(.A(G29gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n478));
  AOI21_X1  g277(.A(G36gat), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G36gat), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n475), .A2(new_n480), .A3(G29gat), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n479), .A2(new_n481), .B1(KEYINPUT15), .B2(new_n466), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n467), .B(new_n473), .C1(new_n479), .C2(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n454), .B1(new_n464), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n460), .A2(new_n463), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(KEYINPUT88), .A3(new_n483), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(KEYINPUT17), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n483), .A2(new_n492), .A3(new_n484), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n464), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT18), .B1(new_n495), .B2(KEYINPUT89), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n489), .A2(new_n498), .A3(new_n490), .A4(new_n494), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n464), .A2(new_n485), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n489), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n490), .B(KEYINPUT13), .Z(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n489), .A2(KEYINPUT18), .A3(new_n490), .A4(new_n494), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT86), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT11), .B(G169gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT12), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n504), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n500), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n497), .B1(new_n496), .B2(new_n499), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n504), .A2(new_n505), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n499), .B2(new_n496), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n513), .A2(new_n514), .B1(new_n516), .B2(new_n511), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n453), .A2(new_n518), .ZN(new_n519));
  AND4_X1   g318(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n520));
  AOI22_X1  g319(.A1(KEYINPUT98), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT8), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n525));
  OR2_X1    g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G99gat), .B(G106gat), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(new_n522), .C1(new_n527), .C2(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(KEYINPUT101), .ZN(new_n535));
  NAND2_X1  g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  OR2_X1    g335(.A1(G71gat), .A2(G78gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(KEYINPUT91), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G57gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G64gat), .ZN(new_n545));
  INV_X1    g344(.A(G64gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G57gat), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n536), .B(new_n537), .C1(new_n543), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n536), .A2(KEYINPUT91), .A3(new_n538), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT91), .B1(new_n536), .B2(new_n538), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(KEYINPUT93), .A3(new_n542), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT92), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n546), .A2(G57gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n556), .A2(new_n557), .B1(new_n537), .B2(new_n536), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n534), .A2(new_n535), .A3(new_n549), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n549), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n533), .B(new_n531), .C1(new_n561), .C2(KEYINPUT101), .ZN(new_n562));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n565), .A2(KEYINPUT103), .ZN(new_n566));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n565), .B2(KEYINPUT103), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n534), .A2(new_n561), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n560), .A2(new_n562), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT102), .B1(new_n575), .B2(new_n564), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT10), .B1(new_n560), .B2(new_n562), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n577), .B(new_n563), .C1(new_n578), .C2(new_n573), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT104), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n571), .A2(new_n576), .A3(KEYINPUT104), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n565), .B1(new_n575), .B2(new_n564), .ZN(new_n585));
  INV_X1    g384(.A(new_n569), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n561), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n464), .B1(new_n561), .B2(new_n589), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT95), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT94), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n594), .B(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n534), .A2(new_n485), .ZN(new_n603));
  NAND3_X1  g402(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n491), .A2(new_n493), .A3(new_n534), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  INV_X1    g409(.A(new_n607), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n605), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT97), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT100), .ZN(new_n619));
  INV_X1    g418(.A(new_n609), .ZN(new_n620));
  INV_X1    g419(.A(new_n612), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n609), .A2(new_n612), .A3(new_n623), .A4(new_n617), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n588), .A2(new_n602), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n519), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n407), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g429(.A(KEYINPUT16), .B(G8gat), .Z(new_n631));
  NAND4_X1  g430(.A1(new_n519), .A2(new_n352), .A3(new_n626), .A4(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n519), .A2(new_n352), .A3(new_n626), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n462), .ZN(new_n634));
  MUX2_X1   g433(.A(new_n632), .B(new_n634), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n636), .A3(new_n450), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n442), .A2(new_n440), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(new_n636), .ZN(G1326gat));
  NAND2_X1  g440(.A1(new_n627), .A2(new_n403), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT43), .B(G22gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  INV_X1    g443(.A(new_n625), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n453), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n588), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n602), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n518), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n646), .A2(new_n476), .A3(new_n628), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT45), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n402), .A2(new_n443), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n449), .A2(new_n452), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(KEYINPUT44), .A3(new_n625), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n453), .B2(new_n645), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n658), .A2(new_n628), .A3(new_n649), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n651), .B1(new_n659), .B2(new_n476), .ZN(G1328gat));
  NAND4_X1  g459(.A1(new_n655), .A2(new_n657), .A3(new_n352), .A4(new_n649), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n480), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n646), .A2(new_n480), .A3(new_n352), .A4(new_n649), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(G1329gat));
  NOR2_X1   g467(.A1(new_n638), .A2(new_n468), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n655), .A2(new_n657), .A3(new_n649), .A4(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n646), .A2(new_n450), .A3(new_n649), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(G43gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g472(.A1(new_n655), .A2(new_n657), .A3(new_n445), .A4(new_n649), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G50gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n403), .A2(new_n469), .A3(new_n625), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n648), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n519), .A2(KEYINPUT107), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n655), .A2(new_n657), .A3(new_n403), .A4(new_n649), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT48), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n681), .A3(G50gat), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n519), .A2(new_n677), .B1(KEYINPUT107), .B2(KEYINPUT48), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n679), .A2(KEYINPUT48), .B1(new_n682), .B2(new_n683), .ZN(G1331gat));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n517), .A2(new_n602), .A3(new_n625), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n654), .A2(new_n685), .A3(new_n588), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n588), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n453), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n628), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n352), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT49), .B(G64gat), .Z(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(G1333gat));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n689), .A3(new_n639), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G71gat), .ZN(new_n698));
  INV_X1    g497(.A(G71gat), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n687), .A2(new_n689), .A3(new_n699), .A4(new_n450), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n698), .B2(new_n700), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(G1334gat));
  NAND2_X1  g503(.A1(new_n690), .A2(new_n403), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G78gat), .ZN(G1335gat));
  INV_X1    g505(.A(new_n602), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n517), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n654), .A2(new_n625), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n646), .A2(KEYINPUT51), .A3(new_n708), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n647), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(G85gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n628), .ZN(new_n715));
  INV_X1    g514(.A(new_n708), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n647), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n658), .A2(new_n628), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n718), .B2(new_n714), .ZN(G1336gat));
  NAND2_X1  g518(.A1(new_n711), .A2(new_n712), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n404), .A2(G92gat), .A3(new_n647), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n655), .A2(new_n657), .A3(new_n352), .A4(new_n717), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G92gat), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n721), .B(KEYINPUT110), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n720), .A2(new_n727), .B1(new_n723), .B2(G92gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(new_n725), .ZN(G1337gat));
  INV_X1    g528(.A(G99gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n730), .A3(new_n450), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n658), .A2(new_n639), .A3(new_n717), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n730), .ZN(G1338gat));
  NOR2_X1   g532(.A1(new_n379), .A2(G106gat), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT51), .B1(new_n646), .B2(new_n708), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n453), .A2(new_n710), .A3(new_n645), .A4(new_n716), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n588), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT53), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n655), .A2(new_n657), .A3(new_n445), .A4(new_n717), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G106gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n655), .A2(new_n657), .A3(new_n403), .A4(new_n717), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n713), .A2(new_n734), .B1(G106gat), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n738), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT54), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n575), .B2(new_n564), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n576), .A2(new_n746), .A3(new_n579), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n745), .B(new_n563), .C1(new_n578), .C2(new_n573), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n586), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(KEYINPUT55), .B1(new_n582), .B2(new_n583), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n747), .A2(new_n749), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT111), .B(KEYINPUT55), .C1(new_n747), .C2(new_n749), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n751), .B(new_n517), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT18), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n759), .A3(new_n499), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT90), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n500), .A3(new_n512), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n502), .A2(new_n503), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n490), .B1(new_n489), .B2(new_n494), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n510), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n767), .B(new_n510), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n588), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n625), .B1(new_n757), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n756), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n747), .A2(KEYINPUT55), .A3(new_n749), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n584), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n625), .A2(new_n762), .A3(new_n769), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n602), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n686), .A2(new_n647), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n403), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n352), .A2(new_n407), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n450), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G113gat), .B1(new_n782), .B2(new_n518), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n407), .B1(new_n778), .B2(new_n779), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n448), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n404), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n517), .A2(new_n219), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT114), .Z(new_n789));
  OAI21_X1  g588(.A(new_n783), .B1(new_n787), .B2(new_n789), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n782), .B2(new_n647), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n647), .A2(new_n230), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n787), .B2(new_n792), .ZN(G1341gat));
  OAI21_X1  g592(.A(G127gat), .B1(new_n782), .B2(new_n602), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n707), .A2(new_n223), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n787), .B2(new_n795), .ZN(G1342gat));
  NOR2_X1   g595(.A1(new_n645), .A2(new_n227), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n404), .A3(new_n797), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n799));
  OAI21_X1  g598(.A(G134gat), .B1(new_n782), .B2(new_n645), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(G1343gat));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n639), .A2(new_n379), .A3(new_n352), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n518), .A2(G141gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n638), .A2(new_n781), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n753), .A2(new_n754), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n517), .A2(new_n584), .A3(new_n808), .A4(new_n774), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n625), .B1(new_n771), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n602), .B1(new_n810), .B2(new_n777), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n779), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n403), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n807), .B1(new_n813), .B2(KEYINPUT57), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n445), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n778), .B2(new_n779), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n517), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n820));
  OAI21_X1  g619(.A(G141gat), .B1(new_n819), .B2(KEYINPUT117), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n803), .B(new_n806), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n819), .A2(G141gat), .B1(new_n824), .B2(new_n806), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n784), .A2(new_n804), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT115), .A3(new_n805), .ZN(new_n828));
  AOI211_X1 g627(.A(new_n823), .B(new_n803), .C1(new_n825), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n819), .A2(G141gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n806), .A2(new_n824), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT116), .B1(new_n832), .B2(KEYINPUT58), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n822), .B1(new_n829), .B2(new_n833), .ZN(G1344gat));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G148gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n815), .B1(new_n812), .B2(new_n403), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n817), .A3(new_n807), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n839), .B2(new_n588), .ZN(new_n840));
  INV_X1    g639(.A(new_n440), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n781), .B(KEYINPUT118), .C1(new_n841), .C2(new_n441), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n588), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT118), .B1(new_n638), .B2(new_n781), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n812), .B2(new_n403), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n445), .A2(KEYINPUT57), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n778), .B2(new_n779), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT119), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n845), .B(new_n851), .C1(new_n846), .C2(new_n848), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(G148gat), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n840), .B1(new_n853), .B2(KEYINPUT59), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n826), .A2(G148gat), .A3(new_n647), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n835), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n855), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n852), .A2(G148gat), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n836), .B1(new_n858), .B2(new_n850), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT120), .B(new_n857), .C1(new_n859), .C2(new_n840), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(G1345gat));
  INV_X1    g660(.A(new_n839), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n205), .A3(new_n602), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n826), .A2(new_n602), .ZN(new_n864));
  AOI21_X1  g663(.A(G155gat), .B1(new_n864), .B2(KEYINPUT121), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n864), .A2(KEYINPUT121), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(G1346gat));
  OAI21_X1  g666(.A(G162gat), .B1(new_n862), .B2(new_n645), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n827), .A2(new_n206), .A3(new_n625), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1347gat));
  AOI21_X1  g669(.A(new_n628), .B1(new_n778), .B2(new_n779), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n451), .A2(new_n404), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n314), .A3(new_n517), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT122), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n352), .A2(new_n407), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n446), .A3(new_n447), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n780), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n518), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT123), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n881), .ZN(G1348gat));
  NOR3_X1   g681(.A1(new_n873), .A2(G176gat), .A3(new_n647), .ZN(new_n883));
  INV_X1    g682(.A(new_n879), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n588), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(G176gat), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT124), .Z(G1349gat));
  NAND3_X1  g686(.A1(new_n874), .A2(new_n303), .A3(new_n707), .ZN(new_n888));
  OAI21_X1  g687(.A(G183gat), .B1(new_n879), .B2(new_n602), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n304), .A3(new_n625), .ZN(new_n892));
  OAI21_X1  g691(.A(G190gat), .B1(new_n879), .B2(new_n645), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n846), .A2(new_n848), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n639), .A2(new_n877), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n517), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G197gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n871), .A2(new_n445), .A3(new_n352), .A4(new_n638), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n904), .A2(G197gat), .A3(new_n518), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1352gat));
  NOR3_X1   g707(.A1(new_n904), .A2(G204gat), .A3(new_n647), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n900), .A2(new_n588), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G204gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n910), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(G1353gat));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n707), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT63), .B1(new_n917), .B2(new_n295), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n904), .A2(G211gat), .A3(new_n602), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT126), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n921), .A3(G211gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n920), .A3(new_n922), .ZN(G1354gat));
  NAND2_X1  g722(.A1(new_n900), .A2(new_n625), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G218gat), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n904), .A2(G218gat), .A3(new_n645), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1355gat));
endmodule


