

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776;

  OR2_X1 U374 ( .A1(n511), .A2(G902), .ZN(n386) );
  NOR2_X1 U375 ( .A1(n374), .A2(n692), .ZN(n637) );
  INV_X2 U376 ( .A(G953), .ZN(n758) );
  BUF_X1 U377 ( .A(G122), .Z(n356) );
  AND2_X1 U378 ( .A1(n446), .A2(n358), .ZN(n353) );
  XNOR2_X2 U379 ( .A(n578), .B(KEYINPUT73), .ZN(n588) );
  XNOR2_X2 U380 ( .A(n604), .B(n603), .ZN(n396) );
  AND2_X2 U381 ( .A1(n600), .A2(n601), .ZN(n604) );
  NOR2_X2 U382 ( .A1(n628), .A2(n717), .ZN(n629) );
  INV_X2 U383 ( .A(G143), .ZN(n482) );
  XNOR2_X2 U384 ( .A(n432), .B(n431), .ZN(n771) );
  XNOR2_X1 U385 ( .A(n386), .B(G472), .ZN(n555) );
  INV_X1 U386 ( .A(KEYINPUT32), .ZN(n431) );
  NOR2_X1 U387 ( .A1(n757), .A2(n404), .ZN(n725) );
  BUF_X1 U388 ( .A(n680), .Z(n354) );
  NAND2_X1 U389 ( .A1(n618), .A2(n434), .ZN(n433) );
  XNOR2_X1 U390 ( .A(n446), .B(KEYINPUT101), .ZN(n686) );
  XNOR2_X1 U391 ( .A(n555), .B(KEYINPUT102), .ZN(n619) );
  XNOR2_X1 U392 ( .A(n537), .B(n490), .ZN(n511) );
  XNOR2_X1 U393 ( .A(n549), .B(n463), .ZN(n517) );
  XNOR2_X1 U394 ( .A(n444), .B(G146), .ZN(n549) );
  XOR2_X1 U395 ( .A(KEYINPUT16), .B(KEYINPUT70), .Z(n544) );
  XOR2_X1 U396 ( .A(G137), .B(KEYINPUT5), .Z(n485) );
  INV_X2 U397 ( .A(KEYINPUT66), .ZN(n453) );
  XNOR2_X1 U398 ( .A(KEYINPUT3), .B(G119), .ZN(n487) );
  XNOR2_X1 U399 ( .A(n639), .B(n640), .ZN(n680) );
  BUF_X1 U400 ( .A(n543), .Z(n355) );
  XNOR2_X1 U401 ( .A(n488), .B(n487), .ZN(n543) );
  XNOR2_X1 U402 ( .A(n542), .B(n544), .ZN(n476) );
  NOR2_X2 U403 ( .A1(n559), .A2(n558), .ZN(n595) );
  NAND2_X2 U404 ( .A1(n390), .A2(n387), .ZN(n757) );
  BUF_X1 U405 ( .A(n748), .Z(n357) );
  XNOR2_X1 U406 ( .A(n476), .B(n543), .ZN(n748) );
  XNOR2_X2 U407 ( .A(n439), .B(n364), .ZN(n755) );
  NOR2_X1 U408 ( .A1(n575), .A2(n360), .ZN(n447) );
  XNOR2_X1 U409 ( .A(n457), .B(n456), .ZN(n706) );
  INV_X1 U410 ( .A(KEYINPUT99), .ZN(n456) );
  NOR2_X1 U411 ( .A1(n757), .A2(n418), .ZN(n401) );
  NOR2_X1 U412 ( .A1(n705), .A2(n704), .ZN(n594) );
  INV_X1 U413 ( .A(KEYINPUT77), .ZN(n378) );
  INV_X1 U414 ( .A(G125), .ZN(n444) );
  XOR2_X1 U415 ( .A(G902), .B(KEYINPUT15), .Z(n653) );
  XOR2_X1 U416 ( .A(KEYINPUT11), .B(G131), .Z(n500) );
  XNOR2_X1 U417 ( .A(G113), .B(G143), .ZN(n499) );
  INV_X1 U418 ( .A(KEYINPUT10), .ZN(n463) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n503) );
  NAND2_X1 U420 ( .A1(G234), .A2(G237), .ZN(n515) );
  XOR2_X1 U421 ( .A(KEYINPUT81), .B(KEYINPUT45), .Z(n651) );
  XNOR2_X1 U422 ( .A(n585), .B(n454), .ZN(n702) );
  XNOR2_X1 U423 ( .A(n455), .B(KEYINPUT38), .ZN(n454) );
  INV_X1 U424 ( .A(KEYINPUT72), .ZN(n455) );
  INV_X1 U425 ( .A(KEYINPUT85), .ZN(n561) );
  AND2_X1 U426 ( .A1(n677), .A2(n623), .ZN(n532) );
  AND2_X1 U427 ( .A1(n394), .A2(n391), .ZN(n390) );
  INV_X1 U428 ( .A(KEYINPUT83), .ZN(n388) );
  NAND2_X1 U429 ( .A1(n521), .A2(G217), .ZN(n460) );
  XOR2_X1 U430 ( .A(KEYINPUT96), .B(G107), .Z(n496) );
  INV_X1 U431 ( .A(n725), .ZN(n440) );
  INV_X1 U432 ( .A(G104), .ZN(n451) );
  XOR2_X1 U433 ( .A(G137), .B(G140), .Z(n533) );
  XNOR2_X1 U434 ( .A(n452), .B(n579), .ZN(n586) );
  NAND2_X1 U435 ( .A1(n619), .A2(n701), .ZN(n452) );
  INV_X1 U436 ( .A(KEYINPUT125), .ZN(n469) );
  AND2_X1 U437 ( .A1(n731), .A2(n758), .ZN(n438) );
  NOR2_X1 U438 ( .A1(n706), .A2(n672), .ZN(n573) );
  OR2_X1 U439 ( .A1(n706), .A2(KEYINPUT71), .ZN(n565) );
  INV_X1 U440 ( .A(KEYINPUT44), .ZN(n415) );
  OR2_X1 U441 ( .A1(G237), .A2(G902), .ZN(n550) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n501) );
  NOR2_X1 U443 ( .A1(n393), .A2(n392), .ZN(n391) );
  INV_X1 U444 ( .A(n684), .ZN(n392) );
  NOR2_X1 U445 ( .A1(n765), .A2(KEYINPUT83), .ZN(n393) );
  XNOR2_X1 U446 ( .A(G119), .B(G128), .ZN(n518) );
  XNOR2_X1 U447 ( .A(n517), .B(n462), .ZN(n756) );
  INV_X1 U448 ( .A(n533), .ZN(n462) );
  NAND2_X1 U449 ( .A1(n373), .A2(n406), .ZN(n405) );
  XNOR2_X1 U450 ( .A(n654), .B(n421), .ZN(n384) );
  INV_X1 U451 ( .A(KEYINPUT80), .ZN(n421) );
  XNOR2_X1 U452 ( .A(n546), .B(n385), .ZN(n547) );
  XNOR2_X1 U453 ( .A(KEYINPUT18), .B(KEYINPUT74), .ZN(n385) );
  INV_X1 U454 ( .A(n549), .ZN(n449) );
  AND2_X1 U455 ( .A1(n619), .A2(n353), .ZN(n556) );
  NAND2_X1 U456 ( .A1(n702), .A2(n701), .ZN(n705) );
  XNOR2_X1 U457 ( .A(n529), .B(n359), .ZN(n473) );
  XNOR2_X1 U458 ( .A(n506), .B(n443), .ZN(n656) );
  XNOR2_X1 U459 ( .A(n507), .B(n505), .ZN(n443) );
  AND2_X1 U460 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U461 ( .A(KEYINPUT0), .ZN(n471) );
  XNOR2_X1 U462 ( .A(n690), .B(n512), .ZN(n623) );
  AND2_X1 U463 ( .A1(n586), .A2(n702), .ZN(n587) );
  INV_X1 U464 ( .A(n686), .ZN(n434) );
  NAND2_X1 U465 ( .A1(n595), .A2(n612), .ZN(n672) );
  NAND2_X1 U466 ( .A1(n620), .A2(KEYINPUT103), .ZN(n429) );
  NOR2_X1 U467 ( .A1(n620), .A2(KEYINPUT103), .ZN(n427) );
  BUF_X1 U468 ( .A(n473), .Z(n446) );
  XNOR2_X1 U469 ( .A(n459), .B(n458), .ZN(n738) );
  XNOR2_X1 U470 ( .A(n497), .B(n362), .ZN(n458) );
  XNOR2_X1 U471 ( .A(n460), .B(n494), .ZN(n459) );
  XNOR2_X1 U472 ( .A(n533), .B(n450), .ZN(n535) );
  XNOR2_X1 U473 ( .A(n534), .B(n451), .ZN(n450) );
  XNOR2_X1 U474 ( .A(n597), .B(n596), .ZN(n775) );
  XNOR2_X1 U475 ( .A(n467), .B(n466), .ZN(n465) );
  INV_X1 U476 ( .A(KEYINPUT36), .ZN(n466) );
  INV_X1 U477 ( .A(KEYINPUT35), .ZN(n634) );
  XNOR2_X1 U478 ( .A(KEYINPUT107), .B(n582), .ZN(n772) );
  AND2_X1 U479 ( .A1(n586), .A2(n585), .ZN(n580) );
  XNOR2_X1 U480 ( .A(n564), .B(KEYINPUT98), .ZN(n679) );
  XNOR2_X1 U481 ( .A(n470), .B(n468), .ZN(n742) );
  XNOR2_X1 U482 ( .A(n741), .B(n469), .ZN(n468) );
  INV_X1 U483 ( .A(KEYINPUT56), .ZN(n379) );
  XNOR2_X1 U484 ( .A(n437), .B(n436), .ZN(G75) );
  XNOR2_X1 U485 ( .A(n732), .B(KEYINPUT119), .ZN(n436) );
  NAND2_X1 U486 ( .A1(n730), .A2(n438), .ZN(n437) );
  AND2_X1 U487 ( .A1(n687), .A2(n367), .ZN(n358) );
  XOR2_X1 U488 ( .A(n528), .B(KEYINPUT25), .Z(n359) );
  NOR2_X1 U489 ( .A1(n573), .A2(n568), .ZN(n360) );
  XOR2_X1 U490 ( .A(G146), .B(n545), .Z(n361) );
  XOR2_X1 U491 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n362) );
  AND2_X1 U492 ( .A1(n430), .A2(n429), .ZN(n363) );
  XOR2_X1 U493 ( .A(G131), .B(G134), .Z(n364) );
  AND2_X1 U494 ( .A1(n622), .A2(n446), .ZN(n365) );
  AND2_X1 U495 ( .A1(n353), .A2(n464), .ZN(n366) );
  AND2_X1 U496 ( .A1(n516), .A2(n609), .ZN(n367) );
  XOR2_X1 U497 ( .A(n491), .B(KEYINPUT65), .Z(n368) );
  XOR2_X1 U498 ( .A(KEYINPUT89), .B(n655), .Z(n743) );
  INV_X1 U499 ( .A(n743), .ZN(n478) );
  XOR2_X1 U500 ( .A(n422), .B(n733), .Z(n369) );
  XOR2_X1 U501 ( .A(n511), .B(KEYINPUT62), .Z(n370) );
  XOR2_X1 U502 ( .A(n658), .B(n657), .Z(n371) );
  XOR2_X1 U503 ( .A(n736), .B(n735), .Z(n372) );
  NAND2_X1 U504 ( .A1(n368), .A2(n419), .ZN(n373) );
  INV_X1 U505 ( .A(n418), .ZN(n406) );
  NOR2_X1 U506 ( .A1(n368), .A2(n419), .ZN(n418) );
  INV_X1 U507 ( .A(KEYINPUT64), .ZN(n419) );
  BUF_X1 U508 ( .A(n693), .Z(n374) );
  BUF_X1 U509 ( .A(n717), .Z(n375) );
  XNOR2_X1 U510 ( .A(n627), .B(n626), .ZN(n717) );
  XNOR2_X1 U511 ( .A(n591), .B(KEYINPUT40), .ZN(n376) );
  BUF_X1 U512 ( .A(n605), .Z(n377) );
  XNOR2_X1 U513 ( .A(n591), .B(KEYINPUT40), .ZN(n774) );
  NAND2_X1 U514 ( .A1(n605), .A2(n677), .ZN(n591) );
  XNOR2_X1 U515 ( .A(n590), .B(n589), .ZN(n605) );
  NAND2_X1 U516 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U517 ( .A(n772), .B(n378), .ZN(n583) );
  XNOR2_X1 U518 ( .A(n380), .B(n379), .ZN(G51) );
  NAND2_X1 U519 ( .A1(n420), .A2(n478), .ZN(n380) );
  XNOR2_X1 U520 ( .A(n423), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U521 ( .A1(n424), .A2(n478), .ZN(n423) );
  XNOR2_X1 U522 ( .A(n425), .B(n370), .ZN(n424) );
  NOR2_X1 U523 ( .A1(n736), .A2(G902), .ZN(n538) );
  XNOR2_X1 U524 ( .A(n472), .B(n471), .ZN(n381) );
  BUF_X1 U525 ( .A(n402), .Z(n382) );
  NAND2_X2 U526 ( .A1(n612), .A2(n611), .ZN(n472) );
  XNOR2_X1 U527 ( .A(G116), .B(n356), .ZN(n495) );
  AND2_X2 U528 ( .A1(n441), .A2(n440), .ZN(n383) );
  AND2_X2 U529 ( .A1(n441), .A2(n440), .ZN(n403) );
  XNOR2_X2 U530 ( .A(n569), .B(KEYINPUT19), .ZN(n612) );
  NAND2_X1 U531 ( .A1(n770), .A2(KEYINPUT44), .ZN(n414) );
  BUF_X1 U532 ( .A(n560), .Z(n585) );
  NAND2_X1 U533 ( .A1(n384), .A2(n401), .ZN(n400) );
  NAND2_X1 U534 ( .A1(n398), .A2(n384), .ZN(n397) );
  INV_X2 U535 ( .A(G122), .ZN(n442) );
  INV_X1 U536 ( .A(n396), .ZN(n389) );
  NAND2_X1 U537 ( .A1(n396), .A2(n395), .ZN(n394) );
  AND2_X1 U538 ( .A1(n765), .A2(KEYINPUT83), .ZN(n395) );
  NAND2_X1 U539 ( .A1(n399), .A2(n397), .ZN(n441) );
  NOR2_X1 U540 ( .A1(n757), .A2(n419), .ZN(n398) );
  NAND2_X1 U541 ( .A1(n400), .A2(n405), .ZN(n399) );
  NAND2_X1 U542 ( .A1(n402), .A2(n653), .ZN(n654) );
  XNOR2_X2 U543 ( .A(n652), .B(n651), .ZN(n402) );
  NAND2_X1 U544 ( .A1(n402), .A2(KEYINPUT2), .ZN(n404) );
  NOR2_X1 U545 ( .A1(n382), .A2(n722), .ZN(n723) );
  NAND2_X1 U546 ( .A1(n382), .A2(n758), .ZN(n747) );
  NAND2_X1 U547 ( .A1(n403), .A2(G475), .ZN(n659) );
  NAND2_X1 U548 ( .A1(n403), .A2(G210), .ZN(n734) );
  NAND2_X1 U549 ( .A1(n383), .A2(G478), .ZN(n737) );
  NAND2_X1 U550 ( .A1(n403), .A2(G472), .ZN(n425) );
  NAND2_X1 U551 ( .A1(n383), .A2(G469), .ZN(n480) );
  NAND2_X1 U552 ( .A1(n383), .A2(G217), .ZN(n470) );
  XNOR2_X1 U553 ( .A(n407), .B(n439), .ZN(n474) );
  XNOR2_X2 U554 ( .A(n492), .B(n483), .ZN(n439) );
  XNOR2_X2 U555 ( .A(n482), .B(G128), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n547), .B(n408), .ZN(n407) );
  XNOR2_X1 U557 ( .A(n545), .B(KEYINPUT17), .ZN(n408) );
  XNOR2_X2 U558 ( .A(n453), .B(G101), .ZN(n545) );
  INV_X1 U559 ( .A(n770), .ZN(n416) );
  XNOR2_X2 U560 ( .A(n636), .B(n635), .ZN(n770) );
  NAND2_X1 U561 ( .A1(n417), .A2(KEYINPUT44), .ZN(n410) );
  NAND2_X1 U562 ( .A1(n671), .A2(n771), .ZN(n417) );
  NOR2_X1 U563 ( .A1(n411), .A2(n409), .ZN(n413) );
  NAND2_X1 U564 ( .A1(n410), .A2(n414), .ZN(n409) );
  NOR2_X1 U565 ( .A1(n417), .A2(n412), .ZN(n411) );
  NAND2_X1 U566 ( .A1(n416), .A2(n415), .ZN(n412) );
  NAND2_X1 U567 ( .A1(n413), .A2(n650), .ZN(n652) );
  NAND2_X1 U568 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U569 ( .A1(n435), .A2(n365), .ZN(n671) );
  XNOR2_X1 U570 ( .A(n734), .B(n369), .ZN(n420) );
  NOR2_X1 U571 ( .A1(n422), .A2(n653), .ZN(n552) );
  XNOR2_X1 U572 ( .A(n475), .B(n474), .ZN(n422) );
  NOR2_X1 U573 ( .A1(n621), .A2(n620), .ZN(n648) );
  NAND2_X1 U574 ( .A1(n363), .A2(n426), .ZN(n435) );
  INV_X1 U575 ( .A(n621), .ZN(n428) );
  NAND2_X1 U576 ( .A1(n621), .A2(KEYINPUT103), .ZN(n430) );
  NOR2_X2 U577 ( .A1(n621), .A2(n433), .ZN(n432) );
  XNOR2_X2 U578 ( .A(n442), .B(G104), .ZN(n542) );
  NOR2_X2 U579 ( .A1(n693), .A2(n577), .ZN(n641) );
  NAND2_X1 U580 ( .A1(n461), .A2(n687), .ZN(n693) );
  XNOR2_X1 U581 ( .A(n548), .B(n449), .ZN(n448) );
  NAND2_X1 U582 ( .A1(n445), .A2(n367), .ZN(n578) );
  XNOR2_X1 U583 ( .A(n641), .B(KEYINPUT106), .ZN(n445) );
  XNOR2_X1 U584 ( .A(n748), .B(n448), .ZN(n475) );
  NAND2_X1 U585 ( .A1(n447), .A2(n481), .ZN(n584) );
  XNOR2_X2 U586 ( .A(n616), .B(KEYINPUT22), .ZN(n621) );
  NOR2_X2 U587 ( .A1(n660), .A2(n743), .ZN(n663) );
  XNOR2_X1 U588 ( .A(n536), .B(n537), .ZN(n736) );
  NOR2_X1 U589 ( .A1(n680), .A2(n667), .ZN(n644) );
  XNOR2_X2 U590 ( .A(n755), .B(n361), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n679), .A2(n677), .ZN(n457) );
  XNOR2_X2 U592 ( .A(n510), .B(KEYINPUT97), .ZN(n677) );
  INV_X1 U593 ( .A(n473), .ZN(n461) );
  XNOR2_X2 U594 ( .A(n538), .B(G469), .ZN(n577) );
  XNOR2_X2 U595 ( .A(KEYINPUT1), .B(n577), .ZN(n692) );
  XNOR2_X2 U596 ( .A(G110), .B(G107), .ZN(n750) );
  NAND2_X1 U597 ( .A1(n532), .A2(n353), .ZN(n570) );
  NAND2_X1 U598 ( .A1(n532), .A2(n366), .ZN(n467) );
  INV_X1 U599 ( .A(n569), .ZN(n464) );
  NAND2_X1 U600 ( .A1(n465), .A2(n617), .ZN(n571) );
  NAND2_X1 U601 ( .A1(n642), .A2(n615), .ZN(n616) );
  XNOR2_X2 U602 ( .A(n472), .B(n471), .ZN(n642) );
  XNOR2_X1 U603 ( .A(n477), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U604 ( .A1(n479), .A2(n478), .ZN(n477) );
  XNOR2_X1 U605 ( .A(n480), .B(n372), .ZN(n479) );
  BUF_X2 U606 ( .A(n555), .Z(n690) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(n560) );
  AND2_X1 U608 ( .A1(n567), .A2(n566), .ZN(n481) );
  INV_X1 U609 ( .A(KEYINPUT67), .ZN(n602) );
  XNOR2_X1 U610 ( .A(G113), .B(G116), .ZN(n486) );
  XNOR2_X1 U611 ( .A(n602), .B(KEYINPUT48), .ZN(n603) );
  INV_X1 U612 ( .A(KEYINPUT86), .ZN(n624) );
  INV_X1 U613 ( .A(KEYINPUT4), .ZN(n483) );
  XNOR2_X1 U614 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U615 ( .A(n355), .B(n489), .ZN(n490) );
  XNOR2_X1 U616 ( .A(n535), .B(n548), .ZN(n536) );
  XNOR2_X1 U617 ( .A(n523), .B(n522), .ZN(n524) );
  AND2_X1 U618 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U619 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n589) );
  XNOR2_X1 U620 ( .A(n659), .B(n371), .ZN(n660) );
  XNOR2_X1 U621 ( .A(n634), .B(KEYINPUT82), .ZN(n635) );
  NAND2_X1 U622 ( .A1(n501), .A2(G210), .ZN(n484) );
  XOR2_X1 U623 ( .A(n485), .B(n484), .Z(n489) );
  INV_X1 U624 ( .A(n486), .ZN(n488) );
  NAND2_X1 U625 ( .A1(n653), .A2(KEYINPUT2), .ZN(n491) );
  XOR2_X1 U626 ( .A(n492), .B(G134), .Z(n494) );
  NAND2_X1 U627 ( .A1(G234), .A2(n758), .ZN(n493) );
  XOR2_X1 U628 ( .A(KEYINPUT8), .B(n493), .Z(n521) );
  XNOR2_X1 U629 ( .A(n496), .B(n495), .ZN(n497) );
  NOR2_X1 U630 ( .A1(n738), .A2(G902), .ZN(n498) );
  XNOR2_X1 U631 ( .A(n498), .B(G478), .ZN(n592) );
  XNOR2_X1 U632 ( .A(n500), .B(n499), .ZN(n507) );
  NAND2_X1 U633 ( .A1(G214), .A2(n501), .ZN(n502) );
  XNOR2_X1 U634 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U635 ( .A(n504), .B(n517), .Z(n506) );
  XNOR2_X1 U636 ( .A(n542), .B(G140), .ZN(n505) );
  NOR2_X1 U637 ( .A1(G902), .A2(n656), .ZN(n509) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(G475), .ZN(n508) );
  XNOR2_X1 U639 ( .A(n509), .B(n508), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n592), .A2(n576), .ZN(n510) );
  INV_X1 U641 ( .A(KEYINPUT6), .ZN(n512) );
  NOR2_X1 U642 ( .A1(G900), .A2(n758), .ZN(n513) );
  NAND2_X1 U643 ( .A1(n513), .A2(G902), .ZN(n514) );
  NAND2_X1 U644 ( .A1(G952), .A2(n758), .ZN(n607) );
  NAND2_X1 U645 ( .A1(n514), .A2(n607), .ZN(n516) );
  XNOR2_X1 U646 ( .A(n515), .B(KEYINPUT14), .ZN(n609) );
  XNOR2_X1 U647 ( .A(n756), .B(KEYINPUT23), .ZN(n525) );
  XOR2_X1 U648 ( .A(KEYINPUT24), .B(G110), .Z(n519) );
  XNOR2_X1 U649 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U650 ( .A(n520), .B(KEYINPUT91), .Z(n523) );
  AND2_X1 U651 ( .A1(n521), .A2(G221), .ZN(n522) );
  XNOR2_X1 U652 ( .A(n525), .B(n524), .ZN(n741) );
  NOR2_X1 U653 ( .A1(n741), .A2(G902), .ZN(n529) );
  INV_X1 U654 ( .A(n653), .ZN(n526) );
  NAND2_X1 U655 ( .A1(n526), .A2(G234), .ZN(n527) );
  XNOR2_X1 U656 ( .A(n527), .B(KEYINPUT20), .ZN(n530) );
  NAND2_X1 U657 ( .A1(n530), .A2(G217), .ZN(n528) );
  NAND2_X1 U658 ( .A1(n530), .A2(G221), .ZN(n531) );
  XOR2_X1 U659 ( .A(KEYINPUT21), .B(n531), .Z(n687) );
  INV_X1 U660 ( .A(n687), .ZN(n613) );
  NAND2_X1 U661 ( .A1(G227), .A2(n758), .ZN(n534) );
  XNOR2_X1 U662 ( .A(KEYINPUT68), .B(n750), .ZN(n548) );
  NAND2_X1 U663 ( .A1(G214), .A2(n550), .ZN(n701) );
  NAND2_X1 U664 ( .A1(n692), .A2(n701), .ZN(n539) );
  NOR2_X1 U665 ( .A1(n570), .A2(n539), .ZN(n541) );
  XNOR2_X1 U666 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n540) );
  XNOR2_X1 U667 ( .A(n541), .B(n540), .ZN(n553) );
  NAND2_X1 U668 ( .A1(G224), .A2(n758), .ZN(n546) );
  NAND2_X1 U669 ( .A1(G210), .A2(n550), .ZN(n551) );
  NOR2_X1 U670 ( .A1(n553), .A2(n585), .ZN(n554) );
  XNOR2_X1 U671 ( .A(n554), .B(KEYINPUT105), .ZN(n765) );
  XOR2_X1 U672 ( .A(KEYINPUT28), .B(n556), .Z(n559) );
  INV_X1 U673 ( .A(n577), .ZN(n557) );
  XOR2_X1 U674 ( .A(n557), .B(KEYINPUT108), .Z(n558) );
  NAND2_X1 U675 ( .A1(n560), .A2(n701), .ZN(n562) );
  XNOR2_X2 U676 ( .A(n562), .B(n561), .ZN(n569) );
  NAND2_X1 U677 ( .A1(n672), .A2(KEYINPUT47), .ZN(n563) );
  XNOR2_X1 U678 ( .A(n563), .B(KEYINPUT76), .ZN(n567) );
  NOR2_X1 U679 ( .A1(n592), .A2(n576), .ZN(n564) );
  NAND2_X1 U680 ( .A1(n565), .A2(KEYINPUT47), .ZN(n566) );
  INV_X1 U681 ( .A(KEYINPUT71), .ZN(n568) );
  XNOR2_X1 U682 ( .A(n692), .B(KEYINPUT87), .ZN(n617) );
  XNOR2_X1 U683 ( .A(n571), .B(KEYINPUT110), .ZN(n766) );
  NOR2_X1 U684 ( .A1(KEYINPUT47), .A2(KEYINPUT71), .ZN(n572) );
  NAND2_X1 U685 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U686 ( .A1(n766), .A2(n574), .ZN(n575) );
  INV_X1 U687 ( .A(n576), .ZN(n593) );
  NOR2_X1 U688 ( .A1(n593), .A2(n592), .ZN(n631) );
  INV_X1 U689 ( .A(KEYINPUT30), .ZN(n579) );
  NAND2_X1 U690 ( .A1(n631), .A2(n581), .ZN(n582) );
  NOR2_X1 U691 ( .A1(n584), .A2(n583), .ZN(n601) );
  NAND2_X1 U692 ( .A1(n588), .A2(n587), .ZN(n590) );
  XOR2_X1 U693 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n597) );
  NAND2_X1 U694 ( .A1(n593), .A2(n592), .ZN(n704) );
  XOR2_X1 U695 ( .A(KEYINPUT41), .B(n594), .Z(n685) );
  NAND2_X1 U696 ( .A1(n595), .A2(n685), .ZN(n596) );
  NAND2_X1 U697 ( .A1(n774), .A2(n775), .ZN(n599) );
  INV_X1 U698 ( .A(KEYINPUT46), .ZN(n598) );
  XNOR2_X1 U699 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U700 ( .A1(n377), .A2(n679), .ZN(n684) );
  NOR2_X1 U701 ( .A1(G898), .A2(n758), .ZN(n606) );
  XNOR2_X1 U702 ( .A(KEYINPUT90), .B(n606), .ZN(n751) );
  NAND2_X1 U703 ( .A1(n751), .A2(G902), .ZN(n608) );
  NAND2_X1 U704 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U705 ( .A(n609), .ZN(n714) );
  NOR2_X1 U706 ( .A1(n613), .A2(n704), .ZN(n614) );
  XNOR2_X1 U707 ( .A(KEYINPUT100), .B(n614), .ZN(n615) );
  INV_X1 U708 ( .A(n623), .ZN(n646) );
  AND2_X1 U709 ( .A1(n646), .A2(n617), .ZN(n618) );
  INV_X1 U710 ( .A(n619), .ZN(n622) );
  INV_X1 U711 ( .A(n692), .ZN(n620) );
  INV_X1 U712 ( .A(KEYINPUT34), .ZN(n630) );
  INV_X1 U713 ( .A(n642), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n637), .A2(n623), .ZN(n627) );
  XOR2_X1 U715 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n625) );
  XNOR2_X1 U716 ( .A(n630), .B(n629), .ZN(n633) );
  INV_X1 U717 ( .A(n631), .ZN(n632) );
  NOR2_X2 U718 ( .A1(n633), .A2(n632), .ZN(n636) );
  XOR2_X1 U719 ( .A(KEYINPUT93), .B(KEYINPUT31), .Z(n640) );
  AND2_X1 U720 ( .A1(n637), .A2(n690), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(KEYINPUT92), .ZN(n697) );
  NAND2_X1 U722 ( .A1(n697), .A2(n381), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n381), .A2(n641), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n690), .A2(n643), .ZN(n667) );
  XNOR2_X1 U725 ( .A(n644), .B(KEYINPUT94), .ZN(n645) );
  OR2_X1 U726 ( .A1(n706), .A2(n645), .ZN(n649) );
  AND2_X1 U727 ( .A1(n646), .A2(n686), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n664) );
  AND2_X1 U729 ( .A1(n649), .A2(n664), .ZN(n650) );
  NOR2_X1 U730 ( .A1(G952), .A2(n758), .ZN(n655) );
  XNOR2_X1 U731 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n656), .B(KEYINPUT88), .ZN(n657) );
  INV_X1 U733 ( .A(KEYINPUT60), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT123), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G60) );
  XNOR2_X1 U736 ( .A(G101), .B(n664), .ZN(G3) );
  XOR2_X1 U737 ( .A(G104), .B(KEYINPUT111), .Z(n666) );
  NAND2_X1 U738 ( .A1(n667), .A2(n677), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n669) );
  NAND2_X1 U741 ( .A1(n667), .A2(n679), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U743 ( .A(G107), .B(n670), .ZN(G9) );
  XNOR2_X1 U744 ( .A(n671), .B(G110), .ZN(G12) );
  XOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .Z(n674) );
  INV_X1 U746 ( .A(n672), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n675), .A2(n679), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n674), .B(n673), .ZN(G30) );
  NAND2_X1 U749 ( .A1(n675), .A2(n677), .ZN(n676) );
  XNOR2_X1 U750 ( .A(n676), .B(G146), .ZN(G48) );
  NAND2_X1 U751 ( .A1(n354), .A2(n677), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n678), .B(G113), .ZN(G15) );
  XOR2_X1 U753 ( .A(G116), .B(KEYINPUT113), .Z(n682) );
  NAND2_X1 U754 ( .A1(n354), .A2(n679), .ZN(n681) );
  XNOR2_X1 U755 ( .A(n682), .B(n681), .ZN(G18) );
  XOR2_X1 U756 ( .A(G134), .B(KEYINPUT115), .Z(n683) );
  XNOR2_X1 U757 ( .A(n684), .B(n683), .ZN(G36) );
  INV_X1 U758 ( .A(n685), .ZN(n718) );
  NOR2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U760 ( .A(KEYINPUT49), .B(n688), .Z(n689) );
  NOR2_X1 U761 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U762 ( .A(KEYINPUT116), .B(n691), .Z(n696) );
  AND2_X1 U763 ( .A1(n374), .A2(n692), .ZN(n694) );
  XNOR2_X1 U764 ( .A(KEYINPUT50), .B(n694), .ZN(n695) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U767 ( .A(KEYINPUT51), .B(n699), .Z(n700) );
  NOR2_X1 U768 ( .A1(n718), .A2(n700), .ZN(n711) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n375), .A2(n709), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U775 ( .A(n712), .B(KEYINPUT52), .ZN(n713) );
  NOR2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U777 ( .A1(G952), .A2(n715), .ZN(n716) );
  XNOR2_X1 U778 ( .A(n716), .B(KEYINPUT117), .ZN(n720) );
  NOR2_X1 U779 ( .A1(n718), .A2(n375), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U781 ( .A(n721), .B(KEYINPUT118), .ZN(n731) );
  XNOR2_X1 U782 ( .A(KEYINPUT2), .B(KEYINPUT75), .ZN(n726) );
  INV_X1 U783 ( .A(n726), .ZN(n722) );
  XNOR2_X1 U784 ( .A(n723), .B(KEYINPUT78), .ZN(n724) );
  NOR2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n729) );
  NAND2_X1 U786 ( .A1(n726), .A2(n757), .ZN(n727) );
  XOR2_X1 U787 ( .A(KEYINPUT79), .B(n727), .Z(n728) );
  NAND2_X1 U788 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U789 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n732) );
  XOR2_X1 U790 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n733) );
  XOR2_X1 U791 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n735) );
  XNOR2_X1 U792 ( .A(n737), .B(KEYINPUT124), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n743), .A2(n740), .ZN(G63) );
  NOR2_X1 U795 ( .A1(n743), .A2(n742), .ZN(G66) );
  NAND2_X1 U796 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U798 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n754) );
  XOR2_X1 U800 ( .A(n357), .B(G101), .Z(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(n752) );
  NOR2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(G69) );
  XNOR2_X1 U804 ( .A(n756), .B(n755), .ZN(n760) );
  XNOR2_X1 U805 ( .A(n757), .B(n760), .ZN(n759) );
  NAND2_X1 U806 ( .A1(n759), .A2(n758), .ZN(n764) );
  XNOR2_X1 U807 ( .A(G227), .B(n760), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(G953), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n764), .A2(n763), .ZN(G72) );
  XNOR2_X1 U811 ( .A(G140), .B(n765), .ZN(G42) );
  XOR2_X1 U812 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n768) );
  XNOR2_X1 U813 ( .A(n766), .B(G125), .ZN(n767) );
  XNOR2_X1 U814 ( .A(n768), .B(n767), .ZN(G27) );
  XOR2_X1 U815 ( .A(n356), .B(KEYINPUT126), .Z(n769) );
  XNOR2_X1 U816 ( .A(n770), .B(n769), .ZN(G24) );
  XNOR2_X1 U817 ( .A(n771), .B(G119), .ZN(G21) );
  XOR2_X1 U818 ( .A(G143), .B(n772), .Z(n773) );
  XNOR2_X1 U819 ( .A(KEYINPUT112), .B(n773), .ZN(G45) );
  XNOR2_X1 U820 ( .A(n376), .B(G131), .ZN(G33) );
  XOR2_X1 U821 ( .A(G137), .B(n775), .Z(n776) );
  XNOR2_X1 U822 ( .A(KEYINPUT127), .B(n776), .ZN(G39) );
endmodule

