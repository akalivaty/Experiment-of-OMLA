//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(new_n458), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  OR2_X1    g044(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(G136), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n462), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n476), .B1(new_n478), .B2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(KEYINPUT69), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n458), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n477), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n463), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n462), .A2(new_n492), .A3(G138), .A4(new_n458), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G88), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(G50), .A3(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(G62), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n506), .B1(new_n511), .B2(G651), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  AOI211_X1 g088(.A(KEYINPUT71), .B(new_n513), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n504), .A2(new_n505), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  OAI221_X1 g092(.A(new_n517), .B1(new_n512), .B2(new_n514), .C1(new_n504), .C2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT73), .B(G89), .Z(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(new_n499), .A3(new_n500), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n496), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  AND4_X1   g103(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n528), .ZN(G168));
  OAI21_X1  g104(.A(G64), .B1(new_n507), .B2(new_n508), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n513), .B1(new_n530), .B2(new_n531), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT74), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n525), .A2(new_n526), .B1(new_n497), .B2(new_n498), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G90), .B1(new_n527), .B2(G52), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n497), .B2(new_n498), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT75), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n507), .A2(new_n508), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n547), .B(new_n544), .C1(new_n548), .C2(new_n542), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(G651), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n538), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n548), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n564));
  AND2_X1   g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT6), .A2(G651), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n500), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n568), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n564), .B1(new_n572), .B2(new_n573), .ZN(G299));
  NAND4_X1  g149(.A1(new_n523), .A2(new_n528), .A3(new_n521), .A4(new_n524), .ZN(G286));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND2_X1  g151(.A1(G166), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G303));
  NAND2_X1  g154(.A1(new_n538), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n581));
  INV_X1    g156(.A(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G543), .B1(new_n565), .B2(new_n566), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(G288));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n548), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n499), .A2(new_n587), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G48), .B2(new_n527), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n538), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n499), .A2(G60), .ZN(new_n594));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n513), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT81), .B(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n538), .A2(G85), .B1(new_n527), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n583), .B2(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n548), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n604), .A2(new_n606), .B1(new_n609), .B2(G651), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n499), .A2(new_n500), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n603), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n603), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G280));
  XOR2_X1   g198(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n618), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n555), .ZN(G323));
  XOR2_X1   g204(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  NAND2_X1  g206(.A1(new_n462), .A2(new_n460), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2100), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n470), .A2(new_n471), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G135), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n458), .A2(G111), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(KEYINPUT85), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(KEYINPUT85), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n478), .A2(G123), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n635), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(G2096), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n636), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT88), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n666), .A3(new_n669), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n668), .A2(new_n670), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n666), .A2(new_n669), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n677), .A2(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n673), .B(new_n675), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT20), .Z(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT90), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n697), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G27), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT103), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n491), .A2(new_n493), .ZN(new_n706));
  INV_X1    g281(.A(new_n489), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n705), .B1(new_n708), .B2(G29), .ZN(new_n709));
  INV_X1    g284(.A(G2078), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NOR2_X1   g287(.A1(G171), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G5), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1961), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G34), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(KEYINPUT24), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(KEYINPUT24), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n703), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G160), .B2(new_n703), .ZN(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n703), .A2(G33), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT99), .B(KEYINPUT25), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n458), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n637), .B2(G139), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n703), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n716), .B(new_n723), .C1(G2072), .C2(new_n731), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n711), .B(new_n732), .C1(G2072), .C2(new_n731), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT30), .B(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n734), .A2(new_n703), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n644), .B2(new_n703), .ZN(new_n738));
  NOR2_X1   g313(.A1(G168), .A2(new_n712), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n712), .B2(G21), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(G1966), .B2(new_n741), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n742), .B1(new_n715), .B2(new_n714), .C1(G1966), .C2(new_n741), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT102), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT102), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n703), .A2(G32), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n470), .A2(G141), .A3(new_n471), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT100), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n460), .A2(G105), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n749), .B(new_n752), .C1(G129), .C2(new_n478), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n703), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n733), .A2(new_n744), .A3(new_n745), .A4(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT104), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n712), .A2(G20), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT106), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT23), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n622), .B2(new_n712), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n703), .A2(G26), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT98), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G128), .B2(new_n478), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n470), .A2(G140), .A3(new_n471), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2067), .ZN(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n618), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT97), .B(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n555), .A2(new_n712), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n712), .B2(G19), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n777), .B(new_n781), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n767), .B(new_n785), .C1(new_n782), .C2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n703), .A2(G35), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G162), .B2(new_n703), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n789));
  INV_X1    g364(.A(G2090), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n788), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n761), .A2(new_n762), .A3(new_n786), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G22), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G166), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n712), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(G288), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n712), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT33), .B(G1976), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n712), .A2(G6), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G305), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT32), .B(G1981), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n803), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n797), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n703), .A2(G25), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n470), .A2(G131), .A3(new_n471), .ZN(new_n814));
  NOR2_X1   g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT92), .ZN(new_n816));
  INV_X1    g391(.A(G2104), .ZN(new_n817));
  INV_X1    g392(.A(G107), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n478), .A2(G119), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n813), .B1(new_n822), .B2(new_n703), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G1991), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT93), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(KEYINPUT93), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n712), .A2(G24), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G290), .B2(G16), .ZN(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n812), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(KEYINPUT96), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n793), .B1(new_n840), .B2(new_n842), .ZN(G311));
  INV_X1    g418(.A(new_n793), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n841), .B1(new_n835), .B2(new_n836), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(G150));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n612), .A2(new_n848), .B1(new_n849), .B2(new_n583), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  INV_X1    g426(.A(G80), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n548), .A2(new_n851), .B1(new_n852), .B2(new_n496), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n513), .B1(new_n853), .B2(KEYINPUT107), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT107), .ZN(new_n855));
  OAI221_X1 g430(.A(new_n855), .B1(new_n852), .B2(new_n496), .C1(new_n548), .C2(new_n851), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n850), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G860), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n550), .A2(new_n552), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT76), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n550), .A2(new_n552), .A3(new_n551), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n854), .A2(new_n856), .ZN(new_n865));
  INV_X1    g440(.A(new_n850), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n861), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n617), .A2(new_n625), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT108), .Z(new_n875));
  OAI21_X1  g450(.A(new_n858), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n860), .B1(new_n875), .B2(new_n876), .ZN(G145));
  AND3_X1   g452(.A1(new_n748), .A2(new_n753), .A3(new_n730), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n730), .B1(new_n748), .B2(new_n753), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n814), .A2(KEYINPUT110), .A3(new_n820), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT110), .B1(new_n814), .B2(new_n820), .ZN(new_n882));
  INV_X1    g457(.A(new_n633), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n885), .B(new_n884), .C1(new_n878), .C2(new_n879), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n775), .A2(new_n708), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n637), .A2(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n478), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n458), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n773), .A2(G164), .A3(new_n774), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n890), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n890), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n889), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n887), .A2(new_n899), .A3(new_n888), .ZN(new_n902));
  INV_X1    g477(.A(new_n644), .ZN(new_n903));
  XOR2_X1   g478(.A(G160), .B(KEYINPUT109), .Z(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n482), .B2(new_n483), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n482), .A2(new_n483), .A3(new_n905), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n910), .A2(new_n644), .A3(new_n906), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n901), .B(new_n902), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n644), .B1(new_n910), .B2(new_n906), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n887), .A2(new_n888), .A3(new_n899), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n899), .B1(new_n887), .B2(new_n888), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g495(.A(new_n869), .B(new_n627), .ZN(new_n921));
  AND2_X1   g496(.A1(G299), .A2(new_n617), .ZN(new_n922));
  NOR2_X1   g497(.A1(G299), .A2(new_n617), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n922), .B2(new_n923), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n622), .A2(new_n618), .ZN(new_n930));
  NAND2_X1  g505(.A1(G299), .A2(new_n617), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT41), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n921), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n926), .B(new_n927), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT42), .B1(new_n936), .B2(new_n925), .ZN(new_n937));
  NAND2_X1  g512(.A1(G166), .A2(new_n799), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n516), .A2(new_n518), .A3(G288), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(G305), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(G305), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n939), .A3(new_n938), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n935), .A2(new_n937), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n935), .B2(new_n937), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n857), .A2(G868), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(G295));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n951), .ZN(G331));
  XNOR2_X1  g530(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n538), .A2(G90), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n527), .A2(G52), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n957), .B(new_n958), .C1(new_n536), .C2(KEYINPUT74), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n533), .A2(new_n534), .ZN(new_n960));
  OAI21_X1  g535(.A(G168), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n535), .A2(G286), .A3(new_n537), .A4(new_n539), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n864), .A2(new_n868), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n867), .B1(new_n553), .B2(new_n554), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n857), .A2(new_n550), .A3(new_n552), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n965), .A2(new_n966), .B1(new_n961), .B2(new_n962), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n924), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n864), .B2(new_n868), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n965), .A2(new_n966), .A3(new_n961), .A4(new_n962), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n929), .A4(new_n932), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT113), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n964), .A2(new_n967), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n933), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n946), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(KEYINPUT114), .A3(new_n918), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n971), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n973), .ZN(new_n979));
  INV_X1    g554(.A(new_n946), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT114), .B1(new_n976), .B2(new_n918), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n978), .A2(new_n946), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n978), .B2(new_n946), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n918), .A4(new_n982), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n956), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n976), .A2(new_n918), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(new_n990), .A3(new_n982), .A4(new_n977), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n982), .B(new_n918), .C1(new_n988), .C2(new_n987), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(KEYINPUT43), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT116), .B1(new_n992), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n999), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n995), .A2(new_n982), .A3(new_n977), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1002), .B(new_n1003), .C1(new_n1006), .C2(new_n956), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1001), .A2(new_n1007), .ZN(G397));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(G40), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n465), .A2(new_n468), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1996), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n754), .B(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n775), .A2(G2067), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n775), .A2(G2067), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n822), .A2(new_n824), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n822), .A2(new_n824), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n941), .A2(new_n830), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G290), .A2(G1986), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1014), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1966), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n706), .B2(new_n707), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1012), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G164), .A2(new_n1009), .A3(G1384), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n722), .A4(new_n1012), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(G168), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT125), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT51), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n1037), .A2(KEYINPUT51), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1036), .A2(G8), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(G8), .A3(G286), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1036), .A2(G8), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(new_n1042), .C1(new_n1043), .C2(new_n1038), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1028), .B2(new_n1012), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n799), .A2(G1976), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G288), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1050), .A2(new_n1046), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G305), .A2(G1981), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT118), .B(G86), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n538), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n591), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n1058), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1048), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1056), .A2(new_n1057), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n1068));
  AOI211_X1 g643(.A(new_n1068), .B(new_n1047), .C1(new_n577), .C2(new_n578), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G303), .A2(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1068), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1384), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n708), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1013), .B1(new_n1075), .B2(new_n1009), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1028), .A2(KEYINPUT45), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n796), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1033), .A2(new_n1034), .A3(new_n1012), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(G2090), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1047), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1067), .B1(new_n1073), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1072), .A3(new_n1070), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1078), .B2(G2078), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1080), .A2(new_n715), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n710), .A4(new_n1077), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1045), .A2(new_n1083), .A3(new_n1085), .A4(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT126), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1067), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1082), .B1(new_n1097), .B2(new_n1069), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1085), .A2(new_n1044), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1087), .A2(G301), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1091), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT54), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1091), .A2(new_n1103), .A3(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1076), .A2(new_n1077), .A3(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT121), .B(G1956), .Z(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1080), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n568), .A2(new_n570), .ZN(new_n1112));
  INV_X1    g687(.A(new_n564), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(KEYINPUT57), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(new_n1114), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1108), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1106), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1077), .A2(new_n1010), .A3(new_n1015), .A4(new_n1012), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1028), .A2(new_n1012), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n555), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(new_n555), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1108), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT61), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1118), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1348), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1080), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1120), .A2(new_n1134), .A3(G2067), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1120), .B2(G2067), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1133), .A2(new_n1135), .A3(KEYINPUT60), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n617), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n617), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1139), .A2(new_n1140), .B1(new_n1138), .B2(new_n1137), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1131), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1129), .A2(new_n1142), .A3(new_n618), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1115), .B(KEYINPUT123), .Z(new_n1147));
  AND2_X1   g722(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1099), .B(new_n1105), .C1(new_n1145), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1098), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1066), .A2(new_n1053), .A3(new_n799), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(G1981), .B2(G305), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1151), .A2(new_n1096), .B1(new_n1153), .B2(new_n1048), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n1085), .A2(new_n1096), .A3(new_n1092), .A4(new_n1098), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1094), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1045), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1095), .A2(new_n1150), .A3(new_n1154), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1084), .A2(KEYINPUT120), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1082), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1160), .A2(new_n1162), .A3(new_n1072), .A4(new_n1070), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1047), .B(G286), .C1(new_n1031), .C2(new_n1035), .ZN(new_n1164));
  AND4_X1   g739(.A1(KEYINPUT63), .A2(new_n1163), .A3(new_n1083), .A4(new_n1164), .ZN(new_n1165));
  AND4_X1   g740(.A1(new_n1085), .A2(new_n1096), .A3(new_n1098), .A4(new_n1164), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1166), .A2(KEYINPUT119), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n1166), .B2(KEYINPUT119), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1026), .B1(new_n1159), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1022), .A2(new_n1014), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1014), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n1023), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT48), .Z(new_n1174));
  AND2_X1   g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT46), .Z(new_n1177));
  AOI21_X1  g752(.A(new_n1172), .B1(new_n1019), .B2(new_n755), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1017), .B1(new_n1181), .B2(new_n1021), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1175), .B(new_n1180), .C1(new_n1014), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1170), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n681), .A2(G319), .A3(new_n664), .ZN(new_n1187));
  NOR2_X1   g761(.A1(G229), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n919), .A2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g763(.A(new_n1186), .B(new_n1189), .C1(new_n985), .C2(new_n991), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n985), .A2(new_n991), .ZN(new_n1191));
  INV_X1    g765(.A(new_n1189), .ZN(new_n1192));
  AOI21_X1  g766(.A(KEYINPUT127), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1190), .A2(new_n1193), .ZN(G308));
  OAI21_X1  g768(.A(new_n1186), .B1(new_n1006), .B2(new_n1189), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1191), .A2(KEYINPUT127), .A3(new_n1192), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(G225));
endmodule


