//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND4_X1  g0008(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT66), .Z(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR3_X1   g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n210), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NOR4_X1   g0022(.A1(new_n213), .A2(new_n215), .A3(new_n219), .A4(new_n222), .ZN(G361));
  XNOR2_X1  g0023(.A(G250), .B(G257), .ZN(new_n224));
  XNOR2_X1  g0024(.A(G264), .B(G270), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n227), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XNOR2_X1  g0033(.A(G107), .B(G116), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(G50), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G68), .ZN(new_n237));
  INV_X1    g0037(.A(G68), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n235), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n218), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G58), .ZN(new_n254));
  OR3_X1    g0054(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT8), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n257), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(G20), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT76), .B1(new_n266), .B2(KEYINPUT7), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT76), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n268), .B(new_n269), .C1(new_n270), .C2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(KEYINPUT7), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G68), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n254), .A2(new_n238), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G58), .A2(G68), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n217), .A2(new_n262), .A3(G159), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT16), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT75), .B1(new_n266), .B2(KEYINPUT7), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT75), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n284), .B(new_n269), .C1(new_n270), .C2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n272), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G68), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n280), .A2(KEYINPUT16), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n246), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n261), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n263), .A2(new_n265), .A3(G226), .A4(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n263), .A2(new_n265), .A3(G223), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G87), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT77), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT77), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n291), .A2(new_n293), .A3(new_n297), .A4(new_n294), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n247), .A2(G274), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT68), .B(G45), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n262), .C2(new_n304), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(G232), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n300), .A2(new_n301), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n295), .B2(KEYINPUT77), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n313), .B2(new_n298), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(G200), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT17), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(KEYINPUT79), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n290), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n287), .A2(new_n288), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n279), .B1(new_n273), .B2(G68), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n245), .C1(KEYINPUT16), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n261), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n269), .B(G20), .C1(new_n263), .C2(new_n265), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n269), .B1(new_n270), .B2(G20), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(KEYINPUT75), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n238), .B1(new_n331), .B2(new_n285), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n280), .A2(KEYINPUT16), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n245), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n323), .B1(new_n334), .B2(new_n281), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n300), .A2(G179), .A3(new_n311), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n300), .B2(new_n311), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT78), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n300), .A2(new_n311), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G169), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n314), .A2(G179), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n335), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT18), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n335), .A2(new_n339), .A3(new_n344), .A4(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n328), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n270), .A2(G222), .A3(new_n292), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n270), .A2(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G223), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n351), .B1(new_n352), .B2(new_n270), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n299), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n307), .A2(new_n308), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n305), .B1(new_n358), .B2(G226), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(G179), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n258), .A2(new_n217), .A3(G1), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n236), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n249), .B2(new_n236), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n202), .A2(G20), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n217), .A2(new_n262), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n217), .A2(G33), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n365), .B1(new_n366), .B2(new_n367), .C1(new_n256), .C2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n364), .B1(new_n369), .B2(new_n245), .ZN(new_n370));
  AOI21_X1  g0170(.A(G169), .B1(new_n356), .B2(new_n359), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n361), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n360), .A2(new_n301), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G200), .B2(new_n360), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT9), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n370), .A2(new_n375), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT10), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n374), .B(new_n380), .C1(new_n376), .C2(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n372), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n263), .A2(new_n265), .A3(G232), .A4(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT72), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n270), .A2(new_n385), .A3(G232), .A4(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n263), .A2(new_n265), .A3(G226), .A4(new_n292), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n307), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n305), .B1(new_n358), .B2(G238), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT13), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n390), .B1(new_n386), .B2(new_n384), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n393), .B(new_n396), .C1(new_n397), .C2(new_n307), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n301), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n260), .A2(new_n401), .ZN(new_n402));
  AND4_X1   g0202(.A1(KEYINPUT70), .A2(new_n247), .A3(G13), .A4(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n404), .A3(new_n238), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT12), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n217), .A2(G68), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT12), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n259), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT73), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n245), .B1(new_n402), .B2(new_n404), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n238), .B1(new_n247), .B2(G20), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT74), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n406), .A2(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT74), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n407), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n368), .B2(new_n352), .C1(new_n236), .C2(new_n367), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n245), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n395), .B2(new_n398), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n400), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n399), .A2(G169), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n395), .A2(new_n398), .A3(G179), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n399), .A2(new_n430), .A3(G169), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n426), .B1(new_n432), .B2(new_n423), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G20), .A2(G77), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(new_n251), .B2(new_n367), .C1(new_n368), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n245), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n402), .A2(new_n404), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n438), .A2(G77), .A3(new_n246), .A4(new_n248), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n437), .B(new_n439), .C1(G77), .C2(new_n438), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n270), .A2(G232), .A3(new_n292), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  INV_X1    g0245(.A(G238), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n444), .B1(new_n445), .B2(new_n270), .C1(new_n353), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n299), .ZN(new_n448));
  INV_X1    g0248(.A(G244), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n306), .B1(new_n449), .B2(new_n357), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G179), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n447), .B2(new_n299), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G169), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n443), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(G200), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(G190), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  AND4_X1   g0265(.A1(new_n350), .A2(new_n382), .A3(new_n433), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n260), .A2(G97), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n246), .B(new_n260), .C1(G1), .C2(new_n262), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G97), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n445), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  XNOR2_X1  g0272(.A(G97), .B(G107), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT6), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n475), .A2(new_n217), .B1(new_n352), .B2(new_n367), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n273), .B2(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n471), .B1(new_n477), .B2(new_n246), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(KEYINPUT80), .B(new_n471), .C1(new_n477), .C2(new_n246), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n247), .B(G45), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n307), .A3(G257), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n247), .A2(G45), .ZN(new_n486));
  OR2_X1    g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G274), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(new_n292), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n498), .B2(new_n299), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n301), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(G200), .B2(new_n499), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n480), .A2(new_n481), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n486), .A2(G250), .ZN(new_n503));
  INV_X1    g0303(.A(G45), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n299), .A2(new_n503), .B1(new_n504), .B2(new_n302), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n270), .A2(G244), .A3(G1698), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n263), .A2(new_n265), .A3(G238), .A4(new_n292), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n509), .B2(new_n299), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n424), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(G190), .B2(new_n510), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n217), .B1(new_n389), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G87), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n445), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n263), .A2(new_n265), .A3(new_n217), .A4(G68), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n513), .B1(new_n368), .B2(new_n516), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n245), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n402), .A2(new_n404), .A3(new_n435), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT82), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(KEYINPUT82), .A3(new_n523), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n526), .A2(new_n527), .B1(G87), .B2(new_n470), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n469), .A2(new_n435), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n527), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT82), .B1(new_n522), .B2(new_n523), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n509), .A2(new_n299), .ZN(new_n534));
  INV_X1    g0334(.A(new_n505), .ZN(new_n535));
  AOI21_X1  g0335(.A(G169), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g0336(.A(G179), .B(new_n505), .C1(new_n509), .C2(new_n299), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n512), .A2(new_n528), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n498), .A2(new_n299), .ZN(new_n540));
  INV_X1    g0340(.A(new_n491), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(G179), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n337), .B2(new_n499), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(new_n478), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n543), .B2(new_n478), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n502), .B(new_n539), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n270), .A2(new_n217), .A3(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n270), .A2(new_n550), .A3(new_n217), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT23), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n445), .A3(G20), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT23), .B1(new_n217), .B2(G107), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT85), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n554), .B1(G20), .B2(new_n507), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g0360(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n552), .A2(new_n561), .A3(new_n559), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n246), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n362), .A2(new_n445), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT25), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n469), .A2(new_n445), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n484), .A2(new_n307), .A3(G264), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n490), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n263), .A2(new_n265), .A3(G250), .A4(new_n292), .ZN(new_n574));
  INV_X1    g0374(.A(G294), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n262), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n299), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n572), .B1(new_n577), .B2(KEYINPUT86), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT86), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n579), .A3(new_n299), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n337), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n490), .A3(new_n571), .ZN(new_n582));
  INV_X1    g0382(.A(G179), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n565), .A2(new_n570), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n489), .A2(new_n299), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(G270), .B1(G274), .B2(new_n489), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n263), .A2(new_n265), .A3(G264), .A4(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(new_n292), .ZN(new_n589));
  INV_X1    g0389(.A(G303), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n270), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n299), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n402), .A2(new_n404), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n247), .B2(G33), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT70), .B1(new_n259), .B2(G20), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n246), .B(new_n596), .C1(new_n597), .C2(new_n403), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n244), .A2(new_n218), .B1(G20), .B2(new_n594), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n496), .B(new_n217), .C1(G33), .C2(new_n516), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT20), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n595), .B(new_n598), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n593), .A2(new_n603), .A3(KEYINPUT21), .A4(G169), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(G179), .A3(new_n592), .A4(new_n587), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n337), .B1(new_n587), .B2(new_n592), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT21), .B1(new_n607), .B2(new_n603), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n603), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT83), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n587), .A2(new_n592), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n424), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n424), .B1(new_n587), .B2(new_n592), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT83), .B1(new_n614), .B2(new_n603), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(G190), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n577), .A2(KEYINPUT86), .ZN(new_n618));
  INV_X1    g0418(.A(new_n572), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n301), .A3(new_n580), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n582), .A2(new_n424), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n552), .A2(new_n561), .A3(new_n559), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n561), .B1(new_n552), .B2(new_n559), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n245), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n625), .A3(new_n569), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n585), .A2(new_n609), .A3(new_n617), .A4(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n467), .A2(new_n547), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT87), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n341), .A2(new_n343), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n335), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(new_n347), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n458), .B1(new_n423), .B2(new_n432), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n400), .A2(new_n423), .A3(new_n425), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n328), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n379), .A2(new_n381), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n372), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n543), .A2(new_n478), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT81), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n543), .A2(new_n544), .A3(new_n478), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n539), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n543), .B(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n480), .A2(new_n481), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .A4(new_n539), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n533), .A2(new_n538), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n578), .A2(new_n580), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G169), .ZN(new_n652));
  INV_X1    g0452(.A(new_n584), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n652), .A2(new_n653), .B1(new_n625), .B2(new_n569), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n607), .A2(new_n603), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n605), .A3(new_n604), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n626), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n650), .B1(new_n547), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n638), .B1(new_n467), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT89), .ZN(G369));
  NAND2_X1  g0463(.A1(new_n259), .A2(new_n217), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(G343), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n654), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n565), .B2(new_n570), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n585), .A2(new_n677), .A3(new_n626), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n609), .A2(new_n674), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n654), .B2(new_n673), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n609), .B(new_n617), .C1(new_n610), .C2(new_n673), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n658), .A2(new_n603), .A3(new_n674), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n517), .A2(G116), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT92), .Z(new_n690));
  INV_X1    g0490(.A(new_n220), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(G1), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n694), .A2(new_n695), .B1(new_n216), .B2(new_n693), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT28), .Z(new_n698));
  INV_X1    g0498(.A(new_n647), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n699), .A2(new_n501), .B1(new_n640), .B2(new_n641), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n585), .A2(new_n609), .A3(new_n617), .A4(new_n626), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n539), .A4(new_n673), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n576), .A2(new_n299), .B1(new_n586), .B2(G264), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n499), .A2(new_n510), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n587), .A2(G179), .A3(new_n592), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n510), .A2(new_n704), .ZN(new_n708));
  INV_X1    g0508(.A(new_n706), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT30), .A4(new_n499), .ZN(new_n710));
  INV_X1    g0510(.A(new_n499), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n510), .A2(G179), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n582), .A4(new_n593), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT31), .B1(new_n714), .B2(new_n674), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n702), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n673), .B1(new_n649), .B2(new_n660), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n647), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n539), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT26), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(KEYINPUT26), .B2(new_n642), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT29), .B(new_n673), .C1(new_n732), .C2(new_n660), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n723), .A2(new_n725), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n722), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n698), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n258), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n247), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n692), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n686), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n684), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n270), .A2(G355), .A3(new_n220), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n242), .A2(new_n504), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n691), .A2(new_n270), .ZN(new_n747));
  INV_X1    g0547(.A(new_n303), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n216), .B2(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n745), .B1(G116), .B2(new_n220), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n218), .B1(G20), .B2(new_n337), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n692), .B(new_n741), .C1(new_n750), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n757));
  INV_X1    g0557(.A(new_n754), .ZN(new_n758));
  INV_X1    g0558(.A(new_n270), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n217), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n301), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G107), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT32), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n759), .B(new_n768), .C1(G87), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n217), .A2(new_n583), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n301), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n774), .A2(G68), .B1(new_n775), .B2(G50), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n765), .A2(KEYINPUT32), .A3(new_n766), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n301), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n217), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(G97), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n772), .A2(G190), .A3(new_n424), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n772), .A2(new_n764), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n254), .B1(new_n783), .B2(new_n352), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT96), .Z(new_n785));
  NAND4_X1  g0585(.A1(new_n771), .A2(new_n776), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n782), .ZN(new_n787));
  INV_X1    g0587(.A(new_n765), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(G322), .B1(new_n788), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(new_n783), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n270), .B1(new_n790), .B2(G311), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n775), .A2(G326), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n774), .A2(new_n794), .B1(new_n770), .B2(G303), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n780), .A2(G294), .B1(new_n762), .B2(G283), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n792), .A2(new_n793), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n758), .B1(new_n786), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n757), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n753), .B(KEYINPUT97), .Z(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n800), .C1(new_n684), .C2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n744), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  AOI21_X1  g0604(.A(new_n673), .B1(new_n441), .B2(new_n442), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n457), .B1(new_n464), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n443), .A2(new_n456), .A3(new_n673), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n723), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n443), .A2(new_n674), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n441), .A2(new_n442), .A3(new_n460), .A4(new_n459), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n810), .B1(new_n457), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n673), .B(new_n814), .C1(new_n649), .C2(new_n660), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n722), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n742), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n722), .A2(new_n809), .A3(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n758), .A2(new_n752), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n742), .B1(new_n820), .B2(G77), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n787), .A2(G143), .B1(new_n790), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(new_n775), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(new_n774), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n366), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT34), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n761), .A2(new_n238), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n270), .B1(new_n765), .B2(new_n830), .C1(new_n779), .C2(new_n254), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(G50), .C2(new_n770), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n826), .A2(new_n827), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n779), .A2(new_n516), .B1(new_n782), .B2(new_n575), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT98), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n823), .A2(new_n590), .B1(new_n761), .B2(new_n515), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n825), .A2(new_n838), .B1(new_n769), .B2(new_n445), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n759), .B1(new_n765), .B2(new_n840), .C1(new_n594), .C2(new_n783), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n837), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n833), .A2(new_n834), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n821), .B1(new_n843), .B2(new_n754), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n814), .B2(new_n752), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n819), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n475), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n218), .A2(new_n217), .A3(new_n594), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n848), .B2(KEYINPUT35), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT36), .ZN(new_n855));
  OR3_X1    g0655(.A1(new_n275), .A2(new_n216), .A3(new_n352), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n247), .B(G13), .C1(new_n856), .C2(new_n237), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n631), .B(KEYINPUT18), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n667), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n807), .B(KEYINPUT100), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n815), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n423), .B(new_n674), .C1(new_n432), .C2(new_n426), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n431), .A2(new_n429), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n430), .B1(new_n399), .B2(G169), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n423), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n423), .A2(new_n674), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n634), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT16), .B1(new_n287), .B2(new_n280), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n323), .B1(new_n334), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n668), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n319), .A2(new_n327), .B1(new_n345), .B2(KEYINPUT18), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n348), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n335), .A2(new_n668), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n877), .A2(new_n878), .A3(new_n324), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n630), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n874), .A2(new_n880), .A3(new_n324), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n879), .A2(new_n345), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n871), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n874), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n349), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n345), .A2(new_n877), .A3(new_n878), .A4(new_n324), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n860), .B1(new_n870), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT101), .B(new_n860), .C1(new_n870), .C2(new_n890), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n336), .A2(new_n338), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n324), .B1(new_n290), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n290), .A2(new_n667), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT102), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n631), .A2(new_n877), .A3(new_n324), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n887), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n328), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n898), .B1(new_n859), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n876), .A2(new_n882), .A3(new_n871), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n895), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n432), .A2(new_n423), .A3(new_n673), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n883), .A2(new_n889), .A3(KEYINPUT39), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n893), .A2(new_n894), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n736), .A2(new_n466), .A3(new_n733), .A4(new_n726), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n638), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n808), .B1(new_n863), .B2(new_n868), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n719), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n883), .A2(new_n889), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n902), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT102), .B1(new_n902), .B2(KEYINPUT37), .ZN(new_n924));
  INV_X1    g0724(.A(new_n887), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n877), .B1(new_n632), .B2(new_n328), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n871), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n919), .B1(new_n928), .B2(new_n889), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n466), .A3(new_n719), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n918), .A2(new_n719), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n907), .B2(new_n908), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(KEYINPUT40), .B1(new_n921), .B2(new_n920), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n467), .B2(new_n720), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(new_n936), .A3(G330), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n917), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n247), .B2(new_n739), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n917), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n858), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NAND2_X1  g0741(.A1(new_n226), .A2(new_n747), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n755), .C1(new_n220), .C2(new_n435), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n742), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT105), .Z(new_n945));
  OAI22_X1  g0745(.A1(new_n825), .A2(new_n766), .B1(new_n769), .B2(new_n254), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(G68), .B2(new_n780), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n782), .A2(new_n366), .B1(new_n765), .B2(new_n824), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n759), .B(new_n948), .C1(G50), .C2(new_n790), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n775), .A2(G143), .B1(new_n762), .B2(G77), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n769), .A2(new_n594), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G107), .A2(new_n780), .B1(new_n775), .B2(G311), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n270), .B1(new_n787), .B2(G303), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G283), .A2(new_n790), .B1(new_n788), .B2(G317), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n774), .A2(G294), .B1(new_n762), .B2(G97), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n951), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n754), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n528), .A2(new_n673), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n533), .A3(new_n538), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n730), .B2(new_n964), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n945), .B1(new_n962), .B2(new_n963), .C1(new_n966), .C2(new_n801), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n679), .B(new_n680), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n686), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n737), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n700), .B1(new_n699), .B2(new_n673), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n645), .A2(new_n647), .A3(new_n674), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n681), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT103), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT103), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n681), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n681), .A2(new_n973), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT44), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n687), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT104), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n970), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(KEYINPUT104), .A3(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n737), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n692), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n741), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n973), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n995), .A2(new_n585), .B1(new_n545), .B2(new_n546), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n679), .A2(new_n973), .A3(new_n680), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(new_n673), .B1(KEYINPUT42), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(KEYINPUT42), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n986), .A2(new_n973), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n967), .B1(new_n994), .B2(new_n1005), .ZN(G387));
  NAND2_X1  g0806(.A1(new_n970), .A2(new_n692), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT111), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(KEYINPUT111), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n969), .A2(new_n737), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n679), .A2(new_n801), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n747), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1016));
  OR3_X1    g0816(.A1(new_n1016), .A2(G50), .A3(new_n251), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(G50), .B2(new_n251), .ZN(new_n1018));
  AOI21_X1  g0818(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1019));
  AND4_X1   g0819(.A1(new_n690), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1015), .B(new_n1020), .C1(new_n231), .C2(new_n748), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n270), .A2(new_n220), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n690), .A2(new_n1022), .B1(G107), .B2(new_n220), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT107), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n755), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n742), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n783), .A2(new_n238), .B1(new_n765), .B2(new_n366), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n759), .B(new_n1027), .C1(G50), .C2(new_n787), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n435), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n780), .A2(new_n1029), .B1(new_n762), .B2(G97), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n775), .A2(G159), .B1(new_n770), .B2(G77), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n256), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n774), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n270), .B1(new_n788), .B2(G326), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n779), .A2(new_n838), .B1(new_n769), .B2(new_n575), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n787), .A2(G317), .B1(new_n790), .B2(G303), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT109), .B(G322), .Z(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n823), .B2(new_n1038), .C1(new_n840), .C2(new_n825), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1035), .B1(new_n594), .B2(new_n761), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT110), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n758), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1026), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n969), .A2(new_n741), .B1(new_n1014), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1013), .A2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n995), .A2(new_n753), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G317), .A2(new_n775), .B1(new_n787), .B2(G311), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n759), .B1(new_n783), .B2(new_n575), .C1(new_n765), .C2(new_n1038), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n763), .B1(new_n825), .B2(new_n590), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n779), .A2(new_n594), .B1(new_n769), .B2(new_n838), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT115), .Z(new_n1060));
  INV_X1    g0860(.A(G143), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n769), .A2(new_n238), .B1(new_n765), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT113), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n270), .B1(new_n515), .B2(new_n761), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT114), .Z(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n775), .B1(new_n787), .B2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n779), .A2(new_n352), .B1(new_n783), .B2(new_n251), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G50), .B2(new_n774), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n754), .B1(new_n1060), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n755), .B1(new_n516), .B2(new_n220), .C1(new_n235), .C2(new_n1015), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1053), .A2(new_n742), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n984), .B(new_n986), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n740), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n970), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n693), .B1(new_n988), .B2(new_n989), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(G390));
  NAND3_X1  g0881(.A1(new_n918), .A2(new_n719), .A3(G330), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n909), .A2(new_n912), .B1(new_n870), .B2(new_n910), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n910), .B1(new_n907), .B2(new_n908), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n869), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n673), .B(new_n814), .C1(new_n732), .C2(new_n660), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n861), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n861), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n869), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n928), .A2(new_n889), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n1093), .A3(new_n910), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n883), .A2(new_n889), .A3(KEYINPUT39), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1093), .B2(new_n895), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n911), .B1(new_n862), .B2(new_n869), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1082), .B(new_n1094), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n740), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1096), .A2(new_n752), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n742), .B1(new_n1032), .B2(new_n820), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n782), .A2(new_n830), .B1(new_n765), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n759), .B(new_n1104), .C1(new_n790), .C2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n769), .A2(new_n366), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G159), .A2(new_n780), .B1(new_n774), .B2(G137), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n775), .A2(G128), .B1(new_n762), .B2(G50), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n759), .B1(new_n769), .B2(new_n515), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT116), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n783), .A2(new_n516), .B1(new_n765), .B2(new_n575), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G116), .B2(new_n787), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n774), .A2(G107), .B1(new_n775), .B2(G283), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n829), .B1(G77), .B2(new_n780), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1112), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1102), .B1(new_n1120), .B2(new_n754), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1100), .B1(new_n1101), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n722), .A2(new_n466), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n915), .A2(new_n638), .A3(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n547), .A2(new_n627), .A3(new_n674), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n714), .A2(new_n674), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT31), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n715), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n814), .B(G330), .C1(new_n1125), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1086), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n1082), .B1(new_n815), .B2(new_n861), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1091), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1131), .A2(new_n1082), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1099), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1090), .A3(new_n1098), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n692), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1122), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(KEYINPUT122), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT57), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n370), .A2(new_n667), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n382), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n382), .B1(new_n370), .B2(new_n667), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n935), .A2(new_n1153), .A3(new_n721), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n931), .B2(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n914), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n931), .A2(G330), .A3(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1153), .B1(new_n935), .B2(new_n721), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1096), .A2(new_n911), .B1(new_n891), .B2(new_n892), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n894), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT119), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1124), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n915), .A2(KEYINPUT119), .A3(new_n638), .A4(new_n1123), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1139), .A2(new_n1166), .A3(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT120), .B1(new_n1139), .B2(new_n1166), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1143), .B(new_n1144), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT120), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1136), .A2(new_n1090), .A3(new_n1098), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1167), .A3(new_n1162), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1143), .B1(new_n1176), .B2(new_n1144), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(KEYINPUT57), .A3(new_n1167), .A4(new_n1162), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n692), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1171), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1162), .A2(new_n741), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n742), .B1(new_n820), .B2(G50), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n759), .A2(new_n304), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n770), .B2(G77), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT117), .Z(new_n1185));
  AOI22_X1  g0985(.A1(new_n780), .A2(G68), .B1(new_n762), .B2(G58), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n516), .B2(new_n825), .C1(new_n594), .C2(new_n823), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n787), .A2(G107), .B1(new_n788), .B2(G283), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n435), .B2(new_n783), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT58), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1183), .B(new_n236), .C1(G33), .C2(G41), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1103), .A2(new_n823), .B1(new_n825), .B2(new_n830), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n787), .A2(G128), .B1(new_n790), .B2(G137), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n769), .B2(new_n1105), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G150), .C2(new_n780), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n762), .A2(G159), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1193), .B1(KEYINPUT58), .B2(new_n1190), .C1(new_n1199), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1182), .B1(new_n1204), .B2(new_n754), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1155), .B2(new_n752), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT118), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1142), .B1(new_n1180), .B2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1178), .A2(new_n692), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1144), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT121), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1212), .A3(new_n1170), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1208), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(KEYINPUT122), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1209), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(G375));
  OAI21_X1  g1017(.A(new_n742), .B1(new_n820), .B2(G68), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n779), .A2(new_n236), .B1(new_n769), .B2(new_n766), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n775), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n759), .B1(new_n788), .B2(G128), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n787), .A2(G137), .B1(new_n790), .B2(G150), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n774), .A2(new_n1106), .B1(new_n762), .B2(G58), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n775), .A2(G294), .B1(new_n790), .B2(G107), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n594), .B2(new_n825), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT123), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n759), .B1(new_n765), .B2(new_n590), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G283), .B2(new_n787), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n780), .A2(new_n1029), .B1(new_n762), .B2(G77), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n516), .C2(new_n769), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1218), .B1(new_n1232), .B2(new_n754), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n869), .B2(new_n752), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1135), .B2(new_n740), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT124), .Z(new_n1236));
  NAND2_X1  g1036(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1137), .A2(new_n993), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(G381));
  NAND4_X1  g1039(.A1(new_n1080), .A2(new_n846), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1013), .A2(new_n803), .A3(new_n1051), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1240), .A2(G387), .A3(G378), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(new_n1242), .ZN(G407));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n670), .A2(new_n671), .A3(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1216), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(G213), .A3(G407), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT125), .ZN(G409));
  NAND2_X1  g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1241), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(G387), .A2(KEYINPUT126), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(G387), .B2(new_n1251), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(new_n1080), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1213), .A2(G378), .A3(new_n1214), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1181), .B(new_n1206), .C1(new_n1176), .C2(new_n992), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1244), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1246), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1237), .B1(new_n1136), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1124), .A2(new_n1135), .A3(KEYINPUT60), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n692), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1236), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n846), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1264), .A2(new_n846), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1246), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1268), .B(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1258), .A2(new_n1268), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1254), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1253), .B(G390), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1258), .A2(new_n1268), .A3(KEYINPUT63), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1272), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(G405));
  NAND3_X1  g1083(.A1(new_n1209), .A2(new_n1244), .A3(new_n1215), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1255), .A2(KEYINPUT127), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1268), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1209), .A2(new_n1289), .A3(new_n1244), .A4(new_n1215), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1254), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1213), .A2(KEYINPUT122), .A3(new_n1214), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT122), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1294), .A2(new_n1295), .A3(G378), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1290), .B1(new_n1296), .B2(new_n1285), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1268), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1278), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1293), .A2(new_n1300), .ZN(G402));
endmodule


