

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578;

  XNOR2_X2 U319 ( .A(n293), .B(KEYINPUT83), .ZN(n432) );
  XNOR2_X2 U320 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n293) );
  XOR2_X1 U321 ( .A(n304), .B(n421), .Z(n526) );
  XNOR2_X2 U322 ( .A(n450), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n410) );
  XNOR2_X1 U324 ( .A(n392), .B(n287), .ZN(n356) );
  XNOR2_X1 U325 ( .A(n343), .B(n342), .ZN(n564) );
  AND2_X1 U326 ( .A1(G232GAT), .A2(G233GAT), .ZN(n287) );
  INV_X1 U327 ( .A(n392), .ZN(n393) );
  XNOR2_X1 U328 ( .A(n394), .B(n393), .ZN(n395) );
  NOR2_X1 U329 ( .A1(n463), .A2(n562), .ZN(n448) );
  XNOR2_X1 U330 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U331 ( .A(n357), .B(n356), .ZN(n363) );
  XNOR2_X1 U332 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U333 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G176GAT), .B(KEYINPUT85), .Z(n289) );
  XNOR2_X1 U335 ( .A(KEYINPUT20), .B(KEYINPUT67), .ZN(n288) );
  XNOR2_X1 U336 ( .A(n289), .B(n288), .ZN(n300) );
  XOR2_X1 U337 ( .A(G190GAT), .B(G134GAT), .Z(n291) );
  XOR2_X1 U338 ( .A(G15GAT), .B(G127GAT), .Z(n372) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n391) );
  XNOR2_X1 U340 ( .A(n372), .B(n391), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U342 ( .A(n292), .B(G99GAT), .Z(n298) );
  XOR2_X1 U343 ( .A(KEYINPUT84), .B(n432), .Z(n295) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(n296), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U349 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n302) );
  XNOR2_X1 U350 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(G169GAT), .B(n303), .Z(n421) );
  XOR2_X1 U353 ( .A(KEYINPUT88), .B(G155GAT), .Z(n306) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U356 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n307) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n446) );
  XOR2_X1 U358 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n310) );
  XNOR2_X1 U359 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n322) );
  XOR2_X1 U361 ( .A(G106GAT), .B(G218GAT), .Z(n312) );
  XOR2_X1 U362 ( .A(G50GAT), .B(G162GAT), .Z(n351) );
  XOR2_X1 U363 ( .A(G148GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U364 ( .A(n351), .B(n390), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(n313), .B(KEYINPUT23), .Z(n320) );
  XOR2_X1 U367 ( .A(G204GAT), .B(G211GAT), .Z(n315) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n412) );
  XOR2_X1 U370 ( .A(n412), .B(KEYINPUT90), .Z(n317) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U373 ( .A(G22GAT), .B(n318), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U375 ( .A(n322), .B(n321), .Z(n323) );
  XOR2_X1 U376 ( .A(n446), .B(n323), .Z(n463) );
  XOR2_X1 U377 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n325) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT71), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n343) );
  XOR2_X1 U380 ( .A(G141GAT), .B(G15GAT), .Z(n327) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G113GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G36GAT), .Z(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n339) );
  XOR2_X1 U385 ( .A(G29GAT), .B(G43GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n361) );
  XOR2_X1 U388 ( .A(G8GAT), .B(KEYINPUT74), .Z(n333) );
  XNOR2_X1 U389 ( .A(G22GAT), .B(G1GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n371) );
  XNOR2_X1 U391 ( .A(n361), .B(n371), .ZN(n337) );
  XOR2_X1 U392 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n335) );
  XNOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT75), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n341) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U399 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n345) );
  XNOR2_X1 U400 ( .A(KEYINPUT11), .B(KEYINPUT66), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n354) );
  XOR2_X1 U402 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n350) );
  INV_X1 U403 ( .A(KEYINPUT79), .ZN(n346) );
  NAND2_X1 U404 ( .A1(n346), .A2(G134GAT), .ZN(n349) );
  INV_X1 U405 ( .A(G134GAT), .ZN(n347) );
  NAND2_X1 U406 ( .A1(n347), .A2(KEYINPUT79), .ZN(n348) );
  NAND2_X1 U407 ( .A1(n349), .A2(n348), .ZN(n438) );
  XNOR2_X1 U408 ( .A(n350), .B(n438), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(n354), .B(n353), .Z(n357) );
  XNOR2_X1 U411 ( .A(G99GAT), .B(G106GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n355), .B(G85GAT), .ZN(n392) );
  XOR2_X1 U413 ( .A(G92GAT), .B(KEYINPUT80), .Z(n359) );
  XNOR2_X1 U414 ( .A(G190GAT), .B(G218GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U416 ( .A(G36GAT), .B(n360), .Z(n420) );
  XNOR2_X1 U417 ( .A(n361), .B(n420), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n556) );
  INV_X1 U419 ( .A(KEYINPUT81), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n556), .B(n364), .ZN(n541) );
  XNOR2_X1 U421 ( .A(n541), .B(KEYINPUT36), .ZN(n485) );
  XOR2_X1 U422 ( .A(G64GAT), .B(G78GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G155GAT), .B(G211GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U425 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n368) );
  XNOR2_X1 U426 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n379) );
  XOR2_X1 U429 ( .A(n372), .B(n371), .Z(n374) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U432 ( .A(G57GAT), .B(KEYINPUT13), .Z(n387) );
  XOR2_X1 U433 ( .A(n375), .B(n387), .Z(n377) );
  XNOR2_X1 U434 ( .A(G183GAT), .B(G71GAT), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n573) );
  NAND2_X1 U437 ( .A1(n485), .A2(n573), .ZN(n381) );
  XOR2_X1 U438 ( .A(KEYINPUT69), .B(KEYINPUT45), .Z(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n399) );
  XOR2_X1 U440 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n383) );
  XNOR2_X1 U441 ( .A(G204GAT), .B(G92GAT), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n398) );
  XOR2_X1 U443 ( .A(KEYINPUT33), .B(KEYINPUT77), .Z(n385) );
  NAND2_X1 U444 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n386), .B(KEYINPUT32), .Z(n389) );
  XOR2_X1 U447 ( .A(G176GAT), .B(G64GAT), .Z(n413) );
  XNOR2_X1 U448 ( .A(n387), .B(n413), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n394) );
  XOR2_X1 U451 ( .A(n398), .B(n397), .Z(n569) );
  NOR2_X1 U452 ( .A1(n399), .A2(n569), .ZN(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT112), .B(n400), .Z(n401) );
  NOR2_X1 U454 ( .A1(n564), .A2(n401), .ZN(n402) );
  XNOR2_X1 U455 ( .A(KEYINPUT113), .B(n402), .ZN(n409) );
  XNOR2_X1 U456 ( .A(n569), .B(KEYINPUT65), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT41), .ZN(n551) );
  NAND2_X1 U458 ( .A1(n551), .A2(n564), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(KEYINPUT46), .ZN(n405) );
  INV_X1 U460 ( .A(n573), .ZN(n470) );
  NAND2_X1 U461 ( .A1(n405), .A2(n470), .ZN(n406) );
  NOR2_X1 U462 ( .A1(n556), .A2(n406), .ZN(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT47), .B(n407), .ZN(n408) );
  AND2_X1 U464 ( .A1(n409), .A2(n408), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n529) );
  XOR2_X1 U466 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U469 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n417) );
  XNOR2_X1 U470 ( .A(G8GAT), .B(KEYINPUT96), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U472 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U474 ( .A(n423), .B(n422), .Z(n518) );
  XOR2_X1 U475 ( .A(n518), .B(KEYINPUT121), .Z(n424) );
  NOR2_X1 U476 ( .A1(n529), .A2(n424), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n425), .B(KEYINPUT54), .ZN(n447) );
  XOR2_X1 U478 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(G57GAT), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U481 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n429) );
  XNOR2_X1 U482 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U484 ( .A(n431), .B(n430), .Z(n444) );
  XOR2_X1 U485 ( .A(n432), .B(KEYINPUT92), .Z(n434) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n442) );
  XOR2_X1 U488 ( .A(G148GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(G127GAT), .B(G120GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n437), .B(G85GAT), .Z(n440) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n525) );
  NAND2_X1 U497 ( .A1(n447), .A2(n525), .ZN(n562) );
  XNOR2_X1 U498 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  NOR2_X1 U499 ( .A1(n526), .A2(n449), .ZN(n450) );
  NAND2_X1 U500 ( .A1(n560), .A2(n541), .ZN(n452) );
  NAND2_X1 U501 ( .A1(n551), .A2(n560), .ZN(n456) );
  XOR2_X1 U502 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n454) );
  XOR2_X1 U503 ( .A(G176GAT), .B(KEYINPUT56), .Z(n453) );
  XNOR2_X1 U504 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U505 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  INV_X1 U506 ( .A(n564), .ZN(n504) );
  NOR2_X1 U507 ( .A1(n504), .A2(n569), .ZN(n490) );
  XNOR2_X1 U508 ( .A(n518), .B(KEYINPUT27), .ZN(n460) );
  XNOR2_X1 U509 ( .A(n463), .B(KEYINPUT28), .ZN(n481) );
  NOR2_X1 U510 ( .A1(n460), .A2(n481), .ZN(n527) );
  NAND2_X1 U511 ( .A1(n526), .A2(n527), .ZN(n457) );
  INV_X1 U512 ( .A(n525), .ZN(n545) );
  NAND2_X1 U513 ( .A1(n457), .A2(n545), .ZN(n469) );
  XOR2_X1 U514 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n459) );
  NAND2_X1 U515 ( .A1(n463), .A2(n526), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n563) );
  NOR2_X1 U517 ( .A1(n563), .A2(n460), .ZN(n544) );
  OR2_X1 U518 ( .A1(n526), .A2(n518), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(n461), .Z(n462) );
  NOR2_X1 U520 ( .A1(n463), .A2(n462), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n465), .B(n464), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n544), .A2(n466), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n467), .A2(n525), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n486) );
  NOR2_X1 U526 ( .A1(n541), .A2(n470), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U528 ( .A1(n486), .A2(n472), .ZN(n505) );
  NAND2_X1 U529 ( .A1(n490), .A2(n505), .ZN(n482) );
  NOR2_X1 U530 ( .A1(n525), .A2(n482), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U534 ( .A1(n518), .A2(n482), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n526), .A2(n482), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  INV_X1 U541 ( .A(n481), .ZN(n522) );
  NOR2_X1 U542 ( .A1(n522), .A2(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n573), .A2(n486), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n485), .A2(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT104), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n489), .ZN(n514) );
  NAND2_X1 U549 ( .A1(n490), .A2(n514), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n491), .ZN(n500) );
  NOR2_X1 U551 ( .A1(n500), .A2(n525), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U554 ( .A1(n500), .A2(n518), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n497) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n500), .A2(n526), .ZN(n498) );
  XOR2_X1 U561 ( .A(n499), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U562 ( .A1(n522), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n507) );
  AND2_X1 U567 ( .A1(n504), .A2(n551), .ZN(n515) );
  NAND2_X1 U568 ( .A1(n515), .A2(n505), .ZN(n510) );
  NOR2_X1 U569 ( .A1(n525), .A2(n510), .ZN(n506) );
  XOR2_X1 U570 ( .A(n507), .B(n506), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n518), .A2(n510), .ZN(n508) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n526), .A2(n510), .ZN(n509) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n521) );
  NOR2_X1 U580 ( .A1(n525), .A2(n521), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n521), .ZN(n519) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n526), .A2(n521), .ZN(n520) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n520), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT115), .Z(n533) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n528) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n531), .B(KEYINPUT114), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n540), .A2(n564), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U598 ( .A1(n551), .A2(n540), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT116), .Z(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n540), .A2(n573), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U609 ( .A1(n529), .A2(n546), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n557), .A2(n564), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n549) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(n550), .Z(n553) );
  NAND2_X1 U616 ( .A1(n557), .A2(n551), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n557), .A2(n573), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT120), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n560), .A2(n564), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n573), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n576) );
  NAND2_X1 U628 ( .A1(n564), .A2(n576), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U634 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U637 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n574), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NAND2_X1 U640 ( .A1(n485), .A2(n576), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

