//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT3), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n462), .A2(new_n463), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND3_X1  g055(.A1(new_n464), .A2(G2105), .A3(new_n467), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n465), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n468), .A2(G136), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n483), .A2(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(new_n467), .A3(new_n471), .A4(new_n465), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(G138), .A3(new_n465), .A4(new_n467), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n464), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT69), .B(G114), .ZN(new_n497));
  OAI211_X1 g072(.A(G2104), .B(new_n496), .C1(new_n497), .C2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT71), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(new_n509), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n504), .A2(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(G88), .B1(new_n513), .B2(G50), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n512), .A2(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n504), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n519), .B(new_n521), .C1(new_n525), .C2(KEYINPUT72), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n511), .A2(new_n529), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n516), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n516), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n513), .A2(G43), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n504), .A2(G81), .A3(new_n510), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT73), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n536), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n513), .A2(G53), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n512), .A2(G91), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n516), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n556), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  XNOR2_X1  g137(.A(G166), .B(new_n562), .ZN(G303));
  NAND2_X1  g138(.A1(new_n512), .A2(G87), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT76), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n510), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(G49), .A2(new_n513), .B1(new_n566), .B2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n510), .A2(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT77), .Z(new_n571));
  AOI21_X1  g146(.A(new_n516), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT78), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n512), .A2(G86), .B1(new_n513), .B2(G48), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G305));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n511), .A2(new_n576), .B1(new_n523), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n580), .A2(new_n581), .B1(new_n516), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n512), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  NAND2_X1  g161(.A1(new_n510), .A2(G66), .ZN(new_n587));
  INV_X1    g162(.A(G79), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n505), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n513), .B2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  OR3_X1    g170(.A1(G168), .A2(KEYINPUT80), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(G168), .B2(new_n595), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n556), .A2(new_n558), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(G868), .C2(new_n598), .ZN(G297));
  OAI211_X1 g174(.A(new_n596), .B(new_n597), .C1(G868), .C2(new_n598), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n544), .A2(new_n595), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n591), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n595), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g182(.A1(new_n476), .A2(G2105), .A3(new_n472), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G2100), .ZN(new_n612));
  INV_X1    g187(.A(G2100), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(KEYINPUT82), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n482), .A2(G123), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n468), .A2(G135), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n465), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n610), .A2(new_n611), .A3(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n619), .A2(G2096), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n614), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT83), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n628), .B(new_n634), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(G14), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n636), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(KEYINPUT18), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n653), .A2(new_n658), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n658), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n661));
  AOI211_X1 g236(.A(new_n657), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n660), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  XOR2_X1   g239(.A(G1991), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1981), .B(G1986), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(new_n670), .ZN(G229));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G20), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT23), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G299), .B2(G16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1956), .ZN(new_n676));
  INV_X1    g251(.A(G2090), .ZN(new_n677));
  NAND2_X1  g252(.A1(G162), .A2(G29), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G29), .B2(G35), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n676), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT95), .Z(new_n684));
  INV_X1    g259(.A(G34), .ZN(new_n685));
  AOI21_X1  g260(.A(G29), .B1(new_n685), .B2(KEYINPUT24), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(KEYINPUT24), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n479), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT91), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(G27), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G164), .B2(new_n688), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G2078), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n468), .A2(G139), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(G115), .A2(G2104), .ZN(new_n703));
  INV_X1    g278(.A(G127), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n472), .B2(new_n704), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n701), .A2(new_n702), .B1(G2105), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G29), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G29), .B2(G33), .ZN(new_n709));
  INV_X1    g284(.A(G2072), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n695), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n482), .A2(G129), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n468), .A2(G141), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n477), .A2(G105), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n712), .A2(new_n713), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G32), .B(new_n717), .S(G29), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT27), .B(G1996), .Z(new_n719));
  AOI211_X1 g294(.A(new_n692), .B(new_n711), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n672), .A2(G21), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G168), .B2(new_n672), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1966), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n710), .B2(new_n709), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n720), .B(new_n724), .C1(G2090), .C2(new_n681), .ZN(new_n725));
  NOR2_X1   g300(.A1(G171), .A2(new_n672), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G5), .B2(new_n672), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT93), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n672), .A2(G19), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n545), .B2(new_n672), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G1341), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n688), .A2(G26), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT28), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n482), .A2(G128), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n465), .A2(G116), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n468), .A2(G140), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2067), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n730), .A2(new_n733), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G4), .A2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n592), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(G1348), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n727), .A2(new_n728), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G11), .ZN(new_n750));
  INV_X1    g325(.A(G28), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT30), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n689), .B2(new_n690), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n749), .B(new_n757), .C1(new_n688), .C2(new_n619), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n694), .A2(G2078), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n718), .A2(new_n719), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n748), .B(new_n761), .C1(G1341), .C2(new_n732), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n684), .A2(new_n725), .A3(new_n744), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n672), .A2(G23), .ZN(new_n764));
  INV_X1    g339(.A(G288), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n672), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT33), .B(G1976), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n672), .A2(G22), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G166), .B2(new_n672), .ZN(new_n770));
  INV_X1    g345(.A(G1971), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G6), .B(G305), .S(G16), .Z(new_n773));
  XOR2_X1   g348(.A(KEYINPUT32), .B(G1981), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n768), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT34), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(KEYINPUT34), .ZN(new_n778));
  MUX2_X1   g353(.A(G24), .B(G290), .S(G16), .Z(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1986), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n688), .A2(G25), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n482), .A2(G119), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n468), .A2(G131), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n465), .A2(G107), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT87), .Z(new_n787));
  OAI21_X1  g362(.A(new_n781), .B1(new_n787), .B2(new_n688), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT35), .B(G1991), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  NAND4_X1  g365(.A1(new_n777), .A2(new_n778), .A3(new_n780), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT36), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n763), .A2(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  INV_X1    g369(.A(G93), .ZN(new_n795));
  INV_X1    g370(.A(G55), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n511), .A2(new_n795), .B1(new_n523), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n516), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G860), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n591), .A2(new_n601), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n544), .A2(KEYINPUT96), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(new_n536), .C1(new_n539), .C2(new_n543), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n800), .B1(new_n807), .B2(new_n809), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n806), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n801), .B1(new_n816), .B2(KEYINPUT39), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n804), .B1(new_n817), .B2(new_n818), .ZN(G145));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n707), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n717), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n741), .ZN(new_n823));
  INV_X1    g398(.A(new_n499), .ZN(new_n824));
  AOI211_X1 g399(.A(KEYINPUT98), .B(new_n492), .C1(new_n493), .C2(KEYINPUT4), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n491), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(KEYINPUT99), .B(new_n824), .C1(new_n825), .C2(new_n828), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n823), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n468), .A2(G142), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n465), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G130), .B2(new_n482), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n609), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n787), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n834), .A2(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n846));
  OR3_X1    g421(.A1(new_n834), .A2(KEYINPUT101), .A3(new_n841), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n843), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n619), .B(G160), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n834), .B2(new_n841), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g430(.A(G288), .B(G305), .Z(new_n856));
  XNOR2_X1  g431(.A(G290), .B(G166), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT103), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n865), .B2(KEYINPUT42), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  NOR2_X1   g443(.A1(G299), .A2(new_n591), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n592), .A2(new_n598), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n814), .A2(new_n604), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n813), .B1(G559), .B2(new_n591), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n869), .B2(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(G299), .A2(new_n591), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n592), .A2(new_n598), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT41), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n872), .A3(new_n873), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n868), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n875), .A2(new_n868), .A3(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n867), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n883), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n866), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(G868), .B2(new_n800), .ZN(G295));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  XNOR2_X1  g466(.A(G295), .B(new_n891), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n894));
  INV_X1    g469(.A(new_n812), .ZN(new_n895));
  AOI21_X1  g470(.A(G301), .B1(new_n895), .B2(new_n810), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n811), .A2(new_n812), .A3(G171), .ZN(new_n897));
  OAI21_X1  g472(.A(G286), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(G171), .B1(new_n811), .B2(new_n812), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(G301), .A3(new_n810), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n900), .A3(G168), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n871), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n881), .B1(new_n898), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n865), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n863), .A2(new_n864), .ZN(new_n908));
  INV_X1    g483(.A(new_n881), .ZN(new_n909));
  INV_X1    g484(.A(new_n901), .ZN(new_n910));
  AOI21_X1  g485(.A(G168), .B1(new_n899), .B2(new_n900), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n902), .ZN(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n893), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT106), .B1(new_n912), .B2(new_n902), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n919), .B(new_n908), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n863), .A2(new_n919), .A3(new_n864), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n905), .A2(new_n906), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n918), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n907), .A2(new_n914), .A3(new_n893), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n907), .A2(new_n914), .A3(new_n931), .A4(new_n893), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n927), .B1(new_n936), .B2(new_n937), .ZN(G397));
  XOR2_X1   g513(.A(KEYINPUT111), .B(G1384), .Z(new_n939));
  AOI21_X1  g514(.A(KEYINPUT45), .B1(new_n833), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n469), .A2(new_n478), .A3(G40), .A4(new_n475), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n741), .A2(G2067), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n736), .A2(new_n949), .A3(new_n740), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n951), .A2(new_n717), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n946), .A2(new_n947), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n947), .B2(new_n946), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT47), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n944), .A2(new_n951), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT114), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n717), .B(new_n945), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n943), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n787), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n959), .A2(new_n789), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n943), .B1(new_n961), .B2(new_n950), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n787), .B(new_n789), .Z(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n944), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(G290), .A2(G1986), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n943), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT48), .Z(new_n967));
  AOI211_X1 g542(.A(new_n955), .B(new_n962), .C1(new_n964), .C2(new_n967), .ZN(new_n968));
  AOI22_X1  g543(.A1(G303), .A2(G8), .B1(KEYINPUT116), .B2(KEYINPUT55), .ZN(new_n969));
  NOR2_X1   g544(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n969), .B(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT118), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n829), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n494), .B2(new_n499), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n942), .B1(KEYINPUT50), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n973), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n677), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n976), .A2(new_n978), .A3(new_n973), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n941), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n831), .A2(KEYINPUT45), .A3(new_n832), .A4(new_n939), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n985), .A2(KEYINPUT115), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(KEYINPUT115), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n982), .B1(new_n988), .B2(new_n771), .ZN(new_n989));
  OAI21_X1  g564(.A(G8), .B1(new_n989), .B2(KEYINPUT119), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n991), .B(new_n982), .C1(new_n988), .C2(new_n771), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n972), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1981), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n573), .A2(new_n994), .A3(new_n574), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n573), .B2(new_n574), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT117), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n829), .A2(new_n975), .A3(new_n942), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1005), .B2(G288), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n765), .A2(G1976), .ZN(new_n1007));
  OR3_X1    g582(.A1(new_n1006), .A2(KEYINPUT52), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n988), .A2(new_n771), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n829), .A2(new_n974), .A3(new_n975), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n941), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n677), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1002), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1016), .B2(new_n971), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n993), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n985), .B(KEYINPUT115), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n984), .A3(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n598), .B(KEYINPUT57), .ZN(new_n1022));
  INV_X1    g597(.A(G1956), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n976), .B2(new_n978), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1021), .A2(KEYINPUT125), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(KEYINPUT61), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1022), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT123), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT125), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1026), .A2(new_n1030), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1001), .A2(new_n949), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1014), .B2(G1348), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(KEYINPUT126), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT126), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1042));
  INV_X1    g617(.A(G1348), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1042), .A2(new_n1043), .B1(new_n1001), .B2(new_n949), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1044), .B2(KEYINPUT60), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1040), .A2(new_n591), .A3(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT126), .B(new_n591), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(KEYINPUT60), .B2(new_n1044), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT61), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n988), .B2(G1996), .ZN(new_n1054));
  INV_X1    g629(.A(new_n984), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n985), .A2(KEYINPUT115), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n985), .A2(KEYINPUT115), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT124), .A3(new_n945), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT58), .B(G1341), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1054), .B(new_n1059), .C1(new_n1001), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n545), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(KEYINPUT59), .A3(new_n545), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1036), .A2(new_n1052), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1044), .A2(new_n591), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1033), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G2078), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT53), .B1(new_n1058), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n728), .B2(new_n1042), .ZN(new_n1073));
  INV_X1    g648(.A(new_n977), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n941), .B1(new_n1074), .B2(KEYINPUT45), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n829), .A2(new_n975), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(KEYINPUT45), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1073), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(G171), .B(KEYINPUT54), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1014), .A2(KEYINPUT120), .A3(new_n690), .ZN(new_n1083));
  INV_X1    g658(.A(G1966), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1042), .B2(G2084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1089), .A2(KEYINPUT127), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1088), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1002), .B1(new_n1093), .B2(G168), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(G168), .B2(new_n1093), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1019), .ZN(new_n1099));
  OR3_X1    g674(.A1(new_n940), .A2(new_n941), .A3(new_n1078), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1073), .B(new_n1080), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1082), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1070), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(KEYINPUT62), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1096), .A2(new_n1105), .A3(new_n1097), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1104), .A2(G171), .A3(new_n1106), .A4(new_n1079), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1018), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1089), .A2(G286), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n993), .A2(new_n1017), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1110), .A2(KEYINPUT121), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT121), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1016), .A2(new_n971), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1010), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1016), .A2(new_n971), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1109), .ZN(new_n1118));
  NOR4_X1   g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1111), .A4(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1112), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n1016), .A3(new_n971), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1004), .A2(new_n1005), .A3(new_n765), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1003), .B1(new_n1122), .B2(new_n996), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT122), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1124), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1119), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(KEYINPUT121), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1126), .B(new_n1127), .C1(new_n1130), .C2(new_n1112), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1108), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G290), .A2(G1986), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1133), .B(new_n1134), .Z(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n943), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT113), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n964), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n968), .B1(new_n1132), .B2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g714(.A1(new_n458), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1141));
  AOI21_X1  g715(.A(new_n1141), .B1(new_n851), .B2(new_n853), .ZN(new_n1142));
  NAND2_X1  g716(.A1(new_n1142), .A2(new_n933), .ZN(G225));
  INV_X1    g717(.A(G225), .ZN(G308));
endmodule


