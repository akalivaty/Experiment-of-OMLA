

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XNOR2_X1 U324 ( .A(n542), .B(n380), .ZN(n387) );
  NOR2_X1 U325 ( .A1(n569), .A2(n509), .ZN(n510) );
  XNOR2_X1 U326 ( .A(n300), .B(n299), .ZN(n304) );
  AND2_X1 U327 ( .A1(G231GAT), .A2(G233GAT), .ZN(n292) );
  AND2_X1 U328 ( .A1(G226GAT), .A2(G233GAT), .ZN(n293) );
  INV_X1 U329 ( .A(KEYINPUT45), .ZN(n505) );
  XNOR2_X1 U330 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U331 ( .A(KEYINPUT27), .ZN(n379) );
  NOR2_X1 U332 ( .A1(n494), .A2(n514), .ZN(n381) );
  XNOR2_X1 U333 ( .A(n379), .B(KEYINPUT97), .ZN(n380) );
  NOR2_X1 U334 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U335 ( .A(n298), .B(n292), .ZN(n299) );
  XNOR2_X1 U336 ( .A(n403), .B(n293), .ZN(n372) );
  NOR2_X1 U337 ( .A1(n546), .A2(n563), .ZN(n548) );
  NOR2_X1 U338 ( .A1(n416), .A2(n579), .ZN(n417) );
  XNOR2_X1 U339 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U340 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U341 ( .A(n451), .B(G29GAT), .ZN(n452) );
  XNOR2_X1 U342 ( .A(n453), .B(n452), .ZN(G1328GAT) );
  XOR2_X1 U343 ( .A(G211GAT), .B(G22GAT), .Z(n295) );
  XOR2_X1 U344 ( .A(G127GAT), .B(G15GAT), .Z(n324) );
  XNOR2_X1 U345 ( .A(n324), .B(KEYINPUT12), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n300) );
  XOR2_X1 U347 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n297) );
  XNOR2_X1 U348 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(G183GAT), .B(G78GAT), .Z(n302) );
  XNOR2_X1 U351 ( .A(G155GAT), .B(G1GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U353 ( .A(n304), .B(n303), .Z(n312) );
  XOR2_X1 U354 ( .A(G71GAT), .B(KEYINPUT70), .Z(n306) );
  XNOR2_X1 U355 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U357 ( .A(KEYINPUT13), .B(n307), .Z(n430) );
  XOR2_X1 U358 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n309) );
  XNOR2_X1 U359 ( .A(G64GAT), .B(G8GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n430), .B(n310), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n574) );
  XOR2_X1 U363 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n314) );
  XNOR2_X1 U364 ( .A(G176GAT), .B(KEYINPUT85), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n332) );
  XOR2_X1 U366 ( .A(G71GAT), .B(G190GAT), .Z(n316) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G99GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U369 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n318) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G169GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U372 ( .A(n320), .B(n319), .Z(n330) );
  XOR2_X1 U373 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(G183GAT), .B(n323), .Z(n373) );
  XNOR2_X1 U377 ( .A(G134GAT), .B(G120GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(KEYINPUT0), .ZN(n351) );
  XOR2_X1 U379 ( .A(n324), .B(n351), .Z(n327) );
  NAND2_X1 U380 ( .A1(G227GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n373), .B(n328), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n516) );
  INV_X1 U385 ( .A(n516), .ZN(n550) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n433) );
  XNOR2_X1 U387 ( .A(G148GAT), .B(G106GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n333), .B(G78GAT), .ZN(n426) );
  XOR2_X1 U389 ( .A(n426), .B(KEYINPUT91), .Z(n335) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U392 ( .A(n433), .B(n336), .Z(n340) );
  XOR2_X1 U393 ( .A(G155GAT), .B(KEYINPUT90), .Z(n338) );
  XNOR2_X1 U394 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n352) );
  XOR2_X1 U396 ( .A(G162GAT), .B(G50GAT), .Z(n399) );
  XNOR2_X1 U397 ( .A(n352), .B(n399), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n350) );
  XOR2_X1 U399 ( .A(G197GAT), .B(KEYINPUT21), .Z(n342) );
  XNOR2_X1 U400 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n343), .B(KEYINPUT89), .Z(n345) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n376) );
  XOR2_X1 U405 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT23), .B(KEYINPUT87), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U408 ( .A(n376), .B(n348), .Z(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n546) );
  XNOR2_X1 U410 ( .A(KEYINPUT28), .B(n546), .ZN(n494) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n371) );
  XOR2_X1 U412 ( .A(KEYINPUT6), .B(G57GAT), .Z(n354) );
  XNOR2_X1 U413 ( .A(G148GAT), .B(G127GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U415 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n356) );
  XNOR2_X1 U416 ( .A(KEYINPUT96), .B(KEYINPUT1), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U418 ( .A(n358), .B(n357), .Z(n369) );
  XOR2_X1 U419 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n360) );
  XNOR2_X1 U420 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n367) );
  XOR2_X1 U422 ( .A(G113GAT), .B(G1GAT), .Z(n441) );
  XOR2_X1 U423 ( .A(G141GAT), .B(G162GAT), .Z(n362) );
  XNOR2_X1 U424 ( .A(G29GAT), .B(G85GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U426 ( .A(n441), .B(n363), .Z(n365) );
  NAND2_X1 U427 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n488) );
  INV_X1 U432 ( .A(n488), .ZN(n544) );
  XOR2_X1 U433 ( .A(G190GAT), .B(G36GAT), .Z(n403) );
  XOR2_X1 U434 ( .A(G8GAT), .B(G169GAT), .Z(n434) );
  XOR2_X1 U435 ( .A(n374), .B(n434), .Z(n378) );
  XNOR2_X1 U436 ( .A(G92GAT), .B(G64GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n375), .B(G176GAT), .ZN(n425) );
  XNOR2_X1 U438 ( .A(n376), .B(n425), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n542) );
  OR2_X1 U440 ( .A1(n544), .A2(n387), .ZN(n514) );
  XOR2_X1 U441 ( .A(KEYINPUT98), .B(n381), .Z(n382) );
  NOR2_X1 U442 ( .A1(n550), .A2(n382), .ZN(n383) );
  XNOR2_X1 U443 ( .A(KEYINPUT99), .B(n383), .ZN(n394) );
  NOR2_X1 U444 ( .A1(n542), .A2(n516), .ZN(n384) );
  NOR2_X1 U445 ( .A1(n546), .A2(n384), .ZN(n385) );
  XOR2_X1 U446 ( .A(KEYINPUT25), .B(n385), .Z(n390) );
  NAND2_X1 U447 ( .A1(n516), .A2(n546), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n386), .B(KEYINPUT26), .ZN(n564) );
  NOR2_X1 U449 ( .A1(n564), .A2(n387), .ZN(n388) );
  XNOR2_X1 U450 ( .A(KEYINPUT100), .B(n388), .ZN(n389) );
  NOR2_X1 U451 ( .A1(n390), .A2(n389), .ZN(n391) );
  NOR2_X1 U452 ( .A1(n488), .A2(n391), .ZN(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT101), .B(n392), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n394), .A2(n393), .ZN(n456) );
  NAND2_X1 U455 ( .A1(n574), .A2(n456), .ZN(n395) );
  XNOR2_X1 U456 ( .A(KEYINPUT104), .B(n395), .ZN(n416) );
  XOR2_X1 U457 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n397) );
  XNOR2_X1 U458 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U460 ( .A(n398), .B(G106GAT), .Z(n401) );
  XNOR2_X1 U461 ( .A(n399), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n407) );
  XNOR2_X1 U463 ( .A(G85GAT), .B(KEYINPUT72), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n402), .B(G99GAT), .ZN(n418) );
  XOR2_X1 U465 ( .A(n418), .B(n403), .Z(n405) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U468 ( .A(n407), .B(n406), .Z(n415) );
  XOR2_X1 U469 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n409) );
  XNOR2_X1 U470 ( .A(KEYINPUT68), .B(G43GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(n410), .ZN(n446) );
  XOR2_X1 U473 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n412) );
  XNOR2_X1 U474 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U476 ( .A(n446), .B(n413), .Z(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n526) );
  XOR2_X1 U478 ( .A(KEYINPUT36), .B(n526), .Z(n579) );
  XNOR2_X1 U479 ( .A(n417), .B(KEYINPUT37), .ZN(n487) );
  XOR2_X1 U480 ( .A(KEYINPUT31), .B(n418), .Z(n420) );
  NAND2_X1 U481 ( .A1(G230GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U483 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n422) );
  XNOR2_X1 U484 ( .A(G120GAT), .B(G204GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U486 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n569) );
  XOR2_X1 U490 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n432) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(G197GAT), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n445) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n436) );
  XNOR2_X1 U494 ( .A(G36GAT), .B(G50GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n438) );
  NAND2_X1 U497 ( .A1(G229GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U500 ( .A(n441), .B(KEYINPUT66), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n565) );
  NOR2_X1 U504 ( .A1(n569), .A2(n565), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n448), .B(KEYINPUT73), .ZN(n458) );
  NOR2_X1 U506 ( .A1(n487), .A2(n458), .ZN(n450) );
  XNOR2_X1 U507 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n473) );
  NOR2_X1 U509 ( .A1(n473), .A2(n544), .ZN(n453) );
  XNOR2_X1 U510 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n451) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n460) );
  NOR2_X1 U512 ( .A1(n526), .A2(n574), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT16), .B(n454), .Z(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT81), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n457), .A2(n456), .ZN(n477) );
  NOR2_X1 U516 ( .A1(n458), .A2(n477), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n465), .A2(n488), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U519 ( .A(G1GAT), .B(n461), .Z(G1324GAT) );
  INV_X1 U520 ( .A(n542), .ZN(n490) );
  NAND2_X1 U521 ( .A1(n490), .A2(n465), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U523 ( .A(G15GAT), .B(KEYINPUT35), .Z(n464) );
  NAND2_X1 U524 ( .A1(n465), .A2(n550), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  XOR2_X1 U526 ( .A(G22GAT), .B(KEYINPUT103), .Z(n467) );
  NAND2_X1 U527 ( .A1(n465), .A2(n494), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(G1327GAT) );
  NOR2_X1 U529 ( .A1(n542), .A2(n473), .ZN(n468) );
  XOR2_X1 U530 ( .A(G36GAT), .B(n468), .Z(G1329GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n470) );
  XNOR2_X1 U532 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n469) );
  XNOR2_X1 U533 ( .A(n470), .B(n469), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n473), .A2(n516), .ZN(n471) );
  XOR2_X1 U535 ( .A(n472), .B(n471), .Z(G1330GAT) );
  INV_X1 U536 ( .A(n494), .ZN(n518) );
  NOR2_X1 U537 ( .A1(n473), .A2(n518), .ZN(n474) );
  XOR2_X1 U538 ( .A(G50GAT), .B(n474), .Z(G1331GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n475) );
  XNOR2_X1 U541 ( .A(n475), .B(n569), .ZN(n552) );
  INV_X1 U542 ( .A(n552), .ZN(n476) );
  NAND2_X1 U543 ( .A1(n476), .A2(n565), .ZN(n486) );
  NOR2_X1 U544 ( .A1(n486), .A2(n477), .ZN(n483) );
  NAND2_X1 U545 ( .A1(n483), .A2(n488), .ZN(n478) );
  XNOR2_X1 U546 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U547 ( .A(G57GAT), .B(n480), .ZN(G1332GAT) );
  NAND2_X1 U548 ( .A1(n490), .A2(n483), .ZN(n481) );
  XNOR2_X1 U549 ( .A(n481), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U550 ( .A1(n483), .A2(n550), .ZN(n482) );
  XNOR2_X1 U551 ( .A(n482), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U552 ( .A(G78GAT), .B(KEYINPUT43), .Z(n485) );
  NAND2_X1 U553 ( .A1(n483), .A2(n494), .ZN(n484) );
  XNOR2_X1 U554 ( .A(n485), .B(n484), .ZN(G1335GAT) );
  NOR2_X1 U555 ( .A1(n487), .A2(n486), .ZN(n495) );
  NAND2_X1 U556 ( .A1(n488), .A2(n495), .ZN(n489) );
  XNOR2_X1 U557 ( .A(G85GAT), .B(n489), .ZN(G1336GAT) );
  NAND2_X1 U558 ( .A1(n495), .A2(n490), .ZN(n491) );
  XNOR2_X1 U559 ( .A(G92GAT), .B(n491), .ZN(G1337GAT) );
  NAND2_X1 U560 ( .A1(n495), .A2(n550), .ZN(n492) );
  XNOR2_X1 U561 ( .A(n492), .B(KEYINPUT110), .ZN(n493) );
  XNOR2_X1 U562 ( .A(G99GAT), .B(n493), .ZN(G1338GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n497) );
  NAND2_X1 U564 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(n498), .ZN(G1339GAT) );
  NOR2_X1 U567 ( .A1(n565), .A2(n552), .ZN(n500) );
  XNOR2_X1 U568 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n499) );
  XNOR2_X1 U569 ( .A(n500), .B(n499), .ZN(n501) );
  NOR2_X1 U570 ( .A1(n526), .A2(n501), .ZN(n502) );
  NAND2_X1 U571 ( .A1(n574), .A2(n502), .ZN(n504) );
  XOR2_X1 U572 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n503) );
  XNOR2_X1 U573 ( .A(n504), .B(n503), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n579), .A2(n574), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(KEYINPUT65), .ZN(n508) );
  NAND2_X1 U576 ( .A1(n508), .A2(n565), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(KEYINPUT114), .ZN(n511) );
  NOR2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT48), .B(n513), .ZN(n541) );
  NOR2_X1 U580 ( .A1(n541), .A2(n514), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(KEYINPUT115), .ZN(n531) );
  NOR2_X1 U582 ( .A1(n516), .A2(n531), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT116), .ZN(n519) );
  NAND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n565), .A2(n527), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1340GAT) );
  NOR2_X1 U588 ( .A1(n552), .A2(n527), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1341GAT) );
  NOR2_X1 U591 ( .A1(n574), .A2(n527), .ZN(n524) );
  XOR2_X1 U592 ( .A(KEYINPUT50), .B(n524), .Z(n525) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(n525), .ZN(G1342GAT) );
  INV_X1 U594 ( .A(n526), .ZN(n560) );
  NOR2_X1 U595 ( .A1(n560), .A2(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(n530), .ZN(G1343GAT) );
  OR2_X1 U599 ( .A1(n564), .A2(n531), .ZN(n539) );
  NOR2_X1 U600 ( .A1(n565), .A2(n539), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(G1344GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n535) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(n537) );
  NOR2_X1 U606 ( .A1(n552), .A2(n539), .ZN(n536) );
  XOR2_X1 U607 ( .A(n537), .B(n536), .Z(G1345GAT) );
  NOR2_X1 U608 ( .A1(n574), .A2(n539), .ZN(n538) );
  XOR2_X1 U609 ( .A(G155GAT), .B(n538), .Z(G1346GAT) );
  NOR2_X1 U610 ( .A1(n560), .A2(n539), .ZN(n540) );
  XOR2_X1 U611 ( .A(G162GAT), .B(n540), .Z(G1347GAT) );
  XNOR2_X1 U612 ( .A(n543), .B(KEYINPUT54), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n563) );
  XNOR2_X1 U614 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n559) );
  NOR2_X1 U617 ( .A1(n565), .A2(n559), .ZN(n551) );
  XOR2_X1 U618 ( .A(G169GAT), .B(n551), .Z(G1348GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n559), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n554) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(KEYINPUT122), .B(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n574), .A2(n559), .ZN(n558) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n558), .Z(G1350GAT) );
  XOR2_X1 U627 ( .A(G190GAT), .B(n561), .Z(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT58), .B(n562), .ZN(G1351GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n570) );
  INV_X1 U630 ( .A(n570), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n565), .A2(n578), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n578), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

