

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767;

  AND2_X1 U366 ( .A1(n364), .A2(n619), .ZN(n628) );
  XNOR2_X1 U367 ( .A(n347), .B(KEYINPUT33), .ZN(n715) );
  NOR2_X1 U368 ( .A1(n580), .A2(n579), .ZN(n582) );
  NOR2_X1 U369 ( .A1(n556), .A2(n543), .ZN(n347) );
  BUF_X1 U370 ( .A(n693), .Z(n348) );
  NOR2_X1 U371 ( .A1(n555), .A2(n554), .ZN(n675) );
  NOR2_X1 U372 ( .A1(n378), .A2(n692), .ZN(n560) );
  XNOR2_X1 U373 ( .A(n589), .B(KEYINPUT1), .ZN(n693) );
  XOR2_X1 U374 ( .A(n491), .B(KEYINPUT92), .Z(n359) );
  XNOR2_X1 U375 ( .A(n346), .B(n518), .ZN(n654) );
  XNOR2_X1 U376 ( .A(n509), .B(n504), .ZN(n346) );
  XNOR2_X1 U377 ( .A(G128), .B(G143), .ZN(n475) );
  XNOR2_X2 U378 ( .A(n402), .B(n401), .ZN(n632) );
  XNOR2_X1 U379 ( .A(n548), .B(n363), .ZN(n549) );
  NOR2_X1 U380 ( .A1(n635), .A2(n738), .ZN(n637) );
  XNOR2_X2 U381 ( .A(G902), .B(KEYINPUT15), .ZN(n621) );
  NOR2_X1 U382 ( .A1(n766), .A2(n765), .ZN(n435) );
  NAND2_X1 U383 ( .A1(n572), .A2(n687), .ZN(n575) );
  XNOR2_X1 U384 ( .A(n513), .B(n512), .ZN(n572) );
  NAND2_X2 U385 ( .A1(n595), .A2(n497), .ZN(n499) );
  XOR2_X1 U386 ( .A(G113), .B(G104), .Z(n451) );
  BUF_X1 U387 ( .A(n628), .Z(n757) );
  BUF_X1 U388 ( .A(G143), .Z(n672) );
  NOR2_X2 U389 ( .A1(n728), .A2(G902), .ZN(n520) );
  INV_X1 U390 ( .A(KEYINPUT76), .ZN(n581) );
  INV_X1 U391 ( .A(G953), .ZN(n480) );
  XNOR2_X1 U392 ( .A(n415), .B(n421), .ZN(n714) );
  INV_X1 U393 ( .A(n693), .ZN(n349) );
  XOR2_X1 U394 ( .A(KEYINPUT65), .B(n623), .Z(n624) );
  XNOR2_X1 U395 ( .A(n476), .B(n449), .ZN(n756) );
  XNOR2_X1 U396 ( .A(n419), .B(n356), .ZN(n414) );
  XNOR2_X1 U397 ( .A(n448), .B(G125), .ZN(n476) );
  XNOR2_X1 U398 ( .A(n470), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U399 ( .A(G122), .B(KEYINPUT101), .ZN(n455) );
  XNOR2_X1 U400 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n424) );
  NOR2_X1 U401 ( .A1(n733), .A2(n738), .ZN(n420) );
  XNOR2_X1 U402 ( .A(n475), .B(KEYINPUT4), .ZN(n503) );
  NAND2_X1 U403 ( .A1(n390), .A2(G469), .ZN(n732) );
  XNOR2_X1 U404 ( .A(n418), .B(n501), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n418), .B(n501), .ZN(n566) );
  NOR2_X1 U406 ( .A1(n657), .A2(n738), .ZN(n659) );
  NAND2_X1 U407 ( .A1(n569), .A2(n568), .ZN(n351) );
  XNOR2_X2 U408 ( .A(n552), .B(n551), .ZN(n569) );
  BUF_X1 U409 ( .A(n558), .Z(n352) );
  XNOR2_X1 U410 ( .A(n351), .B(n570), .ZN(n353) );
  XNOR2_X2 U411 ( .A(n520), .B(G469), .ZN(n589) );
  NAND2_X1 U412 ( .A1(n566), .A2(n535), .ZN(n438) );
  NOR2_X1 U413 ( .A1(n377), .A2(n678), .ZN(n374) );
  OR2_X1 U414 ( .A1(n662), .A2(n660), .ZN(n377) );
  XNOR2_X1 U415 ( .A(n511), .B(G472), .ZN(n512) );
  INV_X1 U416 ( .A(KEYINPUT72), .ZN(n511) );
  INV_X1 U417 ( .A(G146), .ZN(n448) );
  XNOR2_X1 U418 ( .A(n628), .B(n620), .ZN(n371) );
  XNOR2_X1 U419 ( .A(n439), .B(KEYINPUT38), .ZN(n684) );
  OR2_X1 U420 ( .A1(n684), .A2(n429), .ZN(n428) );
  NAND2_X1 U421 ( .A1(n354), .A2(n611), .ZN(n433) );
  NAND2_X1 U422 ( .A1(n621), .A2(KEYINPUT84), .ZN(n367) );
  NOR2_X1 U423 ( .A1(G953), .A2(G237), .ZN(n505) );
  XNOR2_X1 U424 ( .A(G101), .B(KEYINPUT67), .ZN(n474) );
  XNOR2_X1 U425 ( .A(n503), .B(n440), .ZN(n755) );
  XNOR2_X1 U426 ( .A(n502), .B(G137), .ZN(n440) );
  XNOR2_X1 U427 ( .A(G134), .B(G131), .ZN(n502) );
  XNOR2_X1 U428 ( .A(n463), .B(G107), .ZN(n472) );
  INV_X1 U429 ( .A(G122), .ZN(n463) );
  XNOR2_X1 U430 ( .A(n442), .B(n441), .ZN(n527) );
  INV_X1 U431 ( .A(KEYINPUT8), .ZN(n441) );
  NAND2_X1 U432 ( .A1(n480), .A2(G234), .ZN(n442) );
  INV_X1 U433 ( .A(G140), .ZN(n514) );
  XNOR2_X1 U434 ( .A(n755), .B(G146), .ZN(n518) );
  INV_X1 U435 ( .A(KEYINPUT48), .ZN(n430) );
  INV_X1 U436 ( .A(G237), .ZN(n489) );
  INV_X1 U437 ( .A(G902), .ZN(n490) );
  AND2_X1 U438 ( .A1(n422), .A2(n684), .ZN(n690) );
  INV_X1 U439 ( .A(n685), .ZN(n422) );
  XNOR2_X1 U440 ( .A(G110), .B(KEYINPUT95), .ZN(n521) );
  XNOR2_X1 U441 ( .A(G140), .B(KEYINPUT10), .ZN(n449) );
  XNOR2_X1 U442 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U443 ( .A(G119), .ZN(n523) );
  XNOR2_X1 U444 ( .A(G128), .B(G137), .ZN(n524) );
  AND2_X1 U445 ( .A1(n684), .A2(n429), .ZN(n427) );
  AND2_X1 U446 ( .A1(n396), .A2(n675), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n557), .B(KEYINPUT98), .ZN(n705) );
  XNOR2_X1 U448 ( .A(n410), .B(n408), .ZN(n447) );
  XNOR2_X1 U449 ( .A(n409), .B(KEYINPUT28), .ZN(n408) );
  XNOR2_X1 U450 ( .A(n533), .B(n532), .ZN(n696) );
  NOR2_X1 U451 ( .A1(n632), .A2(G902), .ZN(n533) );
  XNOR2_X1 U452 ( .A(n460), .B(G475), .ZN(n425) );
  AND2_X1 U453 ( .A1(n407), .A2(G953), .ZN(n406) );
  XNOR2_X1 U454 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n471) );
  XNOR2_X1 U455 ( .A(n423), .B(n361), .ZN(n456) );
  XNOR2_X1 U456 ( .A(n455), .B(n424), .ZN(n423) );
  XNOR2_X1 U457 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n453) );
  XOR2_X1 U458 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n454) );
  XNOR2_X1 U459 ( .A(KEYINPUT88), .B(KEYINPUT77), .ZN(n478) );
  XOR2_X1 U460 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n479) );
  XNOR2_X1 U461 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n482) );
  XNOR2_X1 U462 ( .A(n571), .B(n570), .ZN(n629) );
  NAND2_X1 U463 ( .A1(G237), .A2(G234), .ZN(n493) );
  NAND2_X1 U464 ( .A1(n587), .A2(n696), .ZN(n604) );
  XNOR2_X1 U465 ( .A(n575), .B(n574), .ZN(n578) );
  INV_X1 U466 ( .A(KEYINPUT113), .ZN(n409) );
  NOR2_X1 U467 ( .A1(n604), .A2(n588), .ZN(n410) );
  XNOR2_X1 U468 ( .A(G478), .B(n465), .ZN(n553) );
  OR2_X1 U469 ( .A1(n696), .A2(n697), .ZN(n692) );
  XNOR2_X1 U470 ( .A(G134), .B(G116), .ZN(n464) );
  XNOR2_X1 U471 ( .A(n516), .B(n517), .ZN(n436) );
  BUF_X1 U472 ( .A(n353), .Z(n739) );
  INV_X1 U473 ( .A(KEYINPUT41), .ZN(n421) );
  NAND2_X1 U474 ( .A1(n690), .A2(n687), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n528), .B(n526), .ZN(n402) );
  XNOR2_X1 U476 ( .A(n756), .B(n525), .ZN(n401) );
  XNOR2_X1 U477 ( .A(n445), .B(n443), .ZN(n736) );
  XNOR2_X1 U478 ( .A(n444), .B(n462), .ZN(n443) );
  XNOR2_X1 U479 ( .A(n461), .B(n446), .ZN(n445) );
  XOR2_X1 U480 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n462) );
  AND2_X1 U481 ( .A1(n618), .A2(n439), .ZN(n638) );
  NAND2_X1 U482 ( .A1(n355), .A2(n397), .ZN(n612) );
  NAND2_X1 U483 ( .A1(n399), .A2(n398), .ZN(n584) );
  NAND2_X1 U484 ( .A1(n400), .A2(n360), .ZN(n398) );
  XNOR2_X1 U485 ( .A(n559), .B(KEYINPUT31), .ZN(n678) );
  NOR2_X1 U486 ( .A1(n597), .A2(n596), .ZN(n673) );
  OR2_X1 U487 ( .A1(n403), .A2(KEYINPUT47), .ZN(n354) );
  AND2_X1 U488 ( .A1(n394), .A2(n428), .ZN(n355) );
  XOR2_X1 U489 ( .A(G119), .B(G116), .Z(n356) );
  OR2_X1 U490 ( .A1(n713), .A2(G953), .ZN(n357) );
  AND2_X1 U491 ( .A1(n404), .A2(n357), .ZN(n358) );
  AND2_X1 U492 ( .A1(n427), .A2(n675), .ZN(n360) );
  AND2_X1 U493 ( .A1(G214), .A2(n505), .ZN(n361) );
  XOR2_X1 U494 ( .A(KEYINPUT106), .B(KEYINPUT6), .Z(n362) );
  XOR2_X1 U495 ( .A(n547), .B(n546), .Z(n363) );
  INV_X1 U496 ( .A(KEYINPUT84), .ZN(n372) );
  XNOR2_X2 U497 ( .A(n608), .B(KEYINPUT19), .ZN(n595) );
  NAND2_X2 U498 ( .A1(n417), .A2(n687), .ZN(n608) );
  XNOR2_X2 U499 ( .A(n412), .B(n359), .ZN(n417) );
  NAND2_X1 U500 ( .A1(n629), .A2(KEYINPUT84), .ZN(n368) );
  XNOR2_X1 U501 ( .A(n431), .B(n430), .ZN(n364) );
  NAND2_X1 U502 ( .A1(n365), .A2(n371), .ZN(n625) );
  NOR2_X1 U503 ( .A1(n366), .A2(n369), .ZN(n365) );
  NAND2_X1 U504 ( .A1(n368), .A2(n367), .ZN(n366) );
  NOR2_X1 U505 ( .A1(n353), .A2(n370), .ZN(n369) );
  NAND2_X1 U506 ( .A1(n622), .A2(n372), .ZN(n370) );
  XNOR2_X1 U507 ( .A(n458), .B(n459), .ZN(n640) );
  BUF_X1 U508 ( .A(n748), .Z(n373) );
  NOR2_X1 U509 ( .A1(n374), .A2(n375), .ZN(n567) );
  AND2_X1 U510 ( .A1(n376), .A2(n598), .ZN(n375) );
  INV_X1 U511 ( .A(n660), .ZN(n376) );
  BUF_X1 U512 ( .A(n589), .Z(n378) );
  NAND2_X1 U513 ( .A1(n414), .A2(n413), .ZN(n380) );
  NAND2_X1 U514 ( .A1(n379), .A2(n473), .ZN(n381) );
  NAND2_X1 U515 ( .A1(n380), .A2(n381), .ZN(n747) );
  INV_X1 U516 ( .A(n414), .ZN(n379) );
  NOR2_X2 U517 ( .A1(n630), .A2(n739), .ZN(n724) );
  XNOR2_X2 U518 ( .A(n499), .B(n498), .ZN(n558) );
  NAND2_X1 U519 ( .A1(n625), .A2(n624), .ZN(n627) );
  OR2_X2 U520 ( .A1(n640), .A2(G902), .ZN(n426) );
  XNOR2_X1 U521 ( .A(n747), .B(n411), .ZN(n488) );
  BUF_X1 U522 ( .A(n755), .Z(n382) );
  BUF_X1 U523 ( .A(n647), .Z(n383) );
  XNOR2_X1 U524 ( .A(n488), .B(n487), .ZN(n647) );
  BUF_X1 U525 ( .A(n543), .Z(n603) );
  XNOR2_X1 U526 ( .A(n588), .B(n362), .ZN(n543) );
  XNOR2_X1 U527 ( .A(n475), .B(KEYINPUT9), .ZN(n444) );
  BUF_X1 U528 ( .A(n595), .Z(n385) );
  INV_X1 U529 ( .A(n439), .ZN(n386) );
  BUF_X1 U530 ( .A(n608), .Z(n387) );
  XNOR2_X1 U531 ( .A(n549), .B(G122), .ZN(G24) );
  BUF_X1 U532 ( .A(n539), .Z(n388) );
  NOR2_X1 U533 ( .A1(n631), .A2(n724), .ZN(n389) );
  NOR2_X2 U534 ( .A1(n631), .A2(n724), .ZN(n390) );
  INV_X1 U535 ( .A(n561), .ZN(n391) );
  NOR2_X2 U536 ( .A1(n631), .A2(n724), .ZN(n734) );
  NAND2_X1 U537 ( .A1(n647), .A2(n621), .ZN(n412) );
  NAND2_X1 U538 ( .A1(n392), .A2(n395), .ZN(n399) );
  NAND2_X1 U539 ( .A1(n393), .A2(n428), .ZN(n392) );
  INV_X1 U540 ( .A(n594), .ZN(n393) );
  INV_X1 U541 ( .A(n594), .ZN(n400) );
  NAND2_X1 U542 ( .A1(n594), .A2(n583), .ZN(n394) );
  NAND2_X1 U543 ( .A1(n428), .A2(n429), .ZN(n396) );
  NAND2_X1 U544 ( .A1(n400), .A2(n427), .ZN(n397) );
  NAND2_X1 U545 ( .A1(n403), .A2(KEYINPUT47), .ZN(n599) );
  NAND2_X1 U546 ( .A1(n673), .A2(n683), .ZN(n403) );
  XNOR2_X1 U547 ( .A(n405), .B(KEYINPUT110), .ZN(n404) );
  NAND2_X1 U548 ( .A1(n576), .A2(n406), .ZN(n405) );
  INV_X1 U549 ( .A(G900), .ZN(n407) );
  INV_X1 U550 ( .A(n572), .ZN(n588) );
  XNOR2_X1 U551 ( .A(n411), .B(n436), .ZN(n519) );
  XNOR2_X2 U552 ( .A(n437), .B(n504), .ZN(n411) );
  INV_X1 U553 ( .A(n473), .ZN(n413) );
  XNOR2_X1 U554 ( .A(n414), .B(n508), .ZN(n509) );
  XNOR2_X2 U555 ( .A(n416), .B(G110), .ZN(n748) );
  XNOR2_X2 U556 ( .A(G104), .B(KEYINPUT89), .ZN(n416) );
  INV_X1 U557 ( .A(n417), .ZN(n439) );
  NAND2_X1 U558 ( .A1(n592), .A2(n386), .ZN(n593) );
  NAND2_X1 U559 ( .A1(n558), .A2(n500), .ZN(n418) );
  XNOR2_X1 U560 ( .A(n420), .B(KEYINPUT122), .ZN(G54) );
  XNOR2_X2 U561 ( .A(n426), .B(n425), .ZN(n554) );
  INV_X1 U562 ( .A(n583), .ZN(n429) );
  NAND2_X1 U563 ( .A1(n434), .A2(n432), .ZN(n431) );
  NOR2_X1 U564 ( .A1(n602), .A2(n433), .ZN(n432) );
  XNOR2_X1 U565 ( .A(n435), .B(KEYINPUT46), .ZN(n434) );
  XNOR2_X2 U566 ( .A(n748), .B(KEYINPUT70), .ZN(n437) );
  INV_X1 U567 ( .A(n388), .ZN(n639) );
  XNOR2_X2 U568 ( .A(n438), .B(KEYINPUT32), .ZN(n539) );
  INV_X1 U569 ( .A(n588), .ZN(n703) );
  XNOR2_X2 U570 ( .A(KEYINPUT107), .B(n466), .ZN(n685) );
  AND2_X2 U571 ( .A1(n554), .A2(n553), .ZN(n466) );
  XNOR2_X2 U572 ( .A(n627), .B(n626), .ZN(n631) );
  XOR2_X1 U573 ( .A(n472), .B(n464), .Z(n446) );
  INV_X1 U574 ( .A(KEYINPUT86), .ZN(n540) );
  INV_X1 U575 ( .A(n681), .ZN(n611) );
  XNOR2_X1 U576 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U577 ( .A(KEYINPUT30), .ZN(n573) );
  XNOR2_X1 U578 ( .A(n573), .B(KEYINPUT112), .ZN(n574) );
  INV_X1 U579 ( .A(KEYINPUT123), .ZN(n636) );
  XNOR2_X1 U580 ( .A(n672), .B(G131), .ZN(n450) );
  XNOR2_X1 U581 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U582 ( .A(n756), .B(n452), .Z(n459) );
  XNOR2_X1 U583 ( .A(n454), .B(n453), .ZN(n457) );
  XOR2_X1 U584 ( .A(n457), .B(n456), .Z(n458) );
  XNOR2_X1 U585 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n460) );
  NAND2_X1 U586 ( .A1(G217), .A2(n527), .ZN(n461) );
  NOR2_X1 U587 ( .A1(G902), .A2(n736), .ZN(n465) );
  NAND2_X1 U588 ( .A1(n621), .A2(G234), .ZN(n467) );
  XNOR2_X1 U589 ( .A(n467), .B(KEYINPUT20), .ZN(n529) );
  NAND2_X1 U590 ( .A1(G221), .A2(n529), .ZN(n468) );
  XNOR2_X1 U591 ( .A(KEYINPUT21), .B(n468), .ZN(n697) );
  NOR2_X1 U592 ( .A1(n685), .A2(n697), .ZN(n469) );
  XNOR2_X1 U593 ( .A(n469), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X2 U594 ( .A(G113), .B(KEYINPUT69), .ZN(n470) );
  XNOR2_X1 U595 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U596 ( .A(n474), .B(KEYINPUT66), .ZN(n504) );
  BUF_X1 U597 ( .A(n503), .Z(n477) );
  XNOR2_X1 U598 ( .A(n477), .B(n476), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n479), .B(n478), .ZN(n484) );
  NAND2_X1 U600 ( .A1(n480), .A2(G224), .ZN(n481) );
  XNOR2_X1 U601 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U602 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U603 ( .A(n486), .B(n485), .ZN(n487) );
  NAND2_X1 U604 ( .A1(n490), .A2(n489), .ZN(n492) );
  NAND2_X1 U605 ( .A1(n492), .A2(G210), .ZN(n491) );
  NAND2_X1 U606 ( .A1(n492), .A2(G214), .ZN(n687) );
  XNOR2_X1 U607 ( .A(n493), .B(KEYINPUT14), .ZN(n495) );
  NAND2_X1 U608 ( .A1(n495), .A2(G902), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n494), .B(KEYINPUT93), .ZN(n576) );
  NOR2_X1 U610 ( .A1(G898), .A2(n480), .ZN(n751) );
  NAND2_X1 U611 ( .A1(n576), .A2(n751), .ZN(n496) );
  NAND2_X1 U612 ( .A1(G952), .A2(n495), .ZN(n713) );
  NAND2_X1 U613 ( .A1(n496), .A2(n357), .ZN(n497) );
  INV_X1 U614 ( .A(KEYINPUT0), .ZN(n498) );
  INV_X1 U615 ( .A(KEYINPUT22), .ZN(n501) );
  XOR2_X1 U616 ( .A(KEYINPUT74), .B(KEYINPUT5), .Z(n507) );
  NAND2_X1 U617 ( .A1(n505), .A2(G210), .ZN(n506) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U619 ( .A1(G902), .A2(n654), .ZN(n513) );
  XNOR2_X1 U620 ( .A(G107), .B(KEYINPUT94), .ZN(n517) );
  NAND2_X1 U621 ( .A1(G227), .A2(n480), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n519), .B(n518), .ZN(n728) );
  XOR2_X1 U623 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n522) );
  XNOR2_X1 U624 ( .A(n522), .B(n521), .ZN(n526) );
  NAND2_X1 U625 ( .A1(G221), .A2(n527), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n529), .A2(G217), .ZN(n531) );
  XOR2_X1 U627 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n530) );
  XNOR2_X1 U628 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U629 ( .A(n696), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n348), .A2(n563), .ZN(n534) );
  AND2_X1 U631 ( .A1(n603), .A2(n534), .ZN(n535) );
  NAND2_X1 U632 ( .A1(n348), .A2(n696), .ZN(n536) );
  NOR2_X1 U633 ( .A1(n703), .A2(n536), .ZN(n537) );
  AND2_X1 U634 ( .A1(n350), .A2(n537), .ZN(n667) );
  INV_X1 U635 ( .A(n667), .ZN(n538) );
  NAND2_X1 U636 ( .A1(n539), .A2(n538), .ZN(n541) );
  XNOR2_X1 U637 ( .A(n541), .B(n540), .ZN(n550) );
  INV_X1 U638 ( .A(n692), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n542), .A2(n349), .ZN(n556) );
  INV_X1 U640 ( .A(n352), .ZN(n561) );
  NOR2_X2 U641 ( .A1(n715), .A2(n561), .ZN(n544) );
  XNOR2_X1 U642 ( .A(n544), .B(KEYINPUT34), .ZN(n545) );
  NOR2_X1 U643 ( .A1(n554), .A2(n553), .ZN(n592) );
  NAND2_X1 U644 ( .A1(n545), .A2(n592), .ZN(n548) );
  XNOR2_X1 U645 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n547) );
  INV_X1 U646 ( .A(KEYINPUT78), .ZN(n546) );
  NAND2_X1 U647 ( .A1(n550), .A2(n549), .ZN(n552) );
  INV_X1 U648 ( .A(KEYINPUT44), .ZN(n551) );
  INV_X1 U649 ( .A(n553), .ZN(n555) );
  AND2_X1 U650 ( .A1(n555), .A2(n554), .ZN(n677) );
  NOR2_X1 U651 ( .A1(n677), .A2(n675), .ZN(n598) );
  NOR2_X1 U652 ( .A1(n556), .A2(n588), .ZN(n557) );
  NAND2_X1 U653 ( .A1(n705), .A2(n391), .ZN(n559) );
  XNOR2_X1 U654 ( .A(n560), .B(KEYINPUT97), .ZN(n580) );
  OR2_X1 U655 ( .A1(n703), .A2(n580), .ZN(n562) );
  NOR2_X1 U656 ( .A1(n562), .A2(n561), .ZN(n662) );
  AND2_X1 U657 ( .A1(n348), .A2(n563), .ZN(n564) );
  AND2_X1 U658 ( .A1(n603), .A2(n564), .ZN(n565) );
  AND2_X1 U659 ( .A1(n350), .A2(n565), .ZN(n660) );
  XNOR2_X1 U660 ( .A(n567), .B(KEYINPUT109), .ZN(n568) );
  NAND2_X1 U661 ( .A1(n569), .A2(n568), .ZN(n571) );
  INV_X1 U662 ( .A(KEYINPUT45), .ZN(n570) );
  XNOR2_X1 U663 ( .A(KEYINPUT79), .B(n358), .ZN(n577) );
  INV_X1 U664 ( .A(n577), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X2 U666 ( .A(n582), .B(n581), .ZN(n594) );
  XOR2_X1 U667 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n583) );
  XNOR2_X1 U668 ( .A(n584), .B(KEYINPUT40), .ZN(n766) );
  NOR2_X1 U669 ( .A1(n697), .A2(n585), .ZN(n586) );
  XNOR2_X1 U670 ( .A(n586), .B(KEYINPUT68), .ZN(n587) );
  INV_X1 U671 ( .A(n378), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n447), .A2(n590), .ZN(n597) );
  NOR2_X1 U673 ( .A1(n597), .A2(n714), .ZN(n591) );
  XNOR2_X1 U674 ( .A(KEYINPUT42), .B(n591), .ZN(n765) );
  NOR2_X1 U675 ( .A1(n594), .A2(n593), .ZN(n671) );
  XNOR2_X1 U676 ( .A(n671), .B(KEYINPUT83), .ZN(n600) );
  INV_X1 U677 ( .A(n385), .ZN(n596) );
  INV_X1 U678 ( .A(n598), .ZN(n683) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n601), .B(KEYINPUT82), .ZN(n602) );
  INV_X1 U681 ( .A(n603), .ZN(n607) );
  INV_X1 U682 ( .A(n675), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n614), .A2(n387), .ZN(n609) );
  XOR2_X1 U686 ( .A(KEYINPUT36), .B(n609), .Z(n610) );
  NOR2_X1 U687 ( .A1(n348), .A2(n610), .ZN(n681) );
  NAND2_X1 U688 ( .A1(n612), .A2(n677), .ZN(n613) );
  XOR2_X1 U689 ( .A(KEYINPUT114), .B(n613), .Z(n767) );
  XOR2_X1 U690 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n617) );
  NOR2_X1 U691 ( .A1(n349), .A2(n614), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n615), .A2(n687), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n617), .B(n616), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n767), .A2(n638), .ZN(n619) );
  INV_X1 U695 ( .A(KEYINPUT75), .ZN(n620) );
  INV_X1 U696 ( .A(n621), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n622), .A2(KEYINPUT2), .ZN(n623) );
  INV_X1 U698 ( .A(KEYINPUT64), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n757), .A2(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n734), .A2(G217), .ZN(n633) );
  XNOR2_X1 U701 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U702 ( .A(G952), .ZN(n634) );
  AND2_X1 U703 ( .A1(n634), .A2(G953), .ZN(n738) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(G66) );
  XOR2_X1 U705 ( .A(n638), .B(G140), .Z(G42) );
  XOR2_X1 U706 ( .A(n639), .B(G119), .Z(G21) );
  NAND2_X1 U707 ( .A1(n389), .A2(G475), .ZN(n642) );
  XNOR2_X1 U708 ( .A(n640), .B(KEYINPUT59), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n642), .B(n641), .ZN(n643) );
  INV_X1 U710 ( .A(n738), .ZN(n650) );
  NAND2_X1 U711 ( .A1(n643), .A2(n650), .ZN(n645) );
  INV_X1 U712 ( .A(KEYINPUT60), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n645), .B(n644), .ZN(G60) );
  NAND2_X1 U714 ( .A1(n390), .A2(G210), .ZN(n649) );
  XOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n646) );
  XNOR2_X1 U716 ( .A(n383), .B(n646), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n649), .B(n648), .ZN(n651) );
  NAND2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n653) );
  INV_X1 U719 ( .A(KEYINPUT56), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n653), .B(n652), .ZN(G51) );
  NAND2_X1 U721 ( .A1(n734), .A2(G472), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT62), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U724 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n659), .B(n658), .ZN(G57) );
  XOR2_X1 U726 ( .A(G101), .B(n660), .Z(G3) );
  NAND2_X1 U727 ( .A1(n662), .A2(n675), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n661), .B(G104), .ZN(G6) );
  XOR2_X1 U729 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n664) );
  NAND2_X1 U730 ( .A1(n662), .A2(n677), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n666) );
  XOR2_X1 U732 ( .A(G107), .B(KEYINPUT115), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(G9) );
  XOR2_X1 U734 ( .A(G110), .B(n667), .Z(G12) );
  XOR2_X1 U735 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n669) );
  NAND2_X1 U736 ( .A1(n673), .A2(n677), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U738 ( .A(G128), .B(n670), .ZN(G30) );
  XOR2_X1 U739 ( .A(n671), .B(n672), .Z(G45) );
  NAND2_X1 U740 ( .A1(n673), .A2(n675), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(G146), .ZN(G48) );
  NAND2_X1 U742 ( .A1(n678), .A2(n675), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(G113), .ZN(G15) );
  XOR2_X1 U744 ( .A(G116), .B(KEYINPUT117), .Z(n680) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(G18) );
  XNOR2_X1 U747 ( .A(G125), .B(n681), .ZN(n682) );
  XNOR2_X1 U748 ( .A(n682), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n688) );
  AND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n715), .A2(n691), .ZN(n710) );
  XOR2_X1 U754 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n695) );
  NAND2_X1 U755 ( .A1(n348), .A2(n692), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n695), .B(n694), .ZN(n701) );
  XOR2_X1 U757 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n699) );
  NAND2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U759 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U763 ( .A(KEYINPUT51), .B(n706), .Z(n707) );
  NOR2_X1 U764 ( .A1(n714), .A2(n707), .ZN(n708) );
  XNOR2_X1 U765 ( .A(n708), .B(KEYINPUT120), .ZN(n709) );
  NOR2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT52), .ZN(n712) );
  NOR2_X1 U768 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U771 ( .A1(n718), .A2(n480), .ZN(n726) );
  INV_X1 U772 ( .A(n739), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n719), .A2(n757), .ZN(n721) );
  XNOR2_X1 U774 ( .A(KEYINPUT81), .B(KEYINPUT2), .ZN(n720) );
  NAND2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U776 ( .A(KEYINPUT80), .B(n722), .Z(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n727), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U780 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n728), .B(KEYINPUT57), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U783 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n389), .A2(G478), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U786 ( .A1(n738), .A2(n737), .ZN(G63) );
  NOR2_X1 U787 ( .A1(n739), .A2(G953), .ZN(n740) );
  XNOR2_X1 U788 ( .A(n740), .B(KEYINPUT125), .ZN(n745) );
  NAND2_X1 U789 ( .A1(G224), .A2(G953), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n741), .B(KEYINPUT61), .ZN(n742) );
  XNOR2_X1 U791 ( .A(KEYINPUT124), .B(n742), .ZN(n743) );
  NAND2_X1 U792 ( .A1(n743), .A2(G898), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n745), .A2(n744), .ZN(n753) );
  XOR2_X1 U794 ( .A(G101), .B(KEYINPUT127), .Z(n746) );
  XNOR2_X1 U795 ( .A(n747), .B(n746), .ZN(n749) );
  XNOR2_X1 U796 ( .A(n373), .B(n749), .ZN(n750) );
  NOR2_X1 U797 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U798 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U799 ( .A(KEYINPUT126), .B(n754), .ZN(G69) );
  XNOR2_X1 U800 ( .A(n756), .B(n382), .ZN(n760) );
  INV_X1 U801 ( .A(n760), .ZN(n758) );
  XNOR2_X1 U802 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U803 ( .A1(n759), .A2(n480), .ZN(n764) );
  XNOR2_X1 U804 ( .A(G227), .B(n760), .ZN(n761) );
  NAND2_X1 U805 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U806 ( .A1(n762), .A2(G953), .ZN(n763) );
  NAND2_X1 U807 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U808 ( .A(G137), .B(n765), .Z(G39) );
  XOR2_X1 U809 ( .A(n766), .B(G131), .Z(G33) );
  XOR2_X1 U810 ( .A(G134), .B(n767), .Z(G36) );
endmodule

