//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n203), .A2(G50), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT67), .B(G244), .Z(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n215), .A2(G77), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT66), .B(G238), .Z(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n202), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n222), .B(new_n223), .C1(new_n217), .C2(new_n216), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G41), .ZN(new_n243));
  INV_X1    g0043(.A(G45), .ZN(new_n244));
  AOI21_X1  g0044(.A(G1), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(new_n247), .A3(G274), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G226), .A2(G1698), .ZN(new_n249));
  INV_X1    g0049(.A(G232), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n249), .B1(new_n250), .B2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n251), .A2(new_n256), .B1(G33), .B2(G97), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n248), .B1(new_n257), .B2(new_n247), .ZN(new_n258));
  INV_X1    g0058(.A(G238), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n247), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n247), .A2(KEYINPUT69), .A3(new_n261), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT13), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n248), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n250), .A2(G1698), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G226), .B2(G1698), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n247), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n268), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n265), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT69), .B1(new_n247), .B2(new_n261), .ZN(new_n280));
  OAI21_X1  g0080(.A(G238), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n267), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G200), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(new_n211), .A3(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n202), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT12), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n211), .A2(new_n253), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n291));
  INV_X1    g0091(.A(G77), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n211), .A2(G33), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n210), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(KEYINPUT11), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n286), .A2(new_n296), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n211), .A2(G1), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G68), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n288), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT11), .B1(new_n294), .B2(new_n296), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n267), .A2(new_n282), .A3(G190), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n284), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n283), .B2(G169), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n267), .A2(new_n282), .A3(G179), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n258), .A2(new_n266), .A3(KEYINPUT13), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n278), .B1(new_n277), .B2(new_n281), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n308), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n304), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n307), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n219), .A2(G1698), .A3(new_n256), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n256), .A2(G232), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G107), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n318), .B(new_n320), .C1(new_n321), .C2(new_n256), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n276), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n264), .A2(new_n265), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n268), .B1(new_n324), .B2(new_n215), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n298), .A2(G77), .A3(new_n300), .ZN(new_n329));
  INV_X1    g0129(.A(new_n286), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n330), .A2(KEYINPUT73), .A3(G77), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n286), .B2(new_n292), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n296), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n338));
  INV_X1    g0138(.A(G87), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT15), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT15), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G87), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n293), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n335), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n334), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n328), .B(new_n348), .C1(G179), .C2(new_n326), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n347), .B1(new_n326), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n323), .B2(new_n325), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n317), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n256), .A2(G222), .A3(new_n319), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n274), .A2(G77), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT70), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT70), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n356), .A2(new_n357), .A3(new_n361), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n276), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT68), .B(G226), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n268), .B1(new_n324), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n247), .B1(new_n360), .B2(new_n362), .ZN(new_n369));
  INV_X1    g0169(.A(new_n367), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT71), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n371), .A3(G200), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  INV_X1    g0173(.A(G50), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n211), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT72), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n337), .A2(new_n344), .B1(G150), .B2(new_n290), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n335), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n298), .A2(G50), .A3(new_n300), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G50), .B2(new_n330), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT9), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n350), .B1(new_n368), .B2(new_n371), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT10), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n385), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT10), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n372), .A4(new_n383), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n336), .A2(new_n299), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n296), .B(new_n286), .C1(new_n391), .C2(KEYINPUT76), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n391), .A2(KEYINPUT76), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n392), .A2(new_n393), .B1(new_n336), .B2(new_n286), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n289), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT75), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(G58), .A3(G68), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n401), .A3(new_n203), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n395), .B(new_n397), .C1(G20), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n272), .A2(new_n273), .A3(new_n404), .A4(G20), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n272), .B2(new_n273), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n254), .A2(KEYINPUT74), .A3(new_n255), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n211), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n409), .B2(new_n404), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n403), .B1(new_n410), .B2(new_n202), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n254), .A2(new_n211), .A3(new_n255), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n404), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n202), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(G20), .ZN(new_n416));
  INV_X1    g0216(.A(new_n397), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n395), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n411), .A2(new_n296), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(G223), .B(new_n319), .C1(new_n272), .C2(new_n273), .ZN(new_n421));
  OAI211_X1 g0221(.A(G226), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT77), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n276), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n247), .A2(G232), .A3(new_n261), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n248), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(G200), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n247), .B1(new_n426), .B2(new_n427), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n248), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n350), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n394), .B(new_n420), .C1(new_n433), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n420), .A2(new_n394), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n327), .B1(new_n434), .B2(new_n431), .ZN(new_n444));
  INV_X1    g0244(.A(G179), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n435), .A2(new_n445), .A3(new_n437), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n434), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT18), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n429), .A2(new_n432), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n451), .B2(new_n327), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n443), .ZN(new_n454));
  INV_X1    g0254(.A(new_n443), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n434), .A2(new_n431), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n456), .A2(G200), .B1(new_n434), .B2(new_n438), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT17), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n442), .A2(new_n450), .A3(new_n454), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n365), .B1(new_n364), .B2(new_n367), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT71), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n327), .ZN(new_n464));
  INV_X1    g0264(.A(new_n381), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(G179), .C2(new_n463), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n355), .A2(new_n390), .A3(new_n460), .A4(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G250), .A2(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT4), .A2(G244), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(G1698), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n256), .A2(new_n473), .B1(G33), .B2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(G244), .B(new_n319), .C1(new_n272), .C2(new_n273), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n276), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n244), .A2(G1), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G257), .A3(new_n247), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n260), .A2(G45), .ZN(new_n486));
  OR2_X1    g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(new_n481), .ZN(new_n488));
  INV_X1    g0288(.A(G274), .ZN(new_n489));
  AND2_X1   g0289(.A1(G1), .A2(G13), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n246), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n479), .A2(KEYINPUT80), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n247), .B1(new_n474), .B2(new_n477), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n485), .A2(new_n492), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(G200), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G190), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n330), .A2(G97), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n260), .A2(G33), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n298), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT7), .B1(new_n274), .B2(new_n211), .ZN(new_n508));
  OAI21_X1  g0308(.A(G107), .B1(new_n508), .B2(new_n405), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  AND2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n321), .A2(KEYINPUT6), .A3(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n507), .B1(new_n517), .B2(new_n296), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n499), .A2(new_n501), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(G20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n290), .A2(G77), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n321), .B1(new_n413), .B2(new_n414), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n296), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n505), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n502), .B1(new_n525), .B2(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n485), .A2(new_n492), .A3(new_n445), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n496), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n327), .B1(new_n496), .B2(new_n497), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n479), .A2(KEYINPUT81), .A3(new_n493), .A4(new_n445), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n527), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n211), .B1(new_n269), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n512), .A2(new_n339), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n211), .B(G68), .C1(new_n272), .C2(new_n273), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n293), .B2(new_n506), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n296), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT15), .B(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n286), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n343), .A2(KEYINPUT82), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n298), .A2(new_n544), .A3(new_n546), .A4(new_n504), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n259), .A2(new_n319), .ZN(new_n549));
  INV_X1    g0349(.A(G244), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G1698), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n551), .C1(new_n272), .C2(new_n273), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n253), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n247), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G250), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n260), .B2(G45), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n247), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n247), .A2(G274), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n486), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n327), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n491), .A2(new_n480), .B1(new_n247), .B2(new_n558), .ZN(new_n563));
  NOR2_X1   g0363(.A1(G238), .A2(G1698), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n550), .B2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n554), .B1(new_n565), .B2(new_n256), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n563), .B(new_n445), .C1(new_n566), .C2(new_n247), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n548), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n525), .A2(G87), .ZN(new_n569));
  OAI21_X1  g0369(.A(G200), .B1(new_n556), .B2(new_n561), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n540), .A2(new_n296), .B1(new_n286), .B2(new_n542), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n563), .B(G190), .C1(new_n566), .C2(new_n247), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n519), .A2(new_n533), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT83), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n519), .A2(new_n533), .A3(KEYINPUT83), .A4(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n286), .A2(new_n553), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n298), .A2(G116), .A3(new_n504), .ZN(new_n581));
  AOI21_X1  g0381(.A(G20), .B1(G33), .B2(G283), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G33), .B2(new_n506), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n553), .A2(G20), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n296), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n580), .B(new_n581), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n488), .A2(new_n276), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G270), .B1(new_n491), .B2(new_n488), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n592));
  OAI211_X1 g0392(.A(G257), .B(new_n319), .C1(new_n272), .C2(new_n273), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n256), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n276), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n589), .A2(G169), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n591), .A2(G179), .A3(new_n596), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(KEYINPUT21), .B1(new_n589), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n589), .B1(G200), .B2(new_n597), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n350), .B2(new_n597), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n589), .A2(new_n597), .A3(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n579), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT25), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n330), .B2(G107), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n321), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n525), .A2(G107), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n211), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT22), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n256), .A2(new_n616), .A3(new_n211), .A4(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT23), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n211), .B2(G107), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n321), .A2(KEYINPUT23), .A3(G20), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n620), .A2(new_n621), .B1(new_n554), .B2(new_n211), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT24), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT24), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n618), .A2(new_n625), .A3(new_n622), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n613), .B1(new_n627), .B2(new_n296), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n484), .A2(G264), .A3(new_n247), .ZN(new_n629));
  NOR2_X1   g0429(.A1(G250), .A2(G1698), .ZN(new_n630));
  INV_X1    g0430(.A(G257), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(G1698), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n256), .B1(G33), .B2(G294), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n492), .B(new_n629), .C1(new_n633), .C2(new_n247), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n352), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT84), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT84), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n637), .A3(new_n352), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n631), .A2(G1698), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(G250), .B2(G1698), .ZN(new_n640));
  INV_X1    g0440(.A(G294), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n640), .A2(new_n274), .B1(new_n253), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(G264), .A2(new_n590), .B1(new_n642), .B2(new_n276), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n350), .A3(new_n492), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n636), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n628), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n618), .A2(new_n625), .A3(new_n622), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n625), .B1(new_n618), .B2(new_n622), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n296), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n612), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n643), .A2(new_n445), .A3(new_n492), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n634), .A2(new_n327), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT85), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n646), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n646), .B2(new_n655), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n470), .A2(new_n608), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT86), .ZN(G372));
  INV_X1    g0461(.A(new_n470), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n600), .A2(new_n605), .A3(new_n655), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n519), .A2(new_n533), .ZN(new_n664));
  INV_X1    g0464(.A(new_n573), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n562), .B(KEYINPUT87), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n548), .A2(new_n567), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n663), .A2(new_n664), .A3(new_n646), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n533), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n672), .A2(KEYINPUT26), .A3(new_n574), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n532), .A2(new_n530), .A3(new_n531), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n668), .A3(new_n527), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n466), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n386), .A2(new_n389), .A3(KEYINPUT89), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT89), .B1(new_n386), .B2(new_n389), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n453), .A2(new_n443), .A3(new_n444), .A4(new_n448), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n453), .B1(new_n452), .B2(new_n443), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n433), .A2(new_n439), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n689), .A2(new_n441), .A3(new_n443), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT17), .B1(new_n455), .B2(new_n457), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n306), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n314), .A2(new_n311), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n316), .B1(new_n694), .B2(new_n309), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n349), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n688), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n682), .B1(new_n685), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n681), .A2(new_n698), .ZN(G369));
  NAND3_X1  g0499(.A1(new_n260), .A2(new_n211), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(G213), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n589), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n606), .B2(KEYINPUT90), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(KEYINPUT90), .B2(new_n606), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n600), .A2(new_n605), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n706), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n705), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n655), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n657), .B2(new_n658), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n659), .B2(new_n650), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n714), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n655), .A2(new_n705), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n710), .A2(new_n705), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n207), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n536), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n214), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n634), .A2(new_n637), .A3(new_n352), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n637), .B1(new_n634), .B2(new_n352), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n634), .A2(G190), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n650), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n628), .A2(new_n653), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT85), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n646), .A2(new_n655), .A3(new_n656), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n705), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n606), .B1(new_n577), .B2(new_n578), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n556), .A2(new_n561), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n643), .A2(new_n479), .A3(new_n493), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n591), .A2(new_n596), .A3(G179), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n629), .B1(new_n633), .B2(new_n247), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n556), .A3(new_n561), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n599), .A2(new_n749), .A3(KEYINPUT30), .A4(new_n500), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n479), .A2(new_n493), .B1(new_n591), .B2(new_n596), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT91), .B1(new_n556), .B2(new_n561), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT91), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n563), .B(new_n753), .C1(new_n566), .C2(new_n247), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n634), .A2(new_n445), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n751), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n747), .A2(new_n750), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT92), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n758), .A2(KEYINPUT92), .A3(KEYINPUT31), .A4(new_n705), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n758), .A2(new_n705), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n761), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n713), .B1(new_n742), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n680), .A2(new_n715), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n677), .A2(KEYINPUT26), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n672), .A2(new_n678), .A3(new_n574), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n670), .B(KEYINPUT93), .Z(new_n773));
  NAND4_X1  g0573(.A1(new_n669), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(KEYINPUT29), .A3(new_n715), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n767), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n731), .B1(new_n776), .B2(G1), .ZN(G364));
  NOR2_X1   g0577(.A1(new_n285), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n260), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n726), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n714), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(G330), .B1(new_n708), .B2(new_n711), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n285), .A2(new_n253), .A3(KEYINPUT95), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT95), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G13), .B2(G33), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n712), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n210), .B1(G20), .B2(new_n327), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n241), .A2(G45), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n407), .A2(new_n408), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n725), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G45), .C2(new_n214), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n725), .A2(new_n274), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G355), .B1(new_n553), .B2(new_n725), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n794), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n792), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n211), .A2(new_n445), .A3(new_n350), .A4(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n211), .A2(new_n445), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G190), .A2(G200), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n274), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n211), .A2(G179), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n809), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n807), .B(new_n813), .C1(G329), .C2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n808), .A2(G190), .A3(G200), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G326), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n808), .A2(new_n350), .A3(G200), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n814), .A2(G190), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n822), .A2(new_n823), .B1(new_n825), .B2(G303), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n350), .A2(G179), .A3(G200), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n211), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n814), .A2(new_n350), .A3(G200), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n829), .A2(G294), .B1(new_n831), .B2(G283), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n817), .A2(new_n820), .A3(new_n826), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(KEYINPUT96), .B(G159), .Z(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n815), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n836), .A2(KEYINPUT32), .B1(new_n339), .B2(new_n824), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G68), .B2(new_n822), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n256), .B1(new_n811), .B2(new_n292), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G58), .B2(new_n804), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n836), .A2(KEYINPUT32), .B1(G107), .B2(new_n831), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G97), .A2(new_n829), .B1(new_n819), .B2(G50), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n838), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n803), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n781), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n802), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n782), .A2(new_n784), .B1(new_n791), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  NOR2_X1   g0648(.A1(new_n788), .A2(new_n792), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n781), .B1(new_n850), .B2(G77), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n811), .A2(new_n553), .B1(new_n815), .B2(new_n812), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n274), .B1(new_n805), .B2(new_n641), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n828), .A2(new_n506), .B1(new_n821), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G303), .A2(new_n819), .B1(new_n825), .B2(G107), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n339), .C2(new_n830), .ZN(new_n858));
  INV_X1    g0658(.A(new_n834), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(new_n810), .B1(new_n804), .B2(G143), .ZN(new_n860));
  INV_X1    g0660(.A(G137), .ZN(new_n861));
  INV_X1    g0661(.A(G150), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n861), .B2(new_n818), .C1(new_n862), .C2(new_n821), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT34), .Z(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n797), .B1(new_n865), .B2(new_n815), .C1(new_n201), .C2(new_n828), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT97), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n374), .A2(new_n824), .B1(new_n830), .B2(new_n202), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n858), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n851), .B1(new_n871), .B2(new_n792), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT98), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n349), .A2(new_n705), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n351), .A2(new_n353), .B1(new_n347), .B2(new_n715), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n349), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n873), .B1(new_n788), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n768), .A2(new_n877), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n874), .A2(new_n876), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n715), .B(new_n880), .C1(new_n671), .C2(new_n679), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n767), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n781), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n767), .A3(new_n881), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  NOR2_X1   g0686(.A1(new_n778), .A2(new_n260), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n409), .A2(new_n404), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n414), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G68), .ZN(new_n891));
  INV_X1    g0691(.A(new_n418), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT16), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n411), .A2(new_n296), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n394), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n703), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n692), .B2(new_n688), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n452), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n897), .A3(new_n440), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n440), .A2(new_n449), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT37), .B1(new_n443), .B2(new_n896), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n900), .A2(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n888), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT99), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n901), .A2(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n897), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n459), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT99), .B(new_n888), .C1(new_n898), .C2(new_n903), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT101), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n765), .A2(new_n759), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n740), .B2(new_n741), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n316), .A2(new_n705), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n695), .A2(new_n306), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n695), .B2(new_n306), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n880), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n914), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n765), .A2(new_n759), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n608), .B2(new_n717), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n316), .B(new_n705), .C1(new_n315), .C2(new_n307), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n695), .A2(new_n306), .A3(new_n917), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n877), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(KEYINPUT101), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n912), .A2(new_n913), .A3(new_n921), .A4(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT102), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(KEYINPUT102), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n443), .A2(new_n896), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT100), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n440), .A2(new_n449), .A3(new_n935), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n935), .B1(new_n692), .B2(new_n688), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n888), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n929), .B1(new_n943), .B2(new_n911), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n916), .A2(new_n920), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n934), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n662), .A2(new_n923), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(G330), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n947), .B2(new_n948), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT39), .B1(new_n943), .B2(new_n911), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n912), .A2(new_n913), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n315), .A2(new_n316), .A3(new_n715), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n688), .A2(new_n896), .ZN(new_n959));
  INV_X1    g0759(.A(new_n954), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n918), .A2(new_n919), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n881), .B2(new_n874), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n770), .B(new_n775), .C1(new_n468), .C2(new_n469), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n698), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n887), .B1(new_n952), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n952), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(new_n553), .A4(new_n213), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT36), .Z(new_n973));
  INV_X1    g0773(.A(new_n214), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n974), .A2(G77), .A3(new_n401), .A4(new_n399), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n374), .A2(G68), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(G1), .A3(new_n285), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n969), .A2(new_n973), .A3(new_n978), .ZN(G367));
  AND2_X1   g0779(.A1(new_n718), .A2(new_n722), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n664), .B1(new_n518), .B2(new_n715), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n675), .A2(new_n527), .A3(new_n676), .A4(new_n705), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n984), .A2(KEYINPUT42), .B1(new_n672), .B2(new_n715), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n723), .A2(new_n721), .ZN(new_n986));
  INV_X1    g0786(.A(new_n983), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(KEYINPUT42), .B2(new_n721), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n670), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n569), .A2(new_n571), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n715), .ZN(new_n992));
  MUX2_X1   g0792(.A(new_n668), .B(new_n990), .S(new_n992), .Z(new_n993));
  AOI22_X1  g0793(.A1(new_n985), .A2(new_n989), .B1(KEYINPUT43), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n719), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n983), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n996), .B(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n726), .B(KEYINPUT41), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n986), .A2(new_n987), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n983), .B1(new_n723), .B2(new_n721), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT103), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n1006), .A3(new_n997), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n776), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n718), .A2(new_n716), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n710), .B2(new_n705), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT104), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n714), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1010), .B(new_n1011), .C1(new_n713), .C2(new_n712), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n723), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n980), .A3(new_n1014), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1008), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1002), .A2(new_n719), .A3(new_n1004), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1007), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1000), .B1(new_n1021), .B2(new_n776), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n999), .B1(new_n1022), .B2(new_n780), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n793), .B1(new_n207), .B2(new_n542), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n234), .A2(new_n725), .A3(new_n797), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n781), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n830), .A2(new_n506), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n641), .A2(new_n821), .B1(new_n818), .B2(new_n812), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n829), .A2(G107), .B1(G283), .B2(new_n810), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(KEYINPUT105), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT105), .B2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n816), .B1(new_n804), .B2(G303), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n797), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n824), .B2(new_n553), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n825), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n859), .A2(new_n822), .B1(new_n819), .B2(G143), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n829), .A2(G68), .B1(new_n825), .B2(G58), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n804), .A2(G150), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G50), .A2(new_n810), .B1(new_n816), .B2(G137), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n830), .A2(new_n292), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n274), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT106), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1031), .A2(new_n1037), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT47), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1026), .B1(new_n1047), .B2(new_n792), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n790), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(new_n993), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1023), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT107), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT107), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1023), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1054), .ZN(G387));
  NOR2_X1   g0855(.A1(new_n1018), .A2(new_n727), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n776), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n728), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1059), .A2(new_n800), .B1(new_n321), .B2(new_n725), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT108), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n231), .A2(new_n244), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n337), .A2(new_n374), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n728), .B(new_n244), .C1(new_n202), .C2(new_n292), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n798), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n845), .B1(new_n1067), .B2(new_n793), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1009), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n1049), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n811), .A2(new_n202), .B1(new_n336), .B2(new_n821), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT109), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n824), .A2(new_n292), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1027), .B(new_n1073), .C1(G159), .C2(new_n819), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n544), .A2(new_n546), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n829), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n805), .A2(new_n374), .B1(new_n815), .B2(new_n862), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n1033), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1072), .A2(new_n1074), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n829), .A2(G283), .B1(new_n825), .B2(G294), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n812), .A2(new_n821), .B1(new_n818), .B2(new_n806), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT110), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(KEYINPUT110), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G303), .A2(new_n810), .B1(new_n804), .B2(G317), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT111), .Z(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1091), .B(new_n1092), .Z(new_n1093));
  INV_X1    g0893(.A(KEYINPUT113), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n797), .B1(G326), .B2(new_n816), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n553), .B2(new_n830), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT114), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1080), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1070), .B1(new_n1100), .B2(new_n792), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1057), .B2(new_n780), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1058), .A2(new_n1102), .ZN(G393));
  INV_X1    g0903(.A(new_n1018), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1005), .A2(new_n997), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1020), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n727), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1021), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n780), .A3(new_n1020), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT118), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n794), .B1(G97), .B2(new_n725), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n238), .A2(new_n798), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n845), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n819), .A2(G150), .B1(new_n804), .B2(G159), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n828), .A2(new_n292), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n202), .A2(new_n824), .B1(new_n830), .B2(new_n339), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(G50), .C2(new_n822), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n337), .A2(new_n810), .B1(new_n816), .B2(G143), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n797), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT116), .Z(new_n1122));
  AOI22_X1  g0922(.A1(new_n819), .A2(G317), .B1(new_n804), .B2(G311), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT52), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n274), .B1(new_n806), .B2(new_n815), .C1(new_n811), .C2(new_n641), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n821), .A2(new_n594), .B1(new_n830), .B2(new_n321), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n828), .A2(new_n553), .B1(new_n824), .B2(new_n854), .ZN(new_n1127));
  OR3_X1    g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1122), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1113), .B1(new_n1049), .B2(new_n983), .C1(new_n1130), .C2(new_n803), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1109), .A2(new_n1110), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1110), .B1(new_n1109), .B2(new_n1131), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1108), .B1(new_n1132), .B2(new_n1133), .ZN(G390));
  INV_X1    g0934(.A(KEYINPUT39), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n912), .B2(new_n913), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1136), .A2(new_n953), .B1(new_n957), .B2(new_n962), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n957), .B1(new_n943), .B2(new_n911), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n774), .A2(new_n715), .A3(new_n876), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1139), .A2(new_n874), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1140), .B2(new_n961), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n961), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n767), .A2(new_n880), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1137), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n923), .A2(G330), .A3(new_n926), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n916), .A2(new_n713), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1142), .B1(new_n1148), .B2(new_n880), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n881), .A2(new_n874), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1142), .B1(new_n767), .B2(new_n880), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1145), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(KEYINPUT119), .B(new_n1151), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1150), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(G330), .B(new_n923), .C1(new_n468), .C2(new_n469), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n965), .A2(new_n1159), .A3(new_n698), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1144), .A2(new_n1146), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n962), .A2(new_n957), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1141), .B1(new_n955), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1153), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1157), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n713), .B(new_n877), .C1(new_n742), .C2(new_n766), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1145), .B1(new_n1167), .B2(new_n1142), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT119), .B1(new_n1168), .B2(new_n1151), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1165), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n965), .A2(new_n1159), .A3(new_n698), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1137), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1164), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1161), .A2(new_n1173), .A3(new_n726), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n811), .A2(new_n1175), .B1(new_n805), .B2(new_n865), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n256), .B1(new_n815), .B2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n821), .A2(new_n861), .B1(new_n830), .B2(new_n374), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n828), .A2(new_n396), .B1(new_n818), .B2(new_n1180), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n824), .A2(new_n862), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT53), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n811), .A2(new_n506), .B1(new_n815), .B2(new_n641), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n274), .B1(new_n805), .B2(new_n553), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n202), .A2(new_n830), .B1(new_n824), .B2(new_n339), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n818), .A2(new_n854), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1189), .B(new_n1117), .C1(G107), .C2(new_n822), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1182), .A2(new_n1184), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n781), .B1(new_n337), .B2(new_n850), .C1(new_n1191), .C2(new_n803), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n955), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n788), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n780), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1174), .A2(new_n1196), .ZN(G378));
  OAI21_X1  g0997(.A(new_n466), .B1(new_n683), .B2(new_n684), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n381), .A2(new_n703), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n466), .B1(new_n381), .B2(new_n703), .C1(new_n683), .C2(new_n684), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n713), .B1(new_n944), .B2(new_n945), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n934), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n928), .A2(KEYINPUT102), .A3(new_n929), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT102), .B1(new_n928), .B2(new_n929), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1206), .B(new_n1205), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n964), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1173), .A2(new_n1171), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1205), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(new_n958), .A3(new_n963), .A4(new_n1210), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1212), .A2(new_n1213), .A3(KEYINPUT57), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n726), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT120), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n958), .B2(new_n963), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1216), .A2(new_n1221), .A3(new_n1210), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1213), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1205), .A2(new_n788), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1033), .A2(new_n243), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G283), .A2(new_n816), .B1(new_n804), .B2(G107), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n202), .B2(new_n828), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(new_n1076), .C2(new_n810), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n506), .A2(new_n821), .B1(new_n818), .B2(new_n553), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1073), .B(new_n1233), .C1(G58), .C2(new_n831), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G50), .B1(new_n253), .B2(new_n243), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1235), .A2(KEYINPUT58), .B1(new_n1229), .B2(new_n1236), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1177), .A2(new_n818), .B1(new_n821), .B2(new_n865), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G137), .A2(new_n810), .B1(new_n804), .B2(G128), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n824), .B2(new_n1175), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G150), .C2(new_n829), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n859), .A2(new_n831), .ZN(new_n1244));
  AOI211_X1 g1044(.A(G33), .B(G41), .C1(new_n816), .C2(G124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1237), .B1(KEYINPUT58), .B2(new_n1235), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n792), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n849), .A2(new_n374), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1228), .A2(new_n781), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1225), .B2(new_n780), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1227), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1000), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT121), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT122), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1158), .B2(new_n779), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1170), .A2(KEYINPUT122), .A3(new_n780), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n818), .A2(new_n641), .B1(new_n824), .B2(new_n506), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1043), .B(new_n1264), .C1(G116), .C2(new_n822), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n256), .B1(new_n816), .B2(G303), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G107), .A2(new_n810), .B1(new_n804), .B2(G283), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1077), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n805), .A2(new_n861), .B1(new_n815), .B2(new_n1180), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(G150), .B2(new_n810), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G132), .A2(new_n819), .B1(new_n825), .B2(G159), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1175), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G50), .A2(new_n829), .B1(new_n822), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1033), .B1(G58), .B2(new_n831), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n803), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n845), .B(new_n1276), .C1(new_n202), .C2(new_n849), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1142), .B2(new_n789), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1262), .A2(new_n1263), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1260), .A2(new_n1280), .ZN(G381));
  NAND3_X1  g1081(.A1(new_n1058), .A2(new_n847), .A3(new_n1102), .ZN(new_n1282));
  OR4_X1    g1082(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT123), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G378), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1174), .A2(KEYINPUT123), .A3(new_n1196), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G387), .A2(G375), .A3(new_n1283), .A4(new_n1287), .ZN(G407));
  INV_X1    g1088(.A(new_n1286), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT123), .B1(new_n1174), .B2(new_n1196), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1254), .A2(new_n704), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  NAND2_X1  g1093(.A1(new_n1256), .A2(new_n726), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1257), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1294), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OR3_X1    g1099(.A1(new_n1299), .A2(new_n885), .A3(new_n1279), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n885), .B1(new_n1299), .B2(new_n1279), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n704), .A2(G213), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1216), .A2(new_n1221), .A3(new_n1210), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1221), .B1(new_n1216), .B2(new_n1210), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1258), .B(new_n1213), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1212), .A2(new_n780), .A3(new_n1217), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1251), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G378), .B(new_n1253), .C1(new_n1219), .C2(new_n1226), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1291), .B2(new_n1309), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1303), .B(new_n1304), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1304), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n704), .A2(G213), .A3(G2897), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1300), .A2(new_n1301), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1307), .A2(new_n1251), .A3(new_n1308), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT124), .B1(new_n1324), .B2(new_n1287), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1316), .A2(new_n1322), .A3(new_n1323), .A4(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(G390), .A2(new_n1023), .A3(new_n1050), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(G390), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1051), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(G390), .A2(new_n1023), .A3(KEYINPUT127), .A4(new_n1050), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1332), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G393), .A2(G396), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1282), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1338), .B(KEYINPUT126), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1052), .A2(new_n1054), .A3(new_n1333), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1330), .A2(new_n1338), .ZN(new_n1341));
  AOI22_X1  g1141(.A1(new_n1336), .A2(new_n1339), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1329), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1342), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT61), .B1(new_n1317), .B2(new_n1321), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1315), .A2(new_n1346), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1344), .A2(new_n1345), .A3(new_n1347), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1343), .A2(new_n1349), .ZN(G405));
  OAI21_X1  g1150(.A(new_n1312), .B1(new_n1254), .B2(new_n1287), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1303), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1302), .B(new_n1312), .C1(new_n1254), .C2(new_n1287), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1352), .A2(new_n1342), .A3(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1342), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(G402));
endmodule


