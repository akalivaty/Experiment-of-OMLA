

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(KEYINPUT28), .ZN(n636) );
  XNOR2_X1 U550 ( .A(n596), .B(KEYINPUT79), .ZN(n512) );
  OR2_X1 U551 ( .A1(n695), .A2(n694), .ZN(n513) );
  NOR2_X1 U552 ( .A1(n725), .A2(n724), .ZN(n514) );
  BUF_X1 U553 ( .A(n628), .Z(n643) );
  NOR2_X1 U554 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U555 ( .A1(n546), .A2(n545), .ZN(n772) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n520), .ZN(n873) );
  NOR2_X1 U557 ( .A1(G651), .A2(n546), .ZN(n769) );
  NOR2_X1 U558 ( .A1(n535), .A2(n534), .ZN(G160) );
  XNOR2_X1 U559 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n516) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XNOR2_X1 U561 ( .A(n516), .B(n515), .ZN(n876) );
  NAND2_X1 U562 ( .A1(G138), .A2(n876), .ZN(n518) );
  INV_X1 U563 ( .A(G2104), .ZN(n519) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n519), .ZN(n877) );
  NAND2_X1 U565 ( .A1(G102), .A2(n877), .ZN(n517) );
  NAND2_X1 U566 ( .A1(n518), .A2(n517), .ZN(n524) );
  INV_X1 U567 ( .A(G2105), .ZN(n520) );
  NOR2_X1 U568 ( .A1(n519), .A2(n520), .ZN(n872) );
  NAND2_X1 U569 ( .A1(G114), .A2(n872), .ZN(n522) );
  NAND2_X1 U570 ( .A1(G126), .A2(n873), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U573 ( .A1(G137), .A2(n876), .ZN(n526) );
  NAND2_X1 U574 ( .A1(G113), .A2(n872), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U576 ( .A(KEYINPUT68), .B(n527), .ZN(n535) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(KEYINPUT23), .Z(n529) );
  NAND2_X1 U578 ( .A1(G101), .A2(n877), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n529), .B(n528), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n873), .A2(G125), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT64), .B(n530), .Z(n531) );
  NOR2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT66), .B(n533), .Z(n534) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n546) );
  NAND2_X1 U585 ( .A1(G49), .A2(n769), .ZN(n536) );
  XNOR2_X1 U586 ( .A(n536), .B(KEYINPUT84), .ZN(n543) );
  INV_X1 U587 ( .A(G651), .ZN(n545) );
  NOR2_X1 U588 ( .A1(G543), .A2(n545), .ZN(n538) );
  XNOR2_X1 U589 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n538), .B(n537), .ZN(n768) );
  NAND2_X1 U591 ( .A1(G87), .A2(n546), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G74), .A2(G651), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U594 ( .A1(n768), .A2(n541), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(G288) );
  NAND2_X1 U596 ( .A1(G65), .A2(n768), .ZN(n544) );
  XOR2_X1 U597 ( .A(KEYINPUT72), .B(n544), .Z(n551) );
  NAND2_X1 U598 ( .A1(G78), .A2(n772), .ZN(n548) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n773) );
  NAND2_X1 U600 ( .A1(G91), .A2(n773), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U602 ( .A(KEYINPUT71), .B(n549), .Z(n550) );
  NOR2_X1 U603 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n769), .A2(G53), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U606 ( .A1(n769), .A2(G52), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n768), .A2(G64), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n561) );
  NAND2_X1 U609 ( .A1(n772), .A2(G77), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n556), .B(KEYINPUT70), .ZN(n558) );
  NAND2_X1 U611 ( .A1(G90), .A2(n773), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U614 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n773), .A2(G89), .ZN(n562) );
  XNOR2_X1 U616 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U617 ( .A1(G76), .A2(n772), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U619 ( .A(KEYINPUT5), .B(n565), .ZN(n571) );
  NAND2_X1 U620 ( .A1(n769), .A2(G51), .ZN(n566) );
  XOR2_X1 U621 ( .A(KEYINPUT81), .B(n566), .Z(n568) );
  NAND2_X1 U622 ( .A1(n768), .A2(G63), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U625 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U626 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G75), .A2(n772), .ZN(n574) );
  NAND2_X1 U629 ( .A1(G88), .A2(n773), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U631 ( .A1(G62), .A2(n768), .ZN(n575) );
  XNOR2_X1 U632 ( .A(KEYINPUT85), .B(n575), .ZN(n576) );
  NOR2_X1 U633 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n769), .A2(G50), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G86), .A2(n773), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G61), .A2(n768), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n772), .A2(G73), .ZN(n582) );
  XOR2_X1 U640 ( .A(KEYINPUT2), .B(n582), .Z(n583) );
  NOR2_X1 U641 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n769), .A2(G48), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U644 ( .A1(G72), .A2(n772), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G85), .A2(n773), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U647 ( .A1(G60), .A2(n768), .ZN(n590) );
  NAND2_X1 U648 ( .A1(G47), .A2(n769), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U650 ( .A1(n592), .A2(n591), .ZN(G290) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n698) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n697) );
  INV_X1 U653 ( .A(n697), .ZN(n614) );
  NAND2_X1 U654 ( .A1(n698), .A2(n614), .ZN(n659) );
  NAND2_X1 U655 ( .A1(G8), .A2(n659), .ZN(n693) );
  NOR2_X1 U656 ( .A1(G1976), .A2(G288), .ZN(n677) );
  NAND2_X1 U657 ( .A1(n677), .A2(KEYINPUT33), .ZN(n593) );
  NOR2_X1 U658 ( .A1(n693), .A2(n593), .ZN(n683) );
  NAND2_X1 U659 ( .A1(G79), .A2(n772), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G54), .A2(n769), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G66), .A2(n768), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n512), .A2(n597), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n773), .A2(G92), .ZN(n598) );
  XOR2_X1 U665 ( .A(KEYINPUT78), .B(n598), .Z(n599) );
  NOR2_X1 U666 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X2 U667 ( .A(KEYINPUT15), .B(n601), .Z(n1001) );
  NAND2_X1 U668 ( .A1(G68), .A2(n772), .ZN(n605) );
  XOR2_X1 U669 ( .A(KEYINPUT12), .B(KEYINPUT75), .Z(n603) );
  NAND2_X1 U670 ( .A1(G81), .A2(n773), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n608) );
  XNOR2_X1 U673 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n606), .B(KEYINPUT13), .ZN(n607) );
  XNOR2_X1 U675 ( .A(n608), .B(n607), .ZN(n611) );
  NAND2_X1 U676 ( .A1(n768), .A2(G56), .ZN(n609) );
  XOR2_X1 U677 ( .A(KEYINPUT14), .B(n609), .Z(n610) );
  NOR2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n769), .A2(G43), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n998) );
  AND2_X1 U681 ( .A1(n698), .A2(n614), .ZN(n641) );
  AND2_X1 U682 ( .A1(n641), .A2(G1996), .ZN(n615) );
  XOR2_X1 U683 ( .A(n615), .B(KEYINPUT26), .Z(n617) );
  NAND2_X1 U684 ( .A1(n659), .A2(G1341), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n621) );
  NOR2_X1 U686 ( .A1(n998), .A2(n621), .ZN(n618) );
  OR2_X1 U687 ( .A1(n1001), .A2(n618), .ZN(n627) );
  INV_X1 U688 ( .A(n1001), .ZN(n619) );
  OR2_X1 U689 ( .A1(n619), .A2(n998), .ZN(n620) );
  OR2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n625) );
  XNOR2_X1 U691 ( .A(KEYINPUT95), .B(n659), .ZN(n628) );
  NAND2_X1 U692 ( .A1(G2067), .A2(n643), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G1348), .A2(n659), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n634) );
  INV_X1 U697 ( .A(G299), .ZN(n995) );
  NAND2_X1 U698 ( .A1(n628), .A2(G2072), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n629), .B(KEYINPUT27), .ZN(n632) );
  INV_X1 U700 ( .A(G1956), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n630), .A2(n643), .ZN(n631) );
  NOR2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U703 ( .A1(n995), .A2(n635), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n635), .A2(n995), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U707 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT29), .B(n640), .Z(n647) );
  NOR2_X1 U709 ( .A1(n641), .A2(G1961), .ZN(n642) );
  XOR2_X1 U710 ( .A(KEYINPUT94), .B(n642), .Z(n645) );
  XNOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .ZN(n960) );
  NAND2_X1 U712 ( .A1(n643), .A2(n960), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n652) );
  NAND2_X1 U714 ( .A1(n652), .A2(G171), .ZN(n646) );
  NAND2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n658) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n693), .ZN(n671) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n659), .ZN(n668) );
  NOR2_X1 U718 ( .A1(n671), .A2(n668), .ZN(n648) );
  NAND2_X1 U719 ( .A1(G8), .A2(n648), .ZN(n650) );
  XNOR2_X1 U720 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X1 U722 ( .A1(G168), .A2(n651), .ZN(n655) );
  NOR2_X1 U723 ( .A1(G171), .A2(n652), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT97), .B(n653), .Z(n654) );
  XOR2_X1 U725 ( .A(KEYINPUT31), .B(n656), .Z(n657) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n669) );
  NAND2_X1 U727 ( .A1(n669), .A2(G286), .ZN(n665) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n693), .ZN(n661) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n659), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n662), .A2(G303), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(KEYINPUT98), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n666), .A2(G8), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT32), .ZN(n675) );
  NAND2_X1 U736 ( .A1(G8), .A2(n668), .ZN(n673) );
  INV_X1 U737 ( .A(n669), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n687) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n988) );
  NAND2_X1 U743 ( .A1(n687), .A2(n988), .ZN(n680) );
  INV_X1 U744 ( .A(n693), .ZN(n678) );
  NAND2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n987) );
  AND2_X1 U746 ( .A1(n678), .A2(n987), .ZN(n679) );
  AND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n681), .A2(KEYINPUT33), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U750 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U751 ( .A1(n684), .A2(n983), .ZN(n690) );
  NOR2_X1 U752 ( .A1(G2090), .A2(G303), .ZN(n685) );
  NAND2_X1 U753 ( .A1(G8), .A2(n685), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n688), .A2(n693), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n695) );
  NOR2_X1 U757 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U758 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT91), .B(G1986), .Z(n696) );
  XNOR2_X1 U761 ( .A(G290), .B(n696), .ZN(n1003) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n737) );
  AND2_X1 U763 ( .A1(n1003), .A2(n737), .ZN(n725) );
  NAND2_X1 U764 ( .A1(G117), .A2(n872), .ZN(n700) );
  NAND2_X1 U765 ( .A1(G129), .A2(n873), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n877), .A2(G105), .ZN(n701) );
  XOR2_X1 U768 ( .A(KEYINPUT38), .B(n701), .Z(n702) );
  NOR2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U770 ( .A(KEYINPUT93), .B(n704), .Z(n706) );
  NAND2_X1 U771 ( .A1(n876), .A2(G141), .ZN(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n887) );
  AND2_X1 U773 ( .A1(n887), .A2(G1996), .ZN(n928) );
  NAND2_X1 U774 ( .A1(G131), .A2(n876), .ZN(n708) );
  NAND2_X1 U775 ( .A1(G107), .A2(n872), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U777 ( .A1(G95), .A2(n877), .ZN(n710) );
  NAND2_X1 U778 ( .A1(G119), .A2(n873), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n859) );
  INV_X1 U781 ( .A(G1991), .ZN(n962) );
  NOR2_X1 U782 ( .A1(n859), .A2(n962), .ZN(n926) );
  OR2_X1 U783 ( .A1(n928), .A2(n926), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n737), .A2(n713), .ZN(n726) );
  XNOR2_X1 U785 ( .A(G2067), .B(KEYINPUT37), .ZN(n734) );
  NAND2_X1 U786 ( .A1(G116), .A2(n872), .ZN(n715) );
  NAND2_X1 U787 ( .A1(G128), .A2(n873), .ZN(n714) );
  NAND2_X1 U788 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U789 ( .A(n716), .B(KEYINPUT35), .ZN(n721) );
  NAND2_X1 U790 ( .A1(G140), .A2(n876), .ZN(n718) );
  NAND2_X1 U791 ( .A1(G104), .A2(n877), .ZN(n717) );
  NAND2_X1 U792 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U793 ( .A(KEYINPUT34), .B(n719), .Z(n720) );
  NAND2_X1 U794 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U795 ( .A(n722), .B(KEYINPUT36), .Z(n886) );
  OR2_X1 U796 ( .A1(n734), .A2(n886), .ZN(n723) );
  XOR2_X1 U797 ( .A(KEYINPUT92), .B(n723), .Z(n949) );
  NAND2_X1 U798 ( .A1(n737), .A2(n949), .ZN(n732) );
  NAND2_X1 U799 ( .A1(n726), .A2(n732), .ZN(n724) );
  NAND2_X1 U800 ( .A1(n513), .A2(n514), .ZN(n740) );
  NOR2_X1 U801 ( .A1(G1996), .A2(n887), .ZN(n942) );
  INV_X1 U802 ( .A(n726), .ZN(n729) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n727) );
  AND2_X1 U804 ( .A1(n962), .A2(n859), .ZN(n927) );
  NOR2_X1 U805 ( .A1(n727), .A2(n927), .ZN(n728) );
  NOR2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U807 ( .A1(n942), .A2(n730), .ZN(n731) );
  XNOR2_X1 U808 ( .A(n731), .B(KEYINPUT39), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n886), .A2(n734), .ZN(n940) );
  NAND2_X1 U811 ( .A1(n735), .A2(n940), .ZN(n736) );
  NAND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U813 ( .A(KEYINPUT99), .B(n738), .Z(n739) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U815 ( .A(n741), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U816 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U817 ( .A(G108), .ZN(G238) );
  INV_X1 U818 ( .A(G120), .ZN(G236) );
  INV_X1 U819 ( .A(G69), .ZN(G235) );
  INV_X1 U820 ( .A(G132), .ZN(G219) );
  NAND2_X1 U821 ( .A1(G7), .A2(G661), .ZN(n742) );
  XNOR2_X1 U822 ( .A(n742), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U823 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n744) );
  INV_X1 U824 ( .A(G223), .ZN(n817) );
  NAND2_X1 U825 ( .A1(G567), .A2(n817), .ZN(n743) );
  XNOR2_X1 U826 ( .A(n744), .B(n743), .ZN(G234) );
  INV_X1 U827 ( .A(G860), .ZN(n767) );
  OR2_X1 U828 ( .A1(n998), .A2(n767), .ZN(G153) );
  INV_X1 U829 ( .A(G171), .ZN(G301) );
  OR2_X1 U830 ( .A1(n1001), .A2(G868), .ZN(n745) );
  XNOR2_X1 U831 ( .A(n745), .B(KEYINPUT80), .ZN(n747) );
  NAND2_X1 U832 ( .A1(G868), .A2(G301), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(G284) );
  XOR2_X1 U834 ( .A(KEYINPUT82), .B(G868), .Z(n748) );
  NOR2_X1 U835 ( .A1(G286), .A2(n748), .ZN(n751) );
  NOR2_X1 U836 ( .A1(G868), .A2(G299), .ZN(n749) );
  XOR2_X1 U837 ( .A(KEYINPUT83), .B(n749), .Z(n750) );
  NOR2_X1 U838 ( .A1(n751), .A2(n750), .ZN(G297) );
  NAND2_X1 U839 ( .A1(n767), .A2(G559), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n752), .A2(n1001), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n753), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U842 ( .A1(G868), .A2(n998), .ZN(n756) );
  NAND2_X1 U843 ( .A1(G868), .A2(n1001), .ZN(n754) );
  NOR2_X1 U844 ( .A1(G559), .A2(n754), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(G282) );
  NAND2_X1 U846 ( .A1(G123), .A2(n873), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n757), .B(KEYINPUT18), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n872), .A2(G111), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U850 ( .A1(G135), .A2(n876), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G99), .A2(n877), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n925) );
  XNOR2_X1 U854 ( .A(n925), .B(G2096), .ZN(n765) );
  INV_X1 U855 ( .A(G2100), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(G156) );
  NAND2_X1 U857 ( .A1(G559), .A2(n1001), .ZN(n766) );
  XOR2_X1 U858 ( .A(n998), .B(n766), .Z(n784) );
  NAND2_X1 U859 ( .A1(n767), .A2(n784), .ZN(n778) );
  NAND2_X1 U860 ( .A1(G67), .A2(n768), .ZN(n771) );
  NAND2_X1 U861 ( .A1(G55), .A2(n769), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G80), .A2(n772), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G93), .A2(n773), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n786) );
  XOR2_X1 U867 ( .A(n778), .B(n786), .Z(G145) );
  XNOR2_X1 U868 ( .A(KEYINPUT19), .B(G288), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n995), .B(G303), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(G305), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n786), .B(n780), .ZN(n781) );
  XNOR2_X1 U872 ( .A(n781), .B(G290), .ZN(n782) );
  XNOR2_X1 U873 ( .A(n783), .B(n782), .ZN(n826) );
  XNOR2_X1 U874 ( .A(n784), .B(n826), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n785), .A2(G868), .ZN(n788) );
  OR2_X1 U876 ( .A1(G868), .A2(n786), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(G295) );
  NAND2_X1 U878 ( .A1(G2078), .A2(G2084), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT20), .B(n789), .Z(n790) );
  NAND2_X1 U880 ( .A1(G2090), .A2(n790), .ZN(n791) );
  XNOR2_X1 U881 ( .A(KEYINPUT21), .B(n791), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n792), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U883 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U884 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U885 ( .A1(G219), .A2(G220), .ZN(n793) );
  XOR2_X1 U886 ( .A(KEYINPUT22), .B(n793), .Z(n794) );
  NOR2_X1 U887 ( .A1(G218), .A2(n794), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G96), .A2(n795), .ZN(n822) );
  NAND2_X1 U889 ( .A1(G2106), .A2(n822), .ZN(n801) );
  NOR2_X1 U890 ( .A1(G235), .A2(G236), .ZN(n796) );
  XNOR2_X1 U891 ( .A(KEYINPUT86), .B(n796), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n797), .A2(G57), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n798), .A2(G238), .ZN(n799) );
  XNOR2_X1 U894 ( .A(n799), .B(KEYINPUT87), .ZN(n823) );
  NAND2_X1 U895 ( .A1(G567), .A2(n823), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U897 ( .A(KEYINPUT88), .B(n802), .Z(G319) );
  NAND2_X1 U898 ( .A1(G661), .A2(G483), .ZN(n803) );
  XNOR2_X1 U899 ( .A(n803), .B(KEYINPUT89), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n804), .A2(G319), .ZN(n805) );
  XOR2_X1 U901 ( .A(KEYINPUT90), .B(n805), .Z(n821) );
  NAND2_X1 U902 ( .A1(G36), .A2(n821), .ZN(G176) );
  XNOR2_X1 U903 ( .A(G2427), .B(G2451), .ZN(n815) );
  XOR2_X1 U904 ( .A(G2430), .B(G2443), .Z(n807) );
  XNOR2_X1 U905 ( .A(KEYINPUT101), .B(G2435), .ZN(n806) );
  XNOR2_X1 U906 ( .A(n807), .B(n806), .ZN(n811) );
  XOR2_X1 U907 ( .A(G2438), .B(G2454), .Z(n809) );
  XNOR2_X1 U908 ( .A(G1341), .B(G1348), .ZN(n808) );
  XNOR2_X1 U909 ( .A(n809), .B(n808), .ZN(n810) );
  XOR2_X1 U910 ( .A(n811), .B(n810), .Z(n813) );
  XNOR2_X1 U911 ( .A(KEYINPUT100), .B(G2446), .ZN(n812) );
  XNOR2_X1 U912 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U913 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n816), .A2(G14), .ZN(n891) );
  XOR2_X1 U915 ( .A(KEYINPUT102), .B(n891), .Z(G401) );
  NAND2_X1 U916 ( .A1(n817), .A2(G2106), .ZN(n818) );
  XOR2_X1 U917 ( .A(KEYINPUT103), .B(n818), .Z(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U919 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U921 ( .A1(n821), .A2(n820), .ZN(G188) );
  NOR2_X1 U922 ( .A1(n823), .A2(n822), .ZN(G325) );
  XOR2_X1 U923 ( .A(KEYINPUT104), .B(G325), .Z(G261) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G57), .ZN(G237) );
  INV_X1 U927 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U928 ( .A(n998), .B(G286), .ZN(n825) );
  XNOR2_X1 U929 ( .A(G171), .B(n1001), .ZN(n824) );
  XNOR2_X1 U930 ( .A(n825), .B(n824), .ZN(n827) );
  XNOR2_X1 U931 ( .A(n827), .B(n826), .ZN(n828) );
  NOR2_X1 U932 ( .A1(G37), .A2(n828), .ZN(G397) );
  XNOR2_X1 U933 ( .A(G1991), .B(G2474), .ZN(n838) );
  XOR2_X1 U934 ( .A(G1986), .B(G1981), .Z(n830) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1961), .ZN(n829) );
  XNOR2_X1 U936 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U937 ( .A(G1976), .B(G1971), .Z(n832) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1956), .ZN(n831) );
  XNOR2_X1 U939 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U940 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U941 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n835) );
  XNOR2_X1 U942 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U944 ( .A(G2678), .B(G2090), .Z(n840) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2084), .ZN(n839) );
  XNOR2_X1 U946 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U947 ( .A(n841), .B(G2100), .Z(n843) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2072), .ZN(n842) );
  XNOR2_X1 U949 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U950 ( .A(G2096), .B(KEYINPUT105), .Z(n845) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U952 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U953 ( .A(n847), .B(n846), .Z(G227) );
  NAND2_X1 U954 ( .A1(G124), .A2(n873), .ZN(n848) );
  XNOR2_X1 U955 ( .A(n848), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U956 ( .A1(G100), .A2(n877), .ZN(n849) );
  XOR2_X1 U957 ( .A(KEYINPUT107), .B(n849), .Z(n850) );
  NAND2_X1 U958 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U959 ( .A1(G136), .A2(n876), .ZN(n853) );
  NAND2_X1 U960 ( .A1(G112), .A2(n872), .ZN(n852) );
  NAND2_X1 U961 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U962 ( .A1(n855), .A2(n854), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n857) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n856) );
  XNOR2_X1 U965 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U966 ( .A(n858), .B(n925), .Z(n861) );
  XNOR2_X1 U967 ( .A(G164), .B(n859), .ZN(n860) );
  XNOR2_X1 U968 ( .A(n861), .B(n860), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G139), .A2(n876), .ZN(n863) );
  NAND2_X1 U970 ( .A1(G103), .A2(n877), .ZN(n862) );
  NAND2_X1 U971 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G115), .A2(n872), .ZN(n865) );
  NAND2_X1 U973 ( .A1(G127), .A2(n873), .ZN(n864) );
  NAND2_X1 U974 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U976 ( .A1(n868), .A2(n867), .ZN(n934) );
  XOR2_X1 U977 ( .A(n869), .B(n934), .Z(n871) );
  XNOR2_X1 U978 ( .A(G160), .B(G162), .ZN(n870) );
  XNOR2_X1 U979 ( .A(n871), .B(n870), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G118), .A2(n872), .ZN(n875) );
  NAND2_X1 U981 ( .A1(G130), .A2(n873), .ZN(n874) );
  NAND2_X1 U982 ( .A1(n875), .A2(n874), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G142), .A2(n876), .ZN(n879) );
  NAND2_X1 U984 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U985 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U986 ( .A(KEYINPUT45), .B(n880), .Z(n881) );
  XNOR2_X1 U987 ( .A(KEYINPUT108), .B(n881), .ZN(n882) );
  NOR2_X1 U988 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U989 ( .A(n885), .B(n884), .Z(n889) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U992 ( .A1(G37), .A2(n890), .ZN(G395) );
  NAND2_X1 U993 ( .A1(n891), .A2(G319), .ZN(n892) );
  NOR2_X1 U994 ( .A1(G397), .A2(n892), .ZN(n895) );
  NOR2_X1 U995 ( .A1(G229), .A2(G227), .ZN(n893) );
  XOR2_X1 U996 ( .A(KEYINPUT49), .B(n893), .Z(n894) );
  NAND2_X1 U997 ( .A1(n895), .A2(n894), .ZN(n896) );
  NOR2_X1 U998 ( .A1(n896), .A2(G395), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n897), .B(KEYINPUT111), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1001 ( .A(G1348), .B(KEYINPUT59), .ZN(n898) );
  XNOR2_X1 U1002 ( .A(n898), .B(G4), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G19), .ZN(n900) );
  XNOR2_X1 U1004 ( .A(G1981), .B(G6), .ZN(n899) );
  NOR2_X1 U1005 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U1006 ( .A1(n902), .A2(n901), .ZN(n905) );
  XOR2_X1 U1007 ( .A(KEYINPUT125), .B(G1956), .Z(n903) );
  XNOR2_X1 U1008 ( .A(G20), .B(n903), .ZN(n904) );
  NOR2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(KEYINPUT60), .B(n906), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(n907), .B(KEYINPUT126), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(G1961), .B(KEYINPUT124), .ZN(n908) );
  XNOR2_X1 U1013 ( .A(n908), .B(G5), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(G1971), .B(G22), .ZN(n910) );
  XNOR2_X1 U1015 ( .A(G1986), .B(G24), .ZN(n909) );
  NOR2_X1 U1016 ( .A1(n910), .A2(n909), .ZN(n913) );
  XNOR2_X1 U1017 ( .A(G1976), .B(KEYINPUT127), .ZN(n911) );
  XNOR2_X1 U1018 ( .A(n911), .B(G23), .ZN(n912) );
  NAND2_X1 U1019 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1020 ( .A(KEYINPUT58), .B(n914), .ZN(n915) );
  NOR2_X1 U1021 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(G21), .B(G1966), .ZN(n919) );
  NOR2_X1 U1024 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1025 ( .A(n921), .B(KEYINPUT61), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(G16), .B(KEYINPUT123), .ZN(n922) );
  NAND2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1028 ( .A1(G11), .A2(n924), .ZN(n956) );
  NOR2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G2084), .B(G160), .Z(n931) );
  XNOR2_X1 U1033 ( .A(KEYINPUT112), .B(n931), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(G2072), .B(n934), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G164), .B(G2078), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n945) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT51), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1047 ( .A(KEYINPUT52), .B(n950), .Z(n951) );
  NOR2_X1 U1048 ( .A1(KEYINPUT55), .A2(n951), .ZN(n952) );
  XOR2_X1 U1049 ( .A(KEYINPUT114), .B(n952), .Z(n953) );
  NAND2_X1 U1050 ( .A1(n953), .A2(G29), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT115), .B(n954), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n982) );
  XOR2_X1 U1053 ( .A(KEYINPUT120), .B(G29), .Z(n980) );
  XOR2_X1 U1054 ( .A(G2090), .B(G35), .Z(n959) );
  XOR2_X1 U1055 ( .A(G34), .B(KEYINPUT54), .Z(n957) );
  XNOR2_X1 U1056 ( .A(n957), .B(G2084), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n977) );
  XNOR2_X1 U1058 ( .A(n960), .B(G27), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(KEYINPUT117), .B(G2072), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(n961), .B(G33), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G25), .B(n962), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n963), .A2(G28), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(G32), .B(G1996), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT116), .B(G2067), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(G26), .B(n968), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n973), .B(KEYINPUT53), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(n975), .B(n974), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT55), .B(n978), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n1011) );
  XOR2_X1 U1077 ( .A(KEYINPUT56), .B(G16), .Z(n1009) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(KEYINPUT121), .ZN(n986) );
  XOR2_X1 U1081 ( .A(KEYINPUT57), .B(n986), .Z(n994) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n991) );
  INV_X1 U1083 ( .A(G1971), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(G166), .A2(n989), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n992), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1007) );
  XNOR2_X1 U1088 ( .A(n995), .B(G1956), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(G171), .B(G1961), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(G1348), .B(n1001), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(n1012), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

