//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT76), .B(G902), .Z(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT78), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(new_n195), .C1(G119), .C2(new_n194), .ZN(new_n196));
  XNOR2_X1  g010(.A(G119), .B(G128), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT24), .B(G110), .Z(new_n198));
  OAI22_X1  g012(.A1(new_n196), .A2(G110), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n204));
  OR3_X1    g018(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n196), .A2(G110), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n196), .A2(KEYINPUT79), .A3(G110), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n198), .A2(new_n197), .ZN(new_n216));
  INV_X1    g030(.A(new_n206), .ZN(new_n217));
  AOI21_X1  g031(.A(G146), .B1(new_n204), .B2(new_n205), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n210), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT80), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(new_n210), .C1(new_n215), .C2(new_n219), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n224), .B(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n227), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(KEYINPUT80), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n231), .B2(new_n188), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  INV_X1    g047(.A(new_n188), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n233), .B(new_n234), .C1(new_n228), .C2(new_n230), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n190), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(KEYINPUT81), .A3(new_n230), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n189), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n236), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT32), .ZN(new_n244));
  NOR2_X1   g058(.A1(G237), .A2(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G210), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n246), .B(KEYINPUT27), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G101), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n192), .A2(G116), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G119), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n250), .B2(new_n252), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT2), .B(G113), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT2), .B(G113), .Z(new_n259));
  XNOR2_X1  g073(.A(G116), .B(G119), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n250), .A2(new_n252), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT70), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n258), .A3(new_n257), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n257), .A3(new_n265), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n258), .B1(new_n263), .B2(new_n257), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n266), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G137), .ZN(new_n278));
  INV_X1    g092(.A(G137), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(KEYINPUT65), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(G134), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT11), .B1(new_n279), .B2(G134), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT65), .B(G137), .ZN(new_n286));
  AND2_X1   g100(.A1(KEYINPUT11), .A2(G134), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G131), .B1(new_n276), .B2(G137), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT66), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n279), .A2(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(G137), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n287), .ZN(new_n293));
  INV_X1    g107(.A(new_n285), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT66), .A4(new_n289), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n284), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n208), .A2(G143), .ZN(new_n300));
  INV_X1    g114(.A(G143), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G146), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT68), .ZN(new_n304));
  XNOR2_X1  g118(.A(G143), .B(G146), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n299), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n302), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT69), .B(KEYINPUT1), .C1(new_n301), .C2(G146), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G128), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT69), .B1(new_n300), .B2(KEYINPUT1), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n293), .A2(new_n294), .A3(new_n289), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n283), .B1(new_n317), .B2(new_n295), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n298), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n293), .B(new_n294), .C1(G134), .C2(new_n279), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n290), .B2(new_n296), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G128), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT64), .B1(new_n305), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(KEYINPUT0), .A2(G128), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT0), .A2(G128), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n309), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n326), .A2(new_n331), .B1(new_n305), .B2(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n274), .B1(new_n321), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n318), .A2(new_n314), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n271), .A2(new_n272), .A3(new_n266), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n272), .B1(new_n271), .B2(new_n266), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n333), .B(new_n335), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT28), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n324), .A2(new_n332), .B1(new_n318), .B2(new_n314), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n274), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT1), .B1(new_n301), .B2(G146), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G128), .A3(new_n310), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n348), .A2(new_n309), .B1(new_n304), .B2(new_n307), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n317), .A2(new_n295), .B1(G131), .B2(new_n322), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n326), .A2(new_n331), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n305), .A2(new_n327), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI22_X1  g167(.A1(new_n297), .A2(new_n349), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n341), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n249), .B1(new_n340), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT67), .B(new_n283), .C1(new_n317), .C2(new_n295), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n333), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n274), .B1(KEYINPUT30), .B2(new_n342), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n365));
  INV_X1    g179(.A(new_n249), .ZN(new_n366));
  AOI211_X1 g180(.A(new_n365), .B(new_n366), .C1(new_n274), .C2(new_n342), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT73), .B1(new_n338), .B2(new_n249), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT31), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n336), .A2(new_n337), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n249), .B1(new_n372), .B2(new_n354), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n365), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n338), .A2(KEYINPUT73), .A3(new_n249), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT31), .A3(new_n364), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n357), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G472), .A2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n244), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n340), .A2(new_n356), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n366), .ZN(new_n383));
  AOI221_X4 g197(.A(new_n370), .B1(new_n362), .B2(new_n363), .C1(new_n374), .C2(new_n375), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT31), .B1(new_n376), .B2(new_n364), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n387), .A3(KEYINPUT75), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n379), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT75), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n244), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n372), .A2(new_n354), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n338), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT28), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(new_n356), .A3(KEYINPUT29), .A4(new_n249), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n188), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n340), .A2(new_n249), .A3(new_n356), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n364), .A2(new_n338), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n400), .B2(new_n366), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G472), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n393), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n401), .A2(new_n399), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT77), .B(G472), .C1(new_n405), .C2(new_n398), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n243), .B1(new_n392), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT93), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(G101), .ZN(new_n411));
  INV_X1    g225(.A(G104), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(new_n412), .B2(G107), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n414));
  INV_X1    g228(.A(G107), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G104), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(G107), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n411), .A2(new_n413), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n418), .A2(KEYINPUT4), .B1(new_n419), .B2(G101), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(KEYINPUT4), .A3(G101), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n268), .A2(new_n422), .A3(new_n273), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n263), .A2(new_n257), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT5), .B1(new_n254), .B2(new_n255), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n426));
  INV_X1    g240(.A(G113), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n424), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT85), .B1(new_n412), .B2(G107), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n415), .A3(G104), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n433), .A3(new_n417), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n430), .A2(new_n411), .B1(new_n434), .B2(G101), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n423), .A2(new_n438), .A3(new_n436), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n443), .A3(new_n439), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n349), .A2(KEYINPUT90), .A3(new_n202), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n308), .A2(new_n202), .A3(new_n313), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n332), .B2(new_n202), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n332), .A2(new_n202), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT89), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G224), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G953), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n456), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n449), .A2(new_n453), .A3(new_n458), .A4(new_n451), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n442), .A2(new_n444), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G902), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n452), .B1(new_n445), .B2(new_n448), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(KEYINPUT7), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n449), .A2(new_n453), .A3(new_n451), .A4(new_n466), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n438), .B(KEYINPUT8), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n424), .B1(new_n428), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT91), .A3(new_n435), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n435), .B2(new_n429), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT91), .B1(new_n474), .B2(new_n435), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n441), .A2(new_n471), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n462), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n410), .B1(new_n461), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n441), .A2(new_n471), .A3(new_n478), .ZN(new_n482));
  INV_X1    g296(.A(new_n452), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n449), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT92), .B1(new_n484), .B2(new_n465), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(new_n467), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n442), .A2(new_n444), .A3(new_n460), .ZN(new_n488));
  INV_X1    g302(.A(new_n410), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G214), .B1(G237), .B2(G902), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT88), .Z(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(G113), .B(G122), .Z(new_n496));
  XOR2_X1   g310(.A(KEYINPUT95), .B(G104), .Z(new_n497));
  XOR2_X1   g311(.A(new_n496), .B(new_n497), .Z(new_n498));
  XNOR2_X1  g312(.A(new_n207), .B(KEYINPUT19), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n208), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n301), .ZN(new_n502));
  NOR2_X1   g316(.A1(KEYINPUT94), .A2(G143), .ZN(new_n503));
  OAI211_X1 g317(.A(G214), .B(new_n245), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n245), .A2(G214), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n501), .B2(new_n301), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n275), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n504), .A2(new_n506), .A3(new_n275), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n500), .B(new_n206), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(KEYINPUT18), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT18), .A2(G131), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n207), .B(new_n208), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n498), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n516));
  INV_X1    g330(.A(new_n218), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n206), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n508), .A2(new_n507), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n504), .A2(new_n506), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT17), .A3(G131), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT96), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT96), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n507), .A2(new_n525), .A3(KEYINPUT17), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n516), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n515), .B1(new_n528), .B2(new_n498), .ZN(new_n529));
  NOR2_X1   g343(.A1(G475), .A2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT20), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n518), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n522), .A2(G131), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n504), .A2(new_n506), .A3(new_n275), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n520), .A3(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n507), .A2(new_n525), .A3(KEYINPUT17), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n525), .B1(new_n507), .B2(KEYINPUT17), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n533), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n498), .A3(new_n514), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n509), .A2(new_n514), .ZN(new_n541));
  INV_X1    g355(.A(new_n498), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n530), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n194), .B2(G143), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n194), .A2(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n301), .A2(G128), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n548), .ZN(new_n553));
  OAI21_X1  g367(.A(G134), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n550), .A3(new_n276), .ZN(new_n555));
  INV_X1    g369(.A(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G116), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n251), .A2(G122), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(new_n415), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G107), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n554), .B(new_n555), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n251), .A2(KEYINPUT14), .A3(G122), .ZN(new_n564));
  OAI211_X1 g378(.A(G107), .B(new_n564), .C1(new_n561), .C2(KEYINPUT14), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n415), .ZN(new_n566));
  INV_X1    g380(.A(new_n555), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n276), .B1(new_n552), .B2(new_n550), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT9), .B(G234), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n570), .A2(new_n187), .A3(G953), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n563), .B2(new_n569), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n188), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G478), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(KEYINPUT97), .B(new_n188), .C1(new_n572), .C2(new_n573), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n574), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G952), .ZN(new_n588));
  AOI211_X1 g402(.A(G953), .B(new_n588), .C1(G234), .C2(G237), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n225), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n540), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n498), .B1(new_n539), .B2(new_n514), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n462), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G475), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n547), .A2(new_n587), .A3(new_n593), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n345), .A2(G128), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n309), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n306), .B1(new_n305), .B2(new_n299), .ZN(new_n601));
  AND4_X1   g415(.A1(new_n306), .A2(new_n299), .A3(new_n300), .A4(new_n302), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n435), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n434), .A2(G101), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n418), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n308), .A3(new_n313), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT86), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n324), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT12), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n314), .A2(KEYINPUT10), .A3(new_n435), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n332), .B1(new_n420), .B2(new_n421), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n350), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n350), .A2(KEYINPUT86), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT12), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n604), .A2(new_n607), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(G110), .B(G140), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n225), .A2(G227), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n616), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n324), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(G469), .B1(new_n634), .B2(G902), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n618), .B1(new_n617), .B2(new_n619), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT87), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT87), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n611), .A2(new_n639), .A3(new_n620), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n640), .A3(new_n630), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n628), .B1(new_n632), .B2(new_n616), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G469), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n188), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n635), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(G221), .B1(new_n570), .B2(G902), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n495), .A2(new_n598), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n408), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(new_n411), .Z(G3));
  AND3_X1   g466(.A1(new_n487), .A2(new_n489), .A3(new_n488), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n489), .B1(new_n487), .B2(new_n488), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n492), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n491), .A2(KEYINPUT99), .A3(new_n492), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n576), .A2(new_n577), .A3(new_n583), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT33), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT33), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n563), .A2(new_n569), .ZN(new_n662));
  INV_X1    g476(.A(new_n571), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(G478), .B(new_n188), .C1(new_n660), .C2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n547), .B2(new_n597), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n657), .A2(new_n658), .A3(new_n593), .A4(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n378), .B2(new_n234), .ZN(new_n671));
  INV_X1    g485(.A(new_n243), .ZN(new_n672));
  INV_X1    g486(.A(new_n648), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n635), .B2(new_n646), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n671), .A2(new_n672), .A3(new_n389), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT34), .B(G104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NAND3_X1  g492(.A1(new_n657), .A2(new_n658), .A3(new_n593), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n547), .A2(new_n597), .A3(new_n586), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NOR2_X1   g497(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n220), .B(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n242), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n223), .A2(new_n227), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n518), .A2(new_n213), .A3(new_n216), .A4(new_n214), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n222), .B1(new_n689), .B2(new_n210), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n230), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n188), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n233), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n687), .B1(new_n696), .B2(new_n190), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n598), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n491), .A3(new_n674), .A4(new_n494), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n671), .A2(new_n389), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT37), .B(G110), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  NAND2_X1  g517(.A1(new_n392), .A2(new_n407), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n649), .A2(new_n697), .ZN(new_n705));
  INV_X1    g519(.A(new_n589), .ZN(new_n706));
  INV_X1    g520(.A(new_n590), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(G900), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT100), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n680), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n657), .A2(new_n658), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n704), .A2(new_n705), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XNOR2_X1  g527(.A(new_n491), .B(KEYINPUT38), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n709), .B(KEYINPUT39), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n674), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n545), .B1(new_n544), .B2(new_n530), .ZN(new_n720));
  AOI211_X1 g534(.A(KEYINPUT20), .B(new_n531), .C1(new_n540), .C2(new_n543), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n539), .A2(new_n514), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n542), .ZN(new_n723));
  AOI21_X1  g537(.A(G902), .B1(new_n723), .B2(new_n540), .ZN(new_n724));
  INV_X1    g538(.A(G475), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n720), .A2(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n587), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n492), .A3(new_n697), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n715), .A2(new_n719), .A3(new_n729), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n376), .A2(new_n364), .B1(new_n366), .B2(new_n395), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n731), .B2(G902), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n392), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n717), .A2(new_n718), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n737));
  INV_X1    g551(.A(new_n668), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n739), .B2(new_n709), .ZN(new_n740));
  INV_X1    g554(.A(new_n709), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n669), .A2(KEYINPUT102), .A3(new_n741), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n657), .A2(new_n658), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n704), .A2(new_n705), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  INV_X1    g559(.A(new_n670), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n611), .A2(new_n620), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n629), .B1(new_n747), .B2(KEYINPUT87), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n642), .B1(new_n748), .B2(new_n640), .ZN(new_n749));
  OAI21_X1  g563(.A(G469), .B1(new_n749), .B2(new_n234), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n648), .A3(new_n646), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n750), .A2(new_n646), .A3(KEYINPUT103), .A4(new_n648), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n408), .A2(new_n746), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NOR2_X1   g573(.A1(new_n679), .A2(new_n680), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n408), .A2(new_n760), .A3(new_n756), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G116), .ZN(G18));
  AOI22_X1  g576(.A1(new_n388), .A2(new_n391), .B1(new_n404), .B2(new_n406), .ZN(new_n763));
  INV_X1    g577(.A(new_n751), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n657), .A2(new_n658), .A3(new_n698), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n192), .ZN(G21));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n593), .A3(new_n754), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n249), .B1(new_n396), .B2(new_n356), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n371), .B2(new_n377), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n771), .B2(new_n380), .ZN(new_n772));
  INV_X1    g586(.A(new_n770), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n384), .B2(new_n385), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT104), .A3(new_n379), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n671), .A2(new_n772), .A3(new_n775), .A4(new_n672), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n657), .A2(new_n658), .A3(new_n728), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G122), .ZN(G24));
  AOI21_X1  g594(.A(KEYINPUT102), .B1(new_n669), .B2(new_n741), .ZN(new_n781));
  AND4_X1   g595(.A1(KEYINPUT102), .A2(new_n726), .A3(new_n738), .A4(new_n741), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT105), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n740), .A2(new_n742), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n697), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n671), .A2(new_n772), .A3(new_n775), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n657), .A2(new_n764), .A3(new_n658), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G125), .ZN(G27));
  NAND3_X1  g606(.A1(new_n481), .A2(new_n490), .A3(new_n492), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n649), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n783), .A3(new_n785), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT42), .B1(new_n408), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n381), .A2(new_n387), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n407), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n672), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n783), .A3(KEYINPUT42), .A4(new_n785), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT106), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n796), .A2(KEYINPUT42), .A3(new_n672), .A4(new_n800), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n763), .A2(new_n795), .A3(new_n243), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(KEYINPUT42), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n275), .ZN(G33));
  AND2_X1   g624(.A1(new_n794), .A2(new_n710), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n704), .A2(new_n811), .A3(new_n672), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G134), .ZN(G36));
  NAND2_X1  g627(.A1(new_n727), .A2(new_n738), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT43), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n697), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(KEYINPUT44), .A3(new_n700), .ZN(new_n817));
  INV_X1    g631(.A(new_n793), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT107), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT107), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT44), .B1(new_n816), .B2(new_n700), .ZN(new_n822));
  INV_X1    g636(.A(new_n646), .ZN(new_n823));
  NAND2_X1  g637(.A1(G469), .A2(G902), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n634), .A2(KEYINPUT45), .ZN(new_n825));
  OAI21_X1  g639(.A(G469), .B1(new_n634), .B2(KEYINPUT45), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT46), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n648), .A3(new_n716), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n820), .A2(new_n821), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G137), .ZN(G39));
  NOR4_X1   g648(.A1(new_n781), .A2(new_n793), .A3(new_n672), .A4(new_n782), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n763), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT108), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n830), .A2(new_n648), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT47), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n830), .A2(KEYINPUT47), .A3(new_n648), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(KEYINPUT108), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT109), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G140), .ZN(G42));
  INV_X1    g661(.A(new_n750), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n848), .A2(new_n823), .A3(KEYINPUT49), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT49), .B1(new_n848), .B2(new_n823), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n814), .A2(new_n493), .A3(new_n673), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n672), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n733), .A2(new_n714), .A3(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n793), .A2(new_n726), .A3(new_n586), .A4(new_n709), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n704), .A2(new_n705), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n789), .A2(new_n794), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n812), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n763), .A2(new_n670), .A3(new_n755), .A4(new_n243), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n672), .A2(new_n671), .A3(new_n772), .A4(new_n775), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n753), .A2(new_n593), .A3(new_n754), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n657), .A2(new_n658), .A3(new_n728), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n861), .A2(new_n862), .B1(new_n763), .B2(new_n765), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n592), .B1(new_n739), .B2(new_n680), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n491), .A3(new_n494), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n675), .A2(new_n866), .B1(new_n699), .B2(new_n700), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n408), .B2(new_n650), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n857), .A2(new_n864), .A3(new_n761), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n809), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT110), .B1(new_n697), .B2(new_n741), .ZN(new_n872));
  INV_X1    g686(.A(new_n687), .ZN(new_n873));
  AND4_X1   g687(.A1(KEYINPUT110), .A2(new_n236), .A3(new_n873), .A4(new_n741), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n674), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT111), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n674), .C1(new_n872), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n733), .A3(new_n778), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n712), .A3(new_n744), .A4(new_n791), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  OR3_X1    g696(.A1(new_n881), .A2(KEYINPUT112), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  INV_X1    g698(.A(new_n705), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n392), .B2(new_n407), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n886), .A2(new_n711), .B1(new_n789), .B2(new_n790), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(KEYINPUT52), .A3(new_n744), .A4(new_n880), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(KEYINPUT112), .A3(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n870), .A2(new_n871), .A3(new_n883), .A4(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n884), .A2(new_n888), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n812), .A2(new_n855), .A3(new_n856), .ZN(new_n892));
  INV_X1    g706(.A(new_n867), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n651), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n765), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n704), .A2(new_n896), .B1(new_n777), .B2(new_n778), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n897), .A2(new_n757), .A3(new_n761), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n895), .A2(new_n898), .A3(new_n804), .A4(new_n808), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT53), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n890), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n871), .B1(new_n891), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT53), .B1(new_n797), .B2(new_n803), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n408), .A2(new_n811), .B1(new_n789), .B2(new_n794), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n868), .A3(new_n855), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n897), .A2(new_n757), .A3(new_n761), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n889), .A3(new_n883), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n902), .A2(KEYINPUT113), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT113), .B1(new_n902), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n818), .A2(new_n764), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n733), .A2(new_n243), .A3(new_n706), .A4(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT116), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n916), .A2(new_n726), .A3(new_n738), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n815), .A2(new_n706), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n918), .A2(new_n788), .A3(new_n914), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n776), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT50), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n492), .B1(KEYINPUT115), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n920), .A2(new_n715), .A3(new_n764), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(KEYINPUT115), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n823), .A2(new_n848), .A3(new_n648), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n842), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n818), .ZN(new_n928));
  OAI221_X1 g742(.A(new_n925), .B1(new_n924), .B2(new_n923), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT114), .B1(new_n917), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT51), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(KEYINPUT51), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n916), .A2(new_n739), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n801), .A2(new_n918), .A3(new_n914), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT48), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n920), .A2(new_n790), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(G952), .A3(new_n225), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n932), .A3(new_n938), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n912), .A2(new_n913), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(G952), .A2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n853), .B1(new_n940), .B2(new_n941), .ZN(G75));
  NAND2_X1  g756(.A1(new_n442), .A2(new_n444), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(new_n460), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n489), .A2(new_n188), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n903), .B2(new_n909), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n948), .B2(KEYINPUT56), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(KEYINPUT117), .B(new_n945), .C1(new_n948), .C2(KEYINPUT56), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n225), .A2(G952), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n945), .B(KEYINPUT119), .Z(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT56), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n884), .A2(new_n888), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT53), .B1(new_n870), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n908), .A2(new_n889), .A3(new_n883), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n946), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT118), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n948), .A2(KEYINPUT118), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n953), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT120), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n953), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G51));
  NAND2_X1  g783(.A1(new_n903), .A2(new_n909), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT54), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n911), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n824), .B(KEYINPUT57), .Z(new_n973));
  AOI21_X1  g787(.A(new_n749), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT121), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n234), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(new_n825), .A3(new_n826), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n974), .B2(KEYINPUT121), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n954), .B1(new_n975), .B2(new_n978), .ZN(G54));
  INV_X1    g793(.A(new_n954), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT58), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n976), .A2(new_n981), .A3(new_n725), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n982), .B2(new_n544), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n544), .B2(new_n982), .ZN(G60));
  INV_X1    g798(.A(new_n972), .ZN(new_n985));
  NAND2_X1  g799(.A1(G478), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT59), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n660), .B2(new_n666), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n980), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n987), .B1(new_n912), .B2(new_n913), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n660), .A2(new_n666), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT60), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n970), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n980), .B1(new_n995), .B2(new_n686), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT122), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT61), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n240), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n999), .B(new_n980), .C1(new_n686), .C2(new_n995), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(G66));
  OAI21_X1  g815(.A(G953), .B1(new_n591), .B2(new_n455), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n907), .A2(new_n894), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n943), .B1(G898), .B2(new_n225), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  OAI21_X1  g821(.A(new_n362), .B1(new_n361), .B2(new_n354), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(new_n499), .Z(new_n1009));
  NAND2_X1  g823(.A1(new_n887), .A2(new_n744), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1010), .A2(KEYINPUT124), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(KEYINPUT124), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n735), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1011), .A2(new_n1015), .A3(new_n735), .A4(new_n1012), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n793), .B1(new_n739), .B2(new_n680), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n408), .A2(new_n674), .A3(new_n716), .A4(new_n1017), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n833), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1014), .A2(new_n846), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1009), .B1(new_n1020), .B2(new_n225), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1021), .A2(KEYINPUT125), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(KEYINPUT125), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1011), .A2(new_n833), .A3(new_n1012), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n831), .A2(new_n801), .A3(new_n862), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n408), .B2(new_n811), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n804), .A2(new_n846), .A3(new_n808), .A4(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1025), .A2(new_n1028), .A3(new_n225), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G900), .A2(G953), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1029), .A2(new_n1009), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1022), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n225), .B1(G227), .B2(G900), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1033), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1022), .A2(new_n1035), .A3(new_n1023), .A4(new_n1031), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1034), .A2(new_n1036), .ZN(G72));
  NAND3_X1  g851(.A1(new_n1025), .A2(new_n1028), .A3(new_n1003), .ZN(new_n1038));
  NAND2_X1  g852(.A1(G472), .A2(G902), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT63), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT127), .ZN(new_n1041));
  AOI211_X1 g855(.A(new_n249), .B(new_n400), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n400), .A2(new_n249), .ZN(new_n1043));
  OR3_X1    g857(.A1(new_n1020), .A2(new_n907), .A3(new_n894), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1043), .B1(new_n1044), .B2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n400), .A2(new_n366), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1040), .B1(new_n1046), .B2(new_n369), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n901), .A2(new_n1047), .ZN(new_n1048));
  NOR4_X1   g862(.A1(new_n1042), .A2(new_n1045), .A3(new_n954), .A4(new_n1048), .ZN(G57));
endmodule


