

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811;

  OR2_X1 U376 ( .A1(n634), .A2(n536), .ZN(n535) );
  XNOR2_X1 U377 ( .A(n387), .B(n590), .ZN(n784) );
  BUF_X1 U378 ( .A(G237), .Z(n355) );
  NOR2_X1 U379 ( .A1(n711), .A2(n723), .ZN(n656) );
  XNOR2_X2 U380 ( .A(n448), .B(n447), .ZN(n711) );
  NOR2_X2 U381 ( .A1(n602), .A2(n601), .ZN(n735) );
  NAND2_X2 U382 ( .A1(n627), .A2(n361), .ZN(n426) );
  NOR2_X2 U383 ( .A1(n745), .A2(n519), .ZN(n520) );
  XNOR2_X2 U384 ( .A(n585), .B(n395), .ZN(n394) );
  XNOR2_X2 U385 ( .A(n595), .B(n594), .ZN(n601) );
  XNOR2_X2 U386 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X2 U387 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U388 ( .A(n406), .B(n571), .ZN(n389) );
  XNOR2_X2 U389 ( .A(n517), .B(G902), .ZN(n668) );
  XNOR2_X1 U390 ( .A(n390), .B(n389), .ZN(n388) );
  XNOR2_X1 U391 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n571) );
  INV_X2 U392 ( .A(KEYINPUT4), .ZN(n407) );
  XNOR2_X1 U393 ( .A(G122), .B(G107), .ZN(n578) );
  INV_X1 U394 ( .A(G953), .ZN(n802) );
  XOR2_X1 U395 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n356) );
  XOR2_X1 U396 ( .A(KEYINPUT30), .B(KEYINPUT109), .Z(n357) );
  XOR2_X1 U397 ( .A(KEYINPUT67), .B(KEYINPUT1), .Z(n358) );
  XNOR2_X2 U398 ( .A(n411), .B(n427), .ZN(n693) );
  AND2_X2 U399 ( .A1(n384), .A2(n417), .ZN(n420) );
  NAND2_X2 U400 ( .A1(n416), .A2(n422), .ZN(n415) );
  AND2_X2 U401 ( .A1(n418), .A2(n423), .ZN(n417) );
  XNOR2_X2 U402 ( .A(n567), .B(n412), .ZN(n597) );
  NAND2_X2 U403 ( .A1(n598), .A2(n736), .ZN(n372) );
  XNOR2_X2 U404 ( .A(n623), .B(KEYINPUT38), .ZN(n598) );
  XOR2_X1 U405 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n572) );
  XNOR2_X1 U406 ( .A(n574), .B(n572), .ZN(n390) );
  XNOR2_X1 U407 ( .A(n370), .B(n391), .ZN(n679) );
  XNOR2_X1 U408 ( .A(n388), .B(n784), .ZN(n370) );
  INV_X1 U409 ( .A(n377), .ZN(n655) );
  NOR2_X2 U410 ( .A1(G953), .A2(G237), .ZN(n584) );
  XNOR2_X1 U411 ( .A(n489), .B(n397), .ZN(n541) );
  INV_X1 U412 ( .A(n811), .ZN(n473) );
  NAND2_X1 U413 ( .A1(n537), .A2(n535), .ZN(n499) );
  AND2_X1 U414 ( .A1(n539), .A2(n538), .ZN(n537) );
  OR2_X1 U415 ( .A1(n779), .A2(G902), .ZN(n382) );
  XNOR2_X1 U416 ( .A(n516), .B(KEYINPUT20), .ZN(n557) );
  NAND2_X1 U417 ( .A1(n436), .A2(n467), .ZN(n531) );
  NAND2_X1 U418 ( .A1(n537), .A2(n535), .ZN(n651) );
  AND2_X1 U419 ( .A1(n450), .A2(n654), .ZN(n449) );
  AND2_X1 U420 ( .A1(n735), .A2(n359), .ZN(n433) );
  XNOR2_X1 U421 ( .A(n409), .B(KEYINPUT105), .ZN(n720) );
  NAND2_X1 U422 ( .A1(n601), .A2(n600), .ZN(n409) );
  NAND2_X1 U423 ( .A1(n749), .A2(n359), .ZN(n745) );
  NOR2_X1 U424 ( .A1(n749), .A2(n514), .ZN(n612) );
  INV_X1 U425 ( .A(n639), .ZN(n359) );
  OR2_X1 U426 ( .A1(n687), .A2(G902), .ZN(n439) );
  NAND2_X1 U427 ( .A1(n557), .A2(G217), .ZN(n381) );
  XNOR2_X1 U428 ( .A(n589), .B(n360), .ZN(n796) );
  XNOR2_X1 U429 ( .A(n566), .B(n360), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n564), .B(n356), .ZN(n378) );
  NAND2_X1 U431 ( .A1(G214), .A2(n576), .ZN(n736) );
  XNOR2_X1 U432 ( .A(n503), .B(G146), .ZN(n569) );
  INV_X1 U433 ( .A(n563), .ZN(n360) );
  XNOR2_X2 U434 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n517) );
  OR2_X1 U435 ( .A1(n355), .A2(G902), .ZN(n576) );
  XNOR2_X1 U436 ( .A(G128), .B(G110), .ZN(n548) );
  XOR2_X1 U437 ( .A(G137), .B(G140), .Z(n563) );
  INV_X1 U438 ( .A(G478), .ZN(n438) );
  INV_X2 U439 ( .A(G125), .ZN(n503) );
  INV_X1 U440 ( .A(KEYINPUT12), .ZN(n395) );
  XOR2_X1 U441 ( .A(G122), .B(G104), .Z(n590) );
  INV_X1 U442 ( .A(KEYINPUT4), .ZN(n797) );
  INV_X1 U443 ( .A(KEYINPUT98), .ZN(n447) );
  XNOR2_X1 U444 ( .A(n455), .B(n674), .ZN(n727) );
  NAND2_X1 U445 ( .A1(n458), .A2(n456), .ZN(n455) );
  AND2_X1 U446 ( .A1(n431), .A2(n666), .ZN(n404) );
  XNOR2_X1 U447 ( .A(n531), .B(n530), .ZN(n501) );
  XNOR2_X1 U448 ( .A(n440), .B(n617), .ZN(n364) );
  NOR2_X1 U449 ( .A1(n661), .A2(n645), .ZN(n646) );
  BUF_X1 U450 ( .A(n711), .Z(n363) );
  NOR2_X1 U451 ( .A1(n463), .A2(n660), .ZN(n662) );
  NAND2_X1 U452 ( .A1(n442), .A2(n441), .ZN(n440) );
  AND2_X1 U453 ( .A1(n443), .A2(n484), .ZN(n442) );
  NAND2_X1 U454 ( .A1(n444), .A2(n486), .ZN(n441) );
  NAND2_X1 U455 ( .A1(n434), .A2(n433), .ZN(n641) );
  NOR2_X1 U456 ( .A1(n607), .A2(n424), .ZN(n422) );
  NAND2_X1 U457 ( .A1(n453), .A2(n376), .ZN(n607) );
  XNOR2_X1 U458 ( .A(n636), .B(KEYINPUT33), .ZN(n743) );
  XNOR2_X1 U459 ( .A(n454), .B(n498), .ZN(n453) );
  NAND2_X1 U460 ( .A1(n408), .A2(n720), .ZN(n620) );
  NAND2_X1 U461 ( .A1(n655), .A2(n612), .ZN(n454) );
  AND2_X1 U462 ( .A1(n642), .A2(n612), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n445), .B(n357), .ZN(n521) );
  BUF_X1 U464 ( .A(n720), .Z(n361) );
  BUF_X1 U465 ( .A(n746), .Z(n398) );
  INV_X1 U466 ( .A(n597), .ZN(n376) );
  XNOR2_X1 U467 ( .A(n597), .B(n358), .ZN(n746) );
  NAND2_X2 U468 ( .A1(n482), .A2(n478), .ZN(n377) );
  XNOR2_X1 U469 ( .A(n439), .B(n437), .ZN(n600) );
  AND2_X1 U470 ( .A1(n428), .A2(n483), .ZN(n482) );
  NOR2_X1 U471 ( .A1(n700), .A2(G902), .ZN(n595) );
  XNOR2_X1 U472 ( .A(n526), .B(n528), .ZN(n687) );
  XNOR2_X1 U473 ( .A(n558), .B(n393), .ZN(n748) );
  XNOR2_X1 U474 ( .A(n383), .B(n796), .ZN(n779) );
  XNOR2_X1 U475 ( .A(n381), .B(n380), .ZN(n379) );
  XNOR2_X1 U476 ( .A(n365), .B(n591), .ZN(n700) );
  XNOR2_X1 U477 ( .A(n411), .B(n399), .ZN(n773) );
  XNOR2_X1 U478 ( .A(n375), .B(n374), .ZN(n399) );
  XNOR2_X1 U479 ( .A(n575), .B(n392), .ZN(n391) );
  XNOR2_X1 U480 ( .A(n509), .B(n545), .ZN(n383) );
  OR2_X1 U481 ( .A1(n633), .A2(KEYINPUT0), .ZN(n536) );
  XNOR2_X1 U482 ( .A(n368), .B(n366), .ZN(n365) );
  XNOR2_X1 U483 ( .A(n394), .B(n588), .ZN(n368) );
  XNOR2_X1 U484 ( .A(n378), .B(n400), .ZN(n410) );
  XNOR2_X1 U485 ( .A(n583), .B(n527), .ZN(n526) );
  XNOR2_X1 U486 ( .A(n533), .B(n561), .ZN(n392) );
  XNOR2_X1 U487 ( .A(n549), .B(n546), .ZN(n509) );
  XNOR2_X1 U488 ( .A(n586), .B(n367), .ZN(n366) );
  XNOR2_X1 U489 ( .A(n570), .B(n505), .ZN(n504) );
  XNOR2_X1 U490 ( .A(n564), .B(n452), .ZN(n374) );
  XNOR2_X1 U491 ( .A(n507), .B(n506), .ZN(n581) );
  INV_X1 U492 ( .A(n736), .ZN(n446) );
  XNOR2_X1 U493 ( .A(n401), .B(G137), .ZN(n400) );
  XNOR2_X1 U494 ( .A(n569), .B(n508), .ZN(n589) );
  XNOR2_X1 U495 ( .A(n559), .B(n560), .ZN(n393) );
  XNOR2_X1 U496 ( .A(n438), .B(KEYINPUT104), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U498 ( .A(n425), .ZN(n386) );
  INV_X1 U499 ( .A(n667), .ZN(n397) );
  XNOR2_X1 U500 ( .A(n550), .B(n515), .ZN(n380) );
  XNOR2_X1 U501 ( .A(n568), .B(KEYINPUT16), .ZN(n387) );
  XOR2_X1 U502 ( .A(G140), .B(KEYINPUT11), .Z(n586) );
  INV_X1 U503 ( .A(KEYINPUT8), .ZN(n506) );
  XOR2_X1 U504 ( .A(G119), .B(KEYINPUT24), .Z(n546) );
  INV_X1 U505 ( .A(KEYINPUT18), .ZN(n505) );
  INV_X2 U506 ( .A(KEYINPUT70), .ZN(n532) );
  XNOR2_X1 U507 ( .A(KEYINPUT90), .B(G104), .ZN(n452) );
  INV_X1 U508 ( .A(G902), .ZN(n480) );
  XNOR2_X1 U509 ( .A(KEYINPUT69), .B(G131), .ZN(n587) );
  NAND2_X1 U510 ( .A1(G953), .A2(G902), .ZN(n630) );
  INV_X1 U511 ( .A(KEYINPUT42), .ZN(n424) );
  INV_X1 U512 ( .A(n499), .ZN(n434) );
  XNOR2_X1 U513 ( .A(n646), .B(KEYINPUT32), .ZN(n811) );
  XNOR2_X1 U514 ( .A(n637), .B(n470), .ZN(n436) );
  XNOR2_X2 U515 ( .A(n614), .B(n606), .ZN(n634) );
  AND2_X1 U516 ( .A1(n362), .A2(n364), .ZN(n477) );
  XNOR2_X1 U517 ( .A(n510), .B(KEYINPUT73), .ZN(n362) );
  XNOR2_X1 U518 ( .A(n364), .B(n691), .ZN(G27) );
  INV_X1 U519 ( .A(n587), .ZN(n367) );
  XNOR2_X2 U520 ( .A(n369), .B(n469), .ZN(n605) );
  NAND2_X1 U521 ( .A1(n679), .A2(n668), .ZN(n369) );
  XNOR2_X2 U522 ( .A(n371), .B(n596), .ZN(n729) );
  NAND2_X1 U523 ( .A1(n734), .A2(n735), .ZN(n371) );
  XNOR2_X2 U524 ( .A(n372), .B(n577), .ZN(n734) );
  NAND2_X1 U525 ( .A1(n414), .A2(n373), .ZN(n413) );
  NAND2_X1 U526 ( .A1(n420), .A2(n373), .ZN(n419) );
  XNOR2_X1 U527 ( .A(n373), .B(G131), .ZN(G33) );
  XNOR2_X2 U528 ( .A(n426), .B(KEYINPUT40), .ZN(n373) );
  XNOR2_X2 U529 ( .A(n407), .B(G101), .ZN(n564) );
  NAND2_X1 U530 ( .A1(n376), .A2(n466), .ZN(n519) );
  NOR2_X1 U531 ( .A1(n377), .A2(n446), .ZN(n445) );
  NOR2_X1 U532 ( .A1(n745), .A2(n377), .ZN(n649) );
  XNOR2_X2 U533 ( .A(n377), .B(KEYINPUT6), .ZN(n642) );
  NAND2_X1 U534 ( .A1(n753), .A2(n450), .ZN(n755) );
  INV_X1 U535 ( .A(n564), .ZN(n561) );
  XNOR2_X2 U536 ( .A(n382), .B(n379), .ZN(n749) );
  AND2_X2 U537 ( .A1(n417), .A2(n415), .ZN(n414) );
  INV_X1 U538 ( .A(n385), .ZN(n384) );
  NAND2_X1 U539 ( .A1(n415), .A2(n386), .ZN(n385) );
  INV_X1 U540 ( .A(n414), .ZN(n496) );
  NAND2_X2 U541 ( .A1(n405), .A2(n404), .ZN(n489) );
  NAND2_X1 U542 ( .A1(n605), .A2(n736), .ZN(n614) );
  INV_X1 U543 ( .A(KEYINPUT46), .ZN(n425) );
  INV_X2 U544 ( .A(n605), .ZN(n623) );
  XNOR2_X1 U545 ( .A(n396), .B(n618), .ZN(n475) );
  NAND2_X1 U546 ( .A1(n476), .A2(n477), .ZN(n396) );
  XNOR2_X2 U547 ( .A(n798), .B(G146), .ZN(n411) );
  XNOR2_X2 U548 ( .A(n583), .B(n587), .ZN(n798) );
  XNOR2_X2 U549 ( .A(n573), .B(G134), .ZN(n583) );
  NAND2_X1 U550 ( .A1(n584), .A2(G210), .ZN(n401) );
  AND2_X2 U551 ( .A1(n403), .A2(n402), .ZN(n405) );
  AND2_X1 U552 ( .A1(n664), .A2(n705), .ZN(n402) );
  NAND2_X1 U553 ( .A1(n429), .A2(n474), .ZN(n403) );
  XNOR2_X1 U554 ( .A(n406), .B(n533), .ZN(n497) );
  XNOR2_X2 U555 ( .A(n532), .B(G119), .ZN(n406) );
  XNOR2_X2 U556 ( .A(n620), .B(n613), .ZN(n488) );
  XNOR2_X1 U557 ( .A(n410), .B(n497), .ZN(n427) );
  XNOR2_X2 U558 ( .A(n534), .B(G116), .ZN(n533) );
  INV_X1 U559 ( .A(G469), .ZN(n412) );
  NAND2_X1 U560 ( .A1(n413), .A2(n425), .ZN(n421) );
  INV_X1 U561 ( .A(n729), .ZN(n416) );
  NAND2_X1 U562 ( .A1(n729), .A2(n424), .ZN(n418) );
  NAND2_X1 U563 ( .A1(n421), .A2(n419), .ZN(n476) );
  NAND2_X1 U564 ( .A1(n607), .A2(n424), .ZN(n423) );
  NAND2_X1 U565 ( .A1(n693), .A2(n562), .ZN(n428) );
  NAND2_X1 U566 ( .A1(n430), .A2(KEYINPUT66), .ZN(n429) );
  NAND2_X1 U567 ( .A1(n518), .A2(n638), .ZN(n430) );
  NAND2_X1 U568 ( .A1(n432), .A2(n665), .ZN(n431) );
  NAND2_X1 U569 ( .A1(n473), .A2(n471), .ZN(n432) );
  NAND2_X1 U570 ( .A1(n435), .A2(KEYINPUT44), .ZN(n666) );
  INV_X1 U571 ( .A(n501), .ZN(n435) );
  NAND2_X1 U572 ( .A1(n488), .A2(n487), .ZN(n443) );
  INV_X1 U573 ( .A(n488), .ZN(n444) );
  NAND2_X1 U574 ( .A1(n451), .A2(n449), .ZN(n448) );
  INV_X1 U575 ( .A(n655), .ZN(n450) );
  XNOR2_X1 U576 ( .A(n499), .B(KEYINPUT89), .ZN(n451) );
  NOR2_X2 U577 ( .A1(n607), .A2(n634), .ZN(n718) );
  XNOR2_X1 U578 ( .A(n457), .B(KEYINPUT83), .ZN(n456) );
  NAND2_X1 U579 ( .A1(n673), .A2(KEYINPUT2), .ZN(n457) );
  INV_X1 U580 ( .A(n459), .ZN(n458) );
  XNOR2_X1 U581 ( .A(n522), .B(n671), .ZN(n676) );
  XNOR2_X1 U582 ( .A(n489), .B(n667), .ZN(n459) );
  INV_X1 U583 ( .A(n494), .ZN(n460) );
  NAND2_X1 U584 ( .A1(n676), .A2(n675), .ZN(n461) );
  NAND2_X1 U585 ( .A1(n676), .A2(n675), .ZN(n678) );
  INV_X1 U586 ( .A(n473), .ZN(n462) );
  XNOR2_X1 U587 ( .A(n641), .B(n640), .ZN(n463) );
  XNOR2_X1 U588 ( .A(n641), .B(n640), .ZN(n661) );
  INV_X1 U589 ( .A(n673), .ZN(n464) );
  NAND2_X1 U590 ( .A1(n475), .A2(n629), .ZN(n672) );
  BUF_X1 U591 ( .A(n734), .Z(n465) );
  XNOR2_X2 U592 ( .A(n461), .B(n677), .ZN(n770) );
  NAND2_X1 U593 ( .A1(n544), .A2(n763), .ZN(n633) );
  NAND2_X1 U594 ( .A1(n481), .A2(n480), .ZN(n479) );
  XNOR2_X1 U595 ( .A(n531), .B(n492), .ZN(n518) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT68), .ZN(n492) );
  INV_X1 U597 ( .A(KEYINPUT68), .ZN(n472) );
  NAND2_X1 U598 ( .A1(n668), .A2(G234), .ZN(n516) );
  AND2_X1 U599 ( .A1(n615), .A2(n616), .ZN(n487) );
  NAND2_X1 U600 ( .A1(n633), .A2(KEYINPUT0), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n802), .A2(G234), .ZN(n507) );
  XNOR2_X1 U602 ( .A(n579), .B(KEYINPUT102), .ZN(n527) );
  INV_X1 U603 ( .A(KEYINPUT10), .ZN(n508) );
  XNOR2_X1 U604 ( .A(G143), .B(G113), .ZN(n588) );
  INV_X1 U605 ( .A(n616), .ZN(n486) );
  INV_X1 U606 ( .A(KEYINPUT91), .ZN(n515) );
  NAND2_X1 U607 ( .A1(n562), .A2(G902), .ZN(n483) );
  XOR2_X1 U608 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n550) );
  INV_X1 U609 ( .A(KEYINPUT23), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n504), .B(n569), .ZN(n575) );
  NAND2_X1 U611 ( .A1(n355), .A2(G234), .ZN(n551) );
  AND2_X1 U612 ( .A1(n485), .A2(n650), .ZN(n484) );
  NAND2_X1 U613 ( .A1(n500), .A2(n486), .ZN(n485) );
  INV_X1 U614 ( .A(KEYINPUT35), .ZN(n530) );
  INV_X1 U615 ( .A(KEYINPUT28), .ZN(n498) );
  XNOR2_X1 U616 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n640) );
  XNOR2_X1 U617 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U618 ( .A(n582), .B(n529), .ZN(n528) );
  XNOR2_X1 U619 ( .A(n580), .B(n578), .ZN(n529) );
  AND2_X1 U620 ( .A1(n766), .A2(G953), .ZN(n783) );
  AND2_X1 U621 ( .A1(n467), .A2(n494), .ZN(n525) );
  NOR2_X1 U622 ( .A1(n745), .A2(n597), .ZN(n654) );
  OR2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n466) );
  AND2_X1 U624 ( .A1(n602), .A2(n601), .ZN(n467) );
  AND2_X1 U625 ( .A1(n541), .A2(n540), .ZN(n468) );
  AND2_X1 U626 ( .A1(G210), .A2(n576), .ZN(n469) );
  XNOR2_X1 U627 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n470) );
  NOR2_X1 U628 ( .A1(n811), .A2(n714), .ZN(n474) );
  NOR2_X1 U629 ( .A1(n714), .A2(n472), .ZN(n471) );
  OR2_X1 U630 ( .A1(n693), .A2(n479), .ZN(n478) );
  INV_X1 U631 ( .A(n562), .ZN(n481) );
  NAND2_X1 U632 ( .A1(n490), .A2(n521), .ZN(n717) );
  AND2_X1 U633 ( .A1(n525), .A2(n520), .ZN(n490) );
  NAND2_X1 U634 ( .A1(n491), .A2(n521), .ZN(n599) );
  AND2_X1 U635 ( .A1(n520), .A2(n737), .ZN(n491) );
  XNOR2_X2 U636 ( .A(n678), .B(n677), .ZN(n493) );
  INV_X1 U637 ( .A(n623), .ZN(n494) );
  XNOR2_X1 U638 ( .A(n464), .B(KEYINPUT82), .ZN(n495) );
  XNOR2_X1 U639 ( .A(n672), .B(KEYINPUT82), .ZN(n801) );
  NAND2_X1 U640 ( .A1(n511), .A2(n611), .ZN(n510) );
  BUF_X1 U641 ( .A(n598), .Z(n737) );
  BUF_X1 U642 ( .A(n614), .Z(n500) );
  XNOR2_X1 U643 ( .A(n651), .B(KEYINPUT89), .ZN(n502) );
  NAND2_X1 U644 ( .A1(n502), .A2(n743), .ZN(n637) );
  NAND2_X1 U645 ( .A1(n513), .A2(n512), .ZN(n511) );
  NAND2_X1 U646 ( .A1(n718), .A2(KEYINPUT47), .ZN(n512) );
  NAND2_X1 U647 ( .A1(n610), .A2(n609), .ZN(n513) );
  NAND2_X1 U648 ( .A1(n748), .A2(n466), .ZN(n514) );
  NAND2_X1 U649 ( .A1(n523), .A2(n670), .ZN(n522) );
  XNOR2_X1 U650 ( .A(n524), .B(KEYINPUT80), .ZN(n523) );
  NAND2_X1 U651 ( .A1(n542), .A2(n541), .ZN(n524) );
  NAND2_X1 U652 ( .A1(n717), .A2(n603), .ZN(n604) );
  XNOR2_X2 U653 ( .A(G113), .B(KEYINPUT3), .ZN(n534) );
  NAND2_X1 U654 ( .A1(n634), .A2(KEYINPUT0), .ZN(n539) );
  INV_X1 U655 ( .A(n495), .ZN(n540) );
  NOR2_X1 U656 ( .A1(n801), .A2(n668), .ZN(n542) );
  AND2_X1 U657 ( .A1(G227), .A2(n802), .ZN(n543) );
  OR2_X1 U658 ( .A1(n632), .A2(n631), .ZN(n544) );
  INV_X1 U659 ( .A(n573), .ZN(n574) );
  INV_X1 U660 ( .A(KEYINPUT65), .ZN(n671) );
  INV_X1 U661 ( .A(KEYINPUT110), .ZN(n577) );
  XNOR2_X1 U662 ( .A(n565), .B(n543), .ZN(n566) );
  XNOR2_X1 U663 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n596) );
  INV_X1 U664 ( .A(KEYINPUT123), .ZN(n778) );
  NAND2_X1 U665 ( .A1(G221), .A2(n581), .ZN(n545) );
  XNOR2_X1 U666 ( .A(n551), .B(KEYINPUT14), .ZN(n763) );
  INV_X1 U667 ( .A(n763), .ZN(n552) );
  NOR2_X1 U668 ( .A1(n552), .A2(n630), .ZN(n553) );
  XOR2_X1 U669 ( .A(KEYINPUT106), .B(n553), .Z(n554) );
  NOR2_X1 U670 ( .A1(G900), .A2(n554), .ZN(n556) );
  INV_X1 U671 ( .A(G952), .ZN(n766) );
  NOR2_X1 U672 ( .A1(G953), .A2(n766), .ZN(n632) );
  AND2_X1 U673 ( .A1(n632), .A2(n763), .ZN(n555) );
  XOR2_X1 U674 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n559) );
  NAND2_X1 U675 ( .A1(n557), .A2(G221), .ZN(n558) );
  INV_X1 U676 ( .A(KEYINPUT21), .ZN(n560) );
  XNOR2_X2 U677 ( .A(G143), .B(G128), .ZN(n573) );
  XNOR2_X1 U678 ( .A(G472), .B(KEYINPUT97), .ZN(n562) );
  XNOR2_X2 U679 ( .A(G107), .B(G110), .ZN(n568) );
  INV_X1 U680 ( .A(n568), .ZN(n565) );
  NAND2_X1 U681 ( .A1(n773), .A2(n480), .ZN(n567) );
  NAND2_X1 U682 ( .A1(G224), .A2(n802), .ZN(n570) );
  XOR2_X1 U683 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n580) );
  XNOR2_X1 U684 ( .A(G116), .B(KEYINPUT7), .ZN(n579) );
  NAND2_X1 U685 ( .A1(G217), .A2(n581), .ZN(n582) );
  INV_X1 U686 ( .A(n600), .ZN(n602) );
  NAND2_X1 U687 ( .A1(n584), .A2(G214), .ZN(n585) );
  XNOR2_X1 U688 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U689 ( .A(KEYINPUT101), .B(KEYINPUT13), .Z(n593) );
  XNOR2_X1 U690 ( .A(KEYINPUT100), .B(G475), .ZN(n592) );
  XNOR2_X1 U691 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U692 ( .A(KEYINPUT95), .B(n748), .ZN(n639) );
  XNOR2_X2 U693 ( .A(n599), .B(KEYINPUT39), .ZN(n627) );
  NOR2_X1 U694 ( .A1(n600), .A2(n601), .ZN(n722) );
  NOR2_X1 U695 ( .A1(n720), .A2(n722), .ZN(n733) );
  NAND2_X1 U696 ( .A1(n733), .A2(KEYINPUT47), .ZN(n603) );
  XOR2_X1 U697 ( .A(KEYINPUT78), .B(n604), .Z(n611) );
  OR2_X1 U698 ( .A1(n720), .A2(n722), .ZN(n608) );
  INV_X1 U699 ( .A(KEYINPUT19), .ZN(n606) );
  NAND2_X1 U700 ( .A1(n608), .A2(n718), .ZN(n610) );
  INV_X1 U701 ( .A(KEYINPUT47), .ZN(n609) );
  INV_X1 U702 ( .A(KEYINPUT112), .ZN(n613) );
  INV_X1 U703 ( .A(n500), .ZN(n615) );
  XNOR2_X1 U704 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n616) );
  INV_X1 U705 ( .A(n746), .ZN(n650) );
  INV_X1 U706 ( .A(KEYINPUT113), .ZN(n617) );
  INV_X1 U707 ( .A(KEYINPUT48), .ZN(n618) );
  NAND2_X1 U708 ( .A1(n398), .A2(n736), .ZN(n619) );
  NOR2_X1 U709 ( .A1(n620), .A2(n619), .ZN(n622) );
  XNOR2_X1 U710 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n621) );
  XNOR2_X1 U711 ( .A(n622), .B(n621), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n624), .A2(n460), .ZN(n626) );
  INV_X1 U713 ( .A(KEYINPUT108), .ZN(n625) );
  XNOR2_X1 U714 ( .A(n626), .B(n625), .ZN(n810) );
  INV_X1 U715 ( .A(n810), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n627), .A2(n722), .ZN(n725) );
  AND2_X1 U717 ( .A1(n628), .A2(n725), .ZN(n629) );
  NOR2_X1 U718 ( .A1(G898), .A2(n630), .ZN(n631) );
  NOR2_X1 U719 ( .A1(n746), .A2(n745), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n635), .A2(n642), .ZN(n636) );
  INV_X1 U721 ( .A(KEYINPUT44), .ZN(n638) );
  NOR2_X1 U722 ( .A1(n746), .A2(n749), .ZN(n643) );
  INV_X1 U723 ( .A(n642), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n643), .A2(n659), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT77), .B(n644), .Z(n645) );
  NOR2_X1 U726 ( .A1(n655), .A2(n749), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n398), .A2(n647), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n463), .A2(n648), .ZN(n714) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n754) );
  NOR2_X1 U730 ( .A1(n499), .A2(n754), .ZN(n653) );
  XNOR2_X1 U731 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n723) );
  NOR2_X1 U733 ( .A1(n733), .A2(n656), .ZN(n658) );
  NOR2_X1 U734 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n657) );
  NOR2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n659), .A2(n398), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n662), .B(KEYINPUT84), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n663), .A2(n749), .ZN(n705) );
  AND2_X1 U739 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n665) );
  INV_X1 U740 ( .A(KEYINPUT45), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT81), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(KEYINPUT2), .ZN(n670) );
  INV_X1 U743 ( .A(n672), .ZN(n673) );
  INV_X1 U744 ( .A(KEYINPUT74), .ZN(n674) );
  INV_X1 U745 ( .A(n727), .ZN(n675) );
  INV_X1 U746 ( .A(KEYINPUT64), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n493), .A2(G210), .ZN(n684) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n682) );
  BUF_X1 U749 ( .A(n679), .Z(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(KEYINPUT79), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X2 U752 ( .A1(n685), .A2(n783), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n686), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U754 ( .A1(n770), .A2(G478), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X2 U756 ( .A1(n689), .A2(n783), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT122), .ZN(G63) );
  XOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .Z(n691) );
  NAND2_X1 U759 ( .A1(n770), .A2(G472), .ZN(n695) );
  XOR2_X1 U760 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n692) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X2 U762 ( .A1(n696), .A2(n783), .ZN(n698) );
  INV_X1 U763 ( .A(KEYINPUT63), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n698), .B(n697), .ZN(G57) );
  NAND2_X1 U765 ( .A1(n493), .A2(G475), .ZN(n702) );
  XNOR2_X1 U766 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X2 U768 ( .A1(n703), .A2(n783), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U770 ( .A(n705), .B(G101), .ZN(G3) );
  NAND2_X1 U771 ( .A1(n363), .A2(n361), .ZN(n706) );
  XNOR2_X1 U772 ( .A(n706), .B(KEYINPUT114), .ZN(n707) );
  XNOR2_X1 U773 ( .A(G104), .B(n707), .ZN(G6) );
  XOR2_X1 U774 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n709) );
  XNOR2_X1 U775 ( .A(G107), .B(KEYINPUT26), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n709), .B(n708), .ZN(n710) );
  XOR2_X1 U777 ( .A(KEYINPUT115), .B(n710), .Z(n713) );
  NAND2_X1 U778 ( .A1(n722), .A2(n363), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n713), .B(n712), .ZN(G9) );
  XOR2_X1 U780 ( .A(G110), .B(n714), .Z(G12) );
  XOR2_X1 U781 ( .A(G128), .B(KEYINPUT29), .Z(n716) );
  NAND2_X1 U782 ( .A1(n718), .A2(n722), .ZN(n715) );
  XNOR2_X1 U783 ( .A(n716), .B(n715), .ZN(G30) );
  XNOR2_X1 U784 ( .A(G143), .B(n717), .ZN(G45) );
  NAND2_X1 U785 ( .A1(n718), .A2(n361), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(G146), .ZN(G48) );
  NAND2_X1 U787 ( .A1(n723), .A2(n361), .ZN(n721) );
  XNOR2_X1 U788 ( .A(n721), .B(G113), .ZN(G15) );
  NAND2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U790 ( .A(n724), .B(G116), .ZN(G18) );
  XNOR2_X1 U791 ( .A(G134), .B(n725), .ZN(G36) );
  NOR2_X1 U792 ( .A1(n468), .A2(KEYINPUT2), .ZN(n726) );
  NOR2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U794 ( .A1(G953), .A2(n728), .ZN(n732) );
  INV_X1 U795 ( .A(n729), .ZN(n758) );
  AND2_X1 U796 ( .A1(n758), .A2(n743), .ZN(n730) );
  XNOR2_X1 U797 ( .A(n730), .B(KEYINPUT119), .ZN(n731) );
  NAND2_X1 U798 ( .A1(n732), .A2(n731), .ZN(n768) );
  NAND2_X1 U799 ( .A1(n608), .A2(n465), .ZN(n742) );
  INV_X1 U800 ( .A(n735), .ZN(n739) );
  NOR2_X1 U801 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U802 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U803 ( .A(KEYINPUT118), .B(n740), .Z(n741) );
  NAND2_X1 U804 ( .A1(n742), .A2(n741), .ZN(n744) );
  NAND2_X1 U805 ( .A1(n744), .A2(n743), .ZN(n761) );
  NAND2_X1 U806 ( .A1(n398), .A2(n745), .ZN(n747) );
  XOR2_X1 U807 ( .A(n747), .B(KEYINPUT50), .Z(n752) );
  NOR2_X1 U808 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U809 ( .A(KEYINPUT49), .B(n750), .Z(n751) );
  NOR2_X1 U810 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U811 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U812 ( .A(n756), .B(KEYINPUT51), .ZN(n757) );
  XNOR2_X1 U813 ( .A(n757), .B(KEYINPUT117), .ZN(n759) );
  NAND2_X1 U814 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U815 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U816 ( .A(KEYINPUT52), .B(n762), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U818 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U820 ( .A(KEYINPUT53), .B(n769), .ZN(G75) );
  BUF_X1 U821 ( .A(n493), .Z(n777) );
  NAND2_X1 U822 ( .A1(n777), .A2(G469), .ZN(n775) );
  XNOR2_X1 U823 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n771) );
  XNOR2_X1 U824 ( .A(n771), .B(KEYINPUT57), .ZN(n772) );
  XNOR2_X1 U825 ( .A(n773), .B(n772), .ZN(n774) );
  XNOR2_X1 U826 ( .A(n775), .B(n774), .ZN(n776) );
  NOR2_X1 U827 ( .A1(n783), .A2(n776), .ZN(G54) );
  NAND2_X1 U828 ( .A1(n777), .A2(G217), .ZN(n781) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(n780) );
  XNOR2_X1 U830 ( .A(n781), .B(n780), .ZN(n782) );
  NOR2_X1 U831 ( .A1(n783), .A2(n782), .ZN(G66) );
  NOR2_X1 U832 ( .A1(G898), .A2(n802), .ZN(n787) );
  XNOR2_X1 U833 ( .A(G101), .B(n784), .ZN(n785) );
  XNOR2_X1 U834 ( .A(n497), .B(n785), .ZN(n786) );
  NOR2_X1 U835 ( .A1(n787), .A2(n786), .ZN(n794) );
  NOR2_X1 U836 ( .A1(G953), .A2(n459), .ZN(n788) );
  XOR2_X1 U837 ( .A(KEYINPUT124), .B(n788), .Z(n792) );
  NAND2_X1 U838 ( .A1(G953), .A2(G224), .ZN(n789) );
  XNOR2_X1 U839 ( .A(KEYINPUT61), .B(n789), .ZN(n790) );
  NAND2_X1 U840 ( .A1(n790), .A2(G898), .ZN(n791) );
  NAND2_X1 U841 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U842 ( .A(n794), .B(n793), .Z(n795) );
  XNOR2_X1 U843 ( .A(KEYINPUT125), .B(n795), .ZN(G69) );
  XOR2_X1 U844 ( .A(n796), .B(KEYINPUT126), .Z(n800) );
  XNOR2_X1 U845 ( .A(n798), .B(n797), .ZN(n799) );
  XNOR2_X1 U846 ( .A(n800), .B(n799), .ZN(n804) );
  XNOR2_X1 U847 ( .A(n495), .B(n804), .ZN(n803) );
  NAND2_X1 U848 ( .A1(n803), .A2(n802), .ZN(n808) );
  XNOR2_X1 U849 ( .A(G227), .B(n804), .ZN(n805) );
  NAND2_X1 U850 ( .A1(n805), .A2(G900), .ZN(n806) );
  NAND2_X1 U851 ( .A1(n806), .A2(G953), .ZN(n807) );
  NAND2_X1 U852 ( .A1(n808), .A2(n807), .ZN(G72) );
  XOR2_X1 U853 ( .A(G122), .B(KEYINPUT127), .Z(n809) );
  XNOR2_X1 U854 ( .A(n501), .B(n809), .ZN(G24) );
  XOR2_X1 U855 ( .A(G140), .B(n810), .Z(G42) );
  XOR2_X1 U856 ( .A(G119), .B(n462), .Z(G21) );
  XOR2_X1 U857 ( .A(n496), .B(G137), .Z(G39) );
endmodule

