//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G250), .B1(G257), .B2(G264), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(KEYINPUT64), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(KEYINPUT64), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(new_n230));
  NAND4_X1  g0030(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n210), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n222), .B1(KEYINPUT0), .B2(new_n214), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT70), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n248), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(G226), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G97), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT76), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT76), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n257), .A2(new_n258), .A3(new_n262), .A4(new_n259), .ZN(new_n263));
  AND2_X1   g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n218), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT13), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n268), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n272), .B2(G238), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n266), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n267), .B1(new_n266), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g0075(.A(G169), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT77), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(G238), .ZN(new_n280));
  INV_X1    g0080(.A(new_n270), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(G1), .A2(G13), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n260), .B2(KEYINPUT76), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n282), .B1(new_n287), .B2(new_n263), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT77), .B1(new_n288), .B2(new_n267), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n267), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n279), .A2(new_n289), .A3(G179), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT14), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(G169), .C1(new_n274), .C2(new_n275), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n277), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n203), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT12), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(new_n218), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT73), .B1(new_n208), .B2(G1), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(new_n207), .A3(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n298), .B1(new_n203), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G20), .A2(G33), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n308), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n217), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(G77), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n299), .A2(new_n218), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT11), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n313), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n307), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n294), .A2(new_n317), .ZN(new_n318));
  AND4_X1   g0118(.A1(G190), .A2(new_n279), .A3(new_n289), .A4(new_n290), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n274), .B2(new_n275), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n316), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n270), .B1(new_n272), .B2(G232), .ZN(new_n323));
  OR2_X1    g0123(.A1(G223), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G226), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G1698), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n324), .B(new_n326), .C1(new_n255), .C2(new_n256), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G87), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n265), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n323), .A2(new_n330), .A3(G179), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n286), .A2(G232), .A3(new_n268), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n281), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n286), .B1(new_n327), .B2(new_n328), .ZN(new_n334));
  OAI21_X1  g0134(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n331), .A2(KEYINPUT79), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT79), .B1(new_n331), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n295), .A2(new_n340), .A3(new_n218), .A4(new_n299), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n305), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT8), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G58), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT71), .ZN(new_n346));
  OR3_X1    g0146(.A1(new_n344), .A2(KEYINPUT71), .A3(G58), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT78), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n295), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n300), .A2(KEYINPUT72), .B1(new_n304), .B2(new_n302), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n354), .B2(new_n341), .ZN(new_n355));
  INV_X1    g0155(.A(new_n352), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT78), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(G58), .B(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(G20), .B1(G159), .B2(new_n308), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT3), .B(G33), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT7), .B1(new_n360), .B2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G68), .ZN(new_n362));
  OR2_X1    g0162(.A1(KEYINPUT64), .A2(G20), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT64), .A2(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n365), .A2(new_n360), .A3(KEYINPUT7), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n359), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n313), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR4_X1   g0169(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT7), .A4(G20), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT7), .B1(new_n365), .B2(new_n360), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G68), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT16), .B1(new_n373), .B2(new_n359), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n353), .B(new_n357), .C1(new_n369), .C2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n338), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n338), .B2(new_n375), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n369), .A2(new_n374), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n323), .A2(new_n330), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G200), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n382), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n357), .A2(new_n353), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n381), .A2(new_n386), .A3(KEYINPUT17), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n375), .B2(new_n385), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n318), .A2(new_n322), .A3(new_n380), .A4(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n308), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n348), .B2(new_n310), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n313), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n354), .A2(G50), .A3(new_n341), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n296), .A2(new_n201), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT9), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n396), .A2(KEYINPUT9), .A3(new_n397), .A4(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n360), .A2(G222), .A3(new_n254), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n360), .A2(G223), .A3(G1698), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n255), .A2(new_n256), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G77), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n265), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n286), .A2(G226), .A3(new_n268), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n281), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G200), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n401), .A2(new_n402), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n407), .B2(new_n265), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n415), .A2(new_n416), .A3(G190), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n415), .B2(G190), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT10), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT74), .B1(new_n412), .B2(new_n384), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n415), .A2(new_n416), .A3(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT10), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n399), .A2(new_n400), .B1(new_n412), .B2(G200), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n402), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n412), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n399), .A3(new_n431), .ZN(new_n432));
  MUX2_X1   g0232(.A(new_n295), .B(new_n306), .S(G77), .Z(new_n433));
  NAND2_X1  g0233(.A1(new_n365), .A2(G77), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n343), .A2(new_n345), .ZN(new_n435));
  INV_X1    g0235(.A(new_n308), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n434), .B1(new_n435), .B2(new_n436), .C1(new_n310), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n313), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n360), .A2(G232), .A3(new_n254), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n360), .A2(G238), .A3(G1698), .ZN(new_n442));
  INV_X1    g0242(.A(G107), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n360), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n265), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n270), .B1(new_n272), .B2(G244), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n440), .B1(new_n448), .B2(G190), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(G200), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n447), .A2(G179), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n447), .A2(new_n428), .B1(new_n433), .B2(new_n439), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n449), .A2(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND4_X1   g0254(.A1(KEYINPUT75), .A2(new_n427), .A3(new_n432), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n432), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n420), .B2(new_n426), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT75), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n393), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G274), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n207), .A2(G45), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n207), .A3(G45), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(G250), .B1(new_n264), .B2(new_n218), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G238), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n472));
  OAI211_X1 g0272(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n265), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G200), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n207), .A2(G33), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n295), .A2(new_n479), .A3(new_n218), .A4(new_n299), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G87), .ZN(new_n484));
  OR2_X1    g0284(.A1(KEYINPUT83), .A2(G87), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT83), .A2(G87), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT19), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n259), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n365), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n363), .A2(G33), .A3(G97), .A4(new_n364), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n489), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n217), .A2(new_n360), .A3(G68), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n313), .B1(new_n296), .B2(new_n437), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n471), .A2(new_n476), .A3(G190), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n478), .A2(new_n484), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n313), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n437), .A2(new_n296), .ZN(new_n500));
  INV_X1    g0300(.A(new_n437), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n481), .A2(new_n501), .A3(new_n482), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n470), .B1(new_n265), .B2(new_n475), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n430), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n477), .A2(new_n428), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G250), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n509));
  OAI211_X1 g0309(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n510));
  INV_X1    g0310(.A(G294), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n284), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n265), .ZN(new_n513));
  OR2_X1    g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n464), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .A3(G274), .A4(new_n286), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  INV_X1    g0318(.A(new_n515), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n462), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G274), .B1(new_n264), .B2(new_n218), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n265), .B1(new_n462), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G264), .ZN(new_n527));
  AND4_X1   g0327(.A1(G190), .A2(new_n513), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G200), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n512), .A2(new_n265), .B1(new_n526), .B2(G264), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n524), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n474), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n208), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT23), .A2(G107), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n443), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n217), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n217), .A2(new_n360), .A3(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n217), .A2(new_n360), .A3(new_n541), .A4(G87), .ZN(new_n542));
  AOI211_X1 g0342(.A(KEYINPUT24), .B(new_n538), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n542), .ZN(new_n545));
  INV_X1    g0345(.A(new_n538), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n313), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n483), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n296), .A2(new_n443), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT25), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n532), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT7), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n217), .B2(new_n405), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n556), .A2(new_n370), .A3(new_n443), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n308), .A2(G77), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n443), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n558), .B1(new_n563), .B2(new_n217), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n313), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n481), .A2(G97), .A3(new_n482), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n295), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n360), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G283), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n360), .A2(G250), .A3(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n265), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n517), .A2(new_n523), .B1(new_n526), .B2(G257), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n428), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n430), .A3(new_n578), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n569), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(G200), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n371), .A2(G107), .A3(new_n372), .ZN(new_n584));
  AND2_X1   g0384(.A1(G97), .A2(G107), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n561), .B1(new_n585), .B2(new_n486), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n559), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n365), .B1(G77), .B2(new_n308), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n567), .B1(new_n589), .B2(new_n313), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n577), .A2(G190), .A3(new_n578), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n583), .A2(new_n590), .A3(new_n566), .A4(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n508), .A2(new_n554), .A3(new_n582), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT86), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n595));
  INV_X1    g0395(.A(new_n256), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT3), .A2(G33), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(G303), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G257), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n265), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n526), .A2(G270), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n524), .A2(new_n601), .A3(G190), .A4(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n301), .A2(KEYINPUT84), .A3(G116), .A4(new_n479), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT84), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n480), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n609), .A2(new_n610), .B1(new_n606), .B2(G20), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(new_n313), .ZN(new_n612));
  NAND2_X1  g0412(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n613));
  INV_X1    g0413(.A(G97), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n574), .B1(new_n614), .B2(G33), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(new_n613), .C1(new_n365), .C2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n313), .B(new_n611), .C1(new_n365), .C2(new_n615), .ZN(new_n617));
  INV_X1    g0417(.A(new_n613), .ZN(new_n618));
  INV_X1    g0418(.A(G13), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(G1), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n208), .A2(G116), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n617), .A2(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n603), .A2(new_n608), .A3(new_n616), .A4(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n517), .A2(new_n523), .B1(new_n526), .B2(G270), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n529), .B1(new_n624), .B2(new_n601), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n594), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n608), .A2(new_n622), .A3(new_n616), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n524), .A2(new_n601), .A3(new_n602), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n628), .A2(new_n630), .A3(KEYINPUT86), .A4(new_n603), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n627), .A2(KEYINPUT21), .A3(G169), .A4(new_n629), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n524), .A2(new_n601), .A3(new_n602), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n627), .A3(G179), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n428), .B1(new_n624), .B2(new_n601), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT21), .B1(new_n637), .B2(new_n627), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n530), .A2(new_n524), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n428), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n530), .A2(new_n430), .A3(new_n524), .ZN(new_n642));
  INV_X1    g0442(.A(new_n313), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n545), .A2(new_n546), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT24), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n545), .A2(new_n544), .A3(new_n546), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n549), .A2(new_n552), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n641), .B(new_n642), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n632), .A2(new_n639), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n460), .A2(new_n593), .A3(new_n650), .ZN(G372));
  NAND2_X1  g0451(.A1(new_n452), .A2(new_n453), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n319), .B2(new_n321), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n391), .B1(new_n318), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n331), .A2(new_n335), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n375), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(new_n376), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n427), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n432), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(KEYINPUT88), .A3(new_n432), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n569), .A2(new_n580), .A3(new_n581), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n508), .A2(new_n666), .A3(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n498), .A2(new_n507), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n582), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n641), .A2(new_n642), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n548), .B2(new_n553), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT87), .B1(new_n636), .B2(new_n638), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n637), .A2(new_n627), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT21), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT87), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n633), .A4(new_n635), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n673), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n671), .B(new_n507), .C1(new_n680), .C2(new_n593), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n665), .B1(new_n460), .B2(new_n682), .ZN(G369));
  NAND2_X1  g0483(.A1(new_n217), .A2(new_n620), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n647), .B2(new_n648), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n673), .B1(new_n554), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n689), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n673), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n639), .A2(new_n689), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n673), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n692), .A2(new_n628), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n674), .A2(new_n679), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n632), .A2(new_n639), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n693), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(G399));
  NOR2_X1   g0506(.A1(new_n212), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n488), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n220), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n579), .A2(new_n640), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n629), .A2(new_n477), .A3(new_n430), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n504), .A2(new_n530), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n430), .A3(new_n629), .ZN(new_n718));
  INV_X1    g0518(.A(new_n579), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT30), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT89), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n717), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n629), .A2(new_n430), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n719), .A3(new_n724), .A4(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n721), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n724), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n579), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n689), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n650), .A2(new_n593), .A3(new_n689), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n720), .A2(new_n716), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n734), .B(new_n692), .C1(new_n736), .C2(new_n725), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n713), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n639), .A2(new_n649), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n592), .A2(new_n582), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n508), .A4(new_n554), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n503), .A2(new_n505), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n667), .A2(new_n670), .B1(new_n506), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n740), .B1(new_n746), .B2(new_n692), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n681), .A2(new_n740), .A3(new_n692), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n739), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n712), .B1(new_n749), .B2(G1), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT90), .Z(G364));
  NOR2_X1   g0551(.A1(new_n365), .A2(new_n619), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G1), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n707), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n211), .A2(new_n360), .ZN(new_n756));
  XOR2_X1   g0556(.A(G355), .B(KEYINPUT91), .Z(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n211), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n248), .A2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n212), .A2(new_n360), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n461), .B2(new_n221), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n283), .B1(new_n208), .B2(G169), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n755), .B1(new_n763), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n217), .A2(new_n430), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n529), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G179), .A2(G200), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n365), .A2(new_n384), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n777), .A2(new_n201), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n774), .A2(new_n384), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n529), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(G68), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n217), .B1(G190), .B2(new_n779), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT93), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT93), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n614), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n529), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n365), .A2(new_n384), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n443), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n485), .A2(new_n487), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n793), .A2(G20), .A3(G190), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n360), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n784), .A2(G200), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n795), .B(new_n799), .C1(new_n800), .C2(G77), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n775), .A2(G200), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G58), .B1(new_n778), .B2(new_n782), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n786), .A2(new_n792), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT94), .B(G326), .Z(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G322), .A2(new_n802), .B1(new_n776), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G311), .A2(new_n800), .B1(new_n785), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n405), .B1(new_n798), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n780), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(G329), .ZN(new_n813));
  INV_X1    g0613(.A(new_n787), .ZN(new_n814));
  INV_X1    g0614(.A(new_n794), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(G294), .B1(new_n815), .B2(G283), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n807), .A2(new_n809), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n804), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n773), .B1(new_n818), .B2(new_n767), .ZN(new_n819));
  INV_X1    g0619(.A(new_n770), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n702), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n755), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n703), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n702), .A2(G330), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT95), .ZN(G396));
  NOR2_X1   g0626(.A1(new_n652), .A2(new_n689), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n449), .A2(new_n450), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n440), .A2(new_n689), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n827), .B1(new_n830), .B2(new_n652), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n674), .A2(new_n679), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n593), .B1(new_n832), .B2(new_n649), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT26), .B1(new_n508), .B2(new_n666), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n669), .A2(new_n582), .A3(new_n668), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n507), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n692), .B(new_n831), .C1(new_n833), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT97), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT97), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n681), .A2(new_n839), .A3(new_n692), .A4(new_n831), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n831), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n682), .B2(new_n689), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n739), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(new_n739), .A3(new_n843), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n755), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n776), .B1(new_n785), .B2(G150), .ZN(new_n849));
  INV_X1    g0649(.A(G143), .ZN(new_n850));
  INV_X1    g0650(.A(new_n802), .ZN(new_n851));
  INV_X1    g0651(.A(new_n800), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n849), .B1(new_n850), .B2(new_n851), .C1(new_n781), .C2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT34), .Z(new_n854));
  AOI21_X1  g0654(.A(new_n405), .B1(new_n812), .B2(G132), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT96), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n815), .A2(G68), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(new_n856), .ZN(new_n860));
  INV_X1    g0660(.A(new_n798), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n814), .A2(G58), .B1(new_n861), .B2(G50), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G283), .A2(new_n785), .B1(new_n776), .B2(G303), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n606), .B2(new_n852), .C1(new_n511), .C2(new_n851), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n815), .A2(G87), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n360), .B1(new_n861), .B2(G107), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n780), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n791), .A2(new_n869), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n854), .A2(new_n863), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n767), .A2(new_n768), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(new_n767), .B1(new_n311), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n831), .A2(new_n769), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n822), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT98), .B1(new_n848), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n847), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n739), .B1(new_n841), .B2(new_n843), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n822), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT98), .ZN(new_n881));
  INV_X1    g0681(.A(new_n876), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  NOR2_X1   g0685(.A1(new_n752), .A2(new_n207), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n318), .B(new_n322), .C1(new_n316), .C2(new_n692), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n294), .A2(new_n317), .A3(new_n689), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n827), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n841), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT100), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n841), .A2(KEYINPUT100), .A3(new_n891), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n381), .A2(new_n386), .A3(new_n387), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n367), .A2(new_n368), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n387), .B1(new_n369), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n656), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n900), .A2(new_n687), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n375), .A2(new_n385), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(new_n687), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n375), .B1(new_n338), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n338), .A2(new_n375), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT18), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n912), .A2(new_n390), .A3(new_n388), .A4(new_n377), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n913), .A2(KEYINPUT101), .A3(new_n903), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT101), .B1(new_n913), .B2(new_n903), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n910), .B(KEYINPUT38), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n896), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n897), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n375), .A2(new_n907), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n657), .A4(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .B1(new_n906), .B2(new_n908), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n658), .B2(new_n392), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n917), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n922), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n318), .A2(new_n689), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n935), .B1(new_n659), .B2(new_n687), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n921), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT103), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n459), .B(new_n938), .C1(new_n748), .C2(new_n747), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n459), .B1(new_n748), .B2(new_n747), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT103), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n665), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n937), .B(new_n942), .Z(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT40), .B1(new_n918), .B2(new_n919), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n692), .B1(new_n722), .B2(new_n730), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT31), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n842), .B1(new_n735), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n947), .A2(new_n889), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n919), .A2(new_n930), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n889), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT40), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n735), .A2(new_n946), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(new_n459), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n953), .A2(new_n955), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n957), .A2(new_n958), .A3(new_n713), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n886), .B1(new_n943), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n943), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n219), .A2(G116), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT35), .B2(new_n587), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT35), .B2(new_n587), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT36), .ZN(new_n966));
  OAI21_X1  g0766(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n967), .A2(new_n220), .B1(G50), .B2(new_n203), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(G1), .A3(new_n619), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT99), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n962), .A2(new_n971), .ZN(G367));
  AND2_X1   g0772(.A1(new_n484), .A2(new_n496), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n507), .A2(new_n973), .A3(new_n692), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n692), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n669), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT104), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n569), .A2(new_n689), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n742), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n666), .A2(new_n689), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n693), .A2(new_n694), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT105), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n582), .B1(new_n983), .B2(new_n649), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n988), .A2(KEYINPUT42), .B1(new_n692), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT42), .B2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(new_n985), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n705), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT106), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n994), .B1(new_n991), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n981), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OR3_X1    g0799(.A1(new_n997), .A2(new_n998), .A3(new_n981), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n707), .B(KEYINPUT41), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n698), .A2(new_n985), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT45), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n697), .A2(new_n992), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT44), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n705), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1003), .A2(new_n705), .A3(new_n1005), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n693), .B(new_n694), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(new_n704), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n749), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1001), .B1(new_n1015), .B2(new_n749), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n754), .B(KEYINPUT107), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n999), .B(new_n1000), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n767), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n790), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(G68), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n794), .A2(new_n311), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n405), .B(new_n1023), .C1(G58), .C2(new_n861), .ZN(new_n1024));
  INV_X1    g0824(.A(G137), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1022), .B(new_n1024), .C1(new_n1025), .C2(new_n780), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n785), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n201), .A2(new_n852), .B1(new_n1027), .B2(new_n781), .ZN(new_n1028));
  INV_X1    g0828(.A(G150), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n850), .A2(new_n777), .B1(new_n851), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n798), .A2(new_n606), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT46), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT108), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n777), .B2(new_n868), .C1(new_n810), .C2(new_n851), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n405), .B1(new_n1032), .B2(KEYINPUT46), .C1(new_n443), .C2(new_n787), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n815), .A2(G97), .ZN(new_n1037));
  INV_X1    g0837(.A(G317), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n780), .ZN(new_n1039));
  INV_X1    g0839(.A(G283), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1040), .A2(new_n852), .B1(new_n1027), .B2(new_n511), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1035), .A2(new_n1036), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1031), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1020), .B1(new_n1043), .B2(KEYINPUT47), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(KEYINPUT47), .B2(new_n1043), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n772), .B1(new_n212), .B2(new_n501), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n243), .A2(new_n760), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n822), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(new_n820), .C2(new_n976), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1019), .A2(new_n1049), .ZN(G387));
  NOR2_X1   g0850(.A1(new_n693), .A2(new_n820), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n709), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n1052), .C1(G68), .C2(G77), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT109), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n435), .A2(G50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n760), .C1(new_n461), .C2(new_n239), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(G107), .B2(new_n211), .C1(new_n709), .C2(new_n756), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n771), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n755), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1037), .B(new_n360), .C1(new_n311), .C2(new_n798), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G150), .B2(new_n812), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1021), .A2(new_n501), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G68), .A2(new_n800), .B1(new_n776), .B2(G159), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G50), .A2(new_n802), .B1(new_n785), .B2(new_n349), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n360), .B1(new_n815), .B2(G116), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G311), .A2(new_n785), .B1(new_n776), .B2(G322), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n810), .B2(new_n852), .C1(new_n1038), .C2(new_n851), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n814), .A2(G283), .B1(new_n861), .B2(G294), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1070), .B1(new_n780), .B2(new_n805), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1069), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1051), .B(new_n1063), .C1(new_n1081), .C2(new_n767), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1012), .A2(new_n749), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT110), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n707), .B(new_n1013), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  NOR2_X1   g0888(.A1(new_n252), .A2(new_n761), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n771), .B1(new_n614), .B2(new_n211), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n755), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G150), .A2(new_n776), .B1(new_n802), .B2(G159), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  AOI21_X1  g0893(.A(new_n405), .B1(new_n861), .B2(G68), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n866), .B(new_n1094), .C1(new_n850), .C2(new_n780), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n201), .A2(new_n1027), .B1(new_n852), .B2(new_n435), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G77), .C2(new_n1021), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n360), .B(new_n795), .C1(G116), .C2(new_n814), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n511), .B2(new_n852), .C1(new_n810), .C2(new_n1027), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n812), .A2(G322), .B1(G283), .B2(new_n861), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT111), .Z(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G311), .A2(new_n802), .B1(new_n776), .B2(G317), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT52), .Z(new_n1104));
  AOI22_X1  g0904(.A1(new_n1093), .A2(new_n1097), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT112), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1020), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1091), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n820), .B2(new_n985), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1010), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n1017), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n708), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1013), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(G390));
  NAND3_X1  g0916(.A1(new_n954), .A2(new_n459), .A3(G330), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n665), .A2(new_n939), .A3(new_n941), .A4(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n632), .A2(new_n639), .A3(new_n649), .ZN(new_n1119));
  AND4_X1   g0919(.A1(new_n582), .A2(new_n508), .A3(new_n554), .A4(new_n592), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n692), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n945), .B1(new_n1121), .B2(KEYINPUT31), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n831), .C1(new_n1122), .C2(new_n737), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n890), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n954), .A2(G330), .A3(new_n831), .A4(new_n889), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT100), .B1(new_n841), .B2(new_n891), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n893), .B(new_n827), .C1(new_n838), .C2(new_n840), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n739), .A2(new_n831), .A3(new_n889), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n689), .B1(new_n743), .B2(new_n745), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n830), .A2(new_n652), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n827), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n947), .A2(G330), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1130), .B(new_n1133), .C1(new_n1134), .C2(new_n889), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1118), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n934), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n896), .B2(new_n935), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1133), .A2(new_n890), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n935), .B(KEYINPUT113), .Z(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n931), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n889), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n935), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n934), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1130), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1142), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1137), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1139), .A2(new_n1130), .A3(new_n1142), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1125), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1153), .A3(new_n1136), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n707), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n1018), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n790), .A2(new_n311), .B1(new_n851), .B2(new_n606), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT114), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n360), .B1(new_n861), .B2(G87), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n859), .B(new_n1159), .C1(new_n511), .C2(new_n780), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G97), .A2(new_n800), .B1(new_n785), .B2(G107), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1040), .B2(new_n777), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1158), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  AOI22_X1  g0964(.A1(G132), .A2(new_n802), .B1(new_n800), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n360), .B1(new_n780), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n861), .A2(G150), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G50), .C2(new_n815), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G128), .A2(new_n776), .B1(new_n785), .B2(G137), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1021), .A2(G159), .ZN(new_n1172));
  AND4_X1   g0972(.A1(new_n1165), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n767), .B1(new_n1163), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n822), .B1(new_n348), .B2(new_n872), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n934), .C2(new_n769), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1156), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1155), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT115), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1155), .A2(new_n1177), .A3(KEYINPUT115), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G378));
  INV_X1    g0983(.A(KEYINPUT118), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n931), .A2(new_n889), .A3(new_n947), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(KEYINPUT40), .A2(new_n1185), .B1(new_n944), .B2(new_n948), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1186), .B2(new_n713), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n953), .A2(KEYINPUT118), .A3(G330), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n399), .A2(new_n907), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n457), .B(new_n1189), .Z(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1187), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1192), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n953), .A2(KEYINPUT118), .A3(G330), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n937), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1193), .A2(new_n937), .A3(new_n1195), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1018), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n872), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n755), .B1(new_n1201), .B2(G50), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G50), .B1(new_n597), .B2(new_n285), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G41), .B(new_n360), .C1(new_n861), .C2(G77), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n815), .A2(G58), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1040), .C2(new_n780), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n614), .A2(new_n1027), .B1(new_n852), .B2(new_n437), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G107), .C2(new_n802), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1022), .B1(new_n606), .B2(new_n777), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT116), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(KEYINPUT116), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1203), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G132), .A2(new_n785), .B1(new_n800), .B2(G137), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1166), .B2(new_n777), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n802), .A2(G128), .B1(new_n861), .B2(new_n1164), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT117), .Z(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G150), .C2(new_n1021), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n815), .A2(G159), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n812), .C2(G124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1214), .B1(new_n1213), .B2(new_n1212), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1202), .B1(new_n1226), .B2(new_n767), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n769), .B2(new_n1192), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1200), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1118), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1154), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1232), .A2(KEYINPUT57), .A3(new_n1199), .A4(new_n1198), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n707), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1193), .A2(new_n937), .A3(new_n1195), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n937), .B1(new_n1195), .B2(new_n1193), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1232), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1230), .B1(new_n1234), .B2(new_n1238), .ZN(G375));
  INV_X1    g1039(.A(new_n1001), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1129), .A2(new_n1118), .A3(new_n1135), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1137), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n890), .A2(new_n768), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n755), .B1(new_n1201), .B2(G68), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n360), .B(new_n1023), .C1(G97), .C2(new_n861), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1066), .B(new_n1245), .C1(new_n810), .C2(new_n780), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G116), .A2(new_n785), .B1(new_n776), .B2(G294), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n443), .B2(new_n852), .C1(new_n1040), .C2(new_n851), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1021), .A2(G50), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n812), .A2(G128), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n405), .B1(new_n861), .B2(G159), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1249), .A2(new_n1205), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G132), .A2(new_n776), .B1(new_n800), .B2(G150), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G137), .A2(new_n802), .B1(new_n785), .B2(new_n1164), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1246), .A2(new_n1248), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1244), .B1(new_n1256), .B2(new_n767), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1243), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1133), .B1(new_n1123), .B2(new_n890), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n889), .B1(new_n947), .B2(G330), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n894), .A2(new_n895), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n1126), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1258), .B1(new_n1263), .B2(new_n1017), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1242), .A2(new_n1265), .ZN(G381));
  NAND3_X1  g1066(.A1(new_n1019), .A2(new_n1049), .A3(new_n1115), .ZN(new_n1267));
  OR2_X1    g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1267), .A2(G384), .A3(G381), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1178), .ZN(new_n1270));
  INV_X1    g1070(.A(G375), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(G407));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1270), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G407), .B(G213), .C1(G343), .C2(new_n1273), .ZN(G409));
  INV_X1    g1074(.A(new_n1232), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1001), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1270), .B1(new_n1277), .B2(new_n1229), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(G375), .B2(new_n1182), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n688), .A2(G213), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1241), .B1(new_n1136), .B2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1129), .A2(new_n1118), .A3(KEYINPUT60), .A4(new_n1135), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1283), .A2(new_n707), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n884), .B(new_n1264), .C1(new_n1282), .C2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G384), .B1(new_n1286), .B2(new_n1265), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1279), .A2(new_n1280), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT123), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1268), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1019), .A2(new_n1049), .A3(new_n1115), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1115), .B1(new_n1019), .B2(new_n1049), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1291), .B(new_n1295), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(G390), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1295), .A2(new_n1291), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT123), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1299), .A2(new_n1267), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1298), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1279), .A2(new_n1304), .A3(new_n1280), .A4(new_n1288), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1290), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  XOR2_X1   g1106(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1307));
  NAND3_X1  g1107(.A1(new_n688), .A2(G213), .A3(G2897), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT120), .B1(new_n1288), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1283), .A2(new_n707), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT60), .B1(new_n1263), .B2(new_n1118), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1311), .B2(new_n1241), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n884), .B1(new_n1312), .B2(new_n1264), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1286), .A2(G384), .A3(new_n1265), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1308), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT120), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1308), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT121), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT121), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1321), .B(new_n1308), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1322));
  OAI22_X1  g1122(.A1(new_n1309), .A2(new_n1317), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT122), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1315), .B(new_n1316), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1288), .B2(new_n1308), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1318), .A2(KEYINPUT121), .A3(new_n1319), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT122), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT57), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1332), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(new_n707), .A3(new_n1233), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1334), .A2(new_n1180), .A3(new_n1181), .A4(new_n1230), .ZN(new_n1335));
  AOI22_X1  g1135(.A1(new_n1335), .A2(new_n1278), .B1(G213), .B2(new_n688), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1307), .B1(new_n1331), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT125), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  OAI211_X1 g1139(.A(KEYINPUT125), .B(new_n1307), .C1(new_n1331), .C2(new_n1336), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1306), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1289), .A2(KEYINPUT63), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1279), .A2(new_n1343), .A3(new_n1280), .A4(new_n1288), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT61), .B1(new_n1342), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(KEYINPUT119), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT119), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1279), .A2(new_n1348), .A3(new_n1280), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1347), .A2(new_n1349), .A3(new_n1330), .A4(new_n1324), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1303), .B1(new_n1345), .B2(new_n1350), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1341), .A2(new_n1351), .ZN(G405));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1270), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1335), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1288), .B1(new_n1354), .B2(KEYINPUT126), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1355), .B1(KEYINPUT126), .B2(new_n1354), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1303), .ZN(new_n1357));
  OR3_X1    g1157(.A1(new_n1354), .A2(KEYINPUT126), .A3(new_n1318), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1356), .A2(new_n1357), .A3(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1357), .B1(new_n1356), .B2(new_n1358), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(G402));
endmodule


