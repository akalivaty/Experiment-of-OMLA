//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n211), .B1(KEYINPUT1), .B2(new_n221), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n221), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G222), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n255), .B1(new_n202), .B2(new_n253), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n226), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(G274), .B1(new_n259), .B2(new_n260), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT68), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(new_n226), .B2(new_n263), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  INV_X1    g0072(.A(new_n268), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n268), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G226), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n266), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G179), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n279), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n260), .ZN(new_n284));
  XOR2_X1   g0084(.A(KEYINPUT8), .B(G58), .Z(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n225), .A2(new_n250), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(new_n206), .A3(new_n250), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n206), .B2(new_n201), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n284), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(G50), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n206), .A2(G1), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n284), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  XOR2_X1   g0107(.A(new_n307), .B(KEYINPUT73), .Z(new_n308));
  NAND2_X1  g0108(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n282), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n279), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G200), .B2(new_n279), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT9), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n301), .B2(new_n308), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n314), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n314), .C1(new_n315), .C2(new_n317), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n311), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n302), .B1(new_n286), .B2(new_n289), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n286), .A2(new_n289), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n306), .ZN(new_n325));
  XNOR2_X1  g0125(.A(G58), .B(G68), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n295), .A2(G159), .B1(new_n326), .B2(G20), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n328), .A2(new_n329), .A3(G20), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  OAI21_X1  g0131(.A(G68), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n251), .A2(new_n222), .A3(new_n224), .A4(new_n252), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(KEYINPUT7), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT16), .B(new_n327), .C1(new_n332), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n284), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(KEYINPUT7), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(new_n331), .A3(new_n206), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G68), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT16), .B1(new_n340), .B2(new_n327), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n325), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n276), .A2(G232), .A3(new_n268), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G223), .A2(G1698), .ZN(new_n345));
  INV_X1    g0145(.A(G226), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(G1698), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n253), .B1(G33), .B2(G87), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n226), .A2(new_n262), .A3(new_n263), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n344), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n267), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n281), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n346), .A2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G223), .B2(G1698), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n359), .A2(new_n338), .B1(new_n250), .B2(new_n215), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n343), .B1(new_n360), .B2(new_n265), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(new_n275), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n356), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n356), .B2(new_n363), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT76), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT76), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n265), .ZN(new_n368));
  AND4_X1   g0168(.A1(new_n362), .A2(new_n368), .A3(new_n275), .A4(new_n344), .ZN(new_n369));
  AOI21_X1  g0169(.A(G169), .B1(new_n361), .B2(new_n275), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT75), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n356), .A2(new_n357), .A3(new_n363), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n342), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT18), .ZN(new_n375));
  INV_X1    g0175(.A(new_n342), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT76), .B1(new_n364), .B2(new_n365), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n372), .A3(new_n367), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n352), .B2(new_n355), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n361), .A2(G190), .A3(new_n275), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n382), .B1(new_n342), .B2(new_n385), .ZN(new_n386));
  AND4_X1   g0186(.A1(G190), .A2(new_n368), .A3(new_n275), .A4(new_n344), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n361), .B2(new_n275), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT64), .B(G20), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n331), .B1(new_n338), .B2(new_n392), .ZN(new_n393));
  NOR4_X1   g0193(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT7), .A4(G20), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n393), .A2(new_n394), .A3(new_n213), .ZN(new_n395));
  INV_X1    g0195(.A(new_n327), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n284), .A3(new_n335), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n390), .A2(KEYINPUT17), .A3(new_n398), .A4(new_n325), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n375), .A2(new_n381), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n253), .A2(G232), .A3(new_n254), .ZN(new_n403));
  INV_X1    g0203(.A(G107), .ZN(new_n404));
  OAI221_X1 g0204(.A(new_n403), .B1(new_n404), .B2(new_n253), .C1(new_n256), .C2(new_n214), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n265), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n277), .A2(G244), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n406), .A2(new_n275), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n362), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT15), .B(G87), .Z(new_n410));
  NAND2_X1  g0210(.A1(new_n290), .A2(new_n410), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n411), .B1(new_n202), .B2(new_n392), .C1(new_n296), .C2(new_n287), .ZN(new_n412));
  INV_X1    g0212(.A(new_n302), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n412), .A2(new_n284), .B1(new_n202), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n413), .B2(new_n284), .ZN(new_n416));
  INV_X1    g0216(.A(new_n305), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n302), .A2(KEYINPUT74), .A3(new_n260), .A4(new_n283), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G77), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n406), .A2(new_n275), .A3(new_n407), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n281), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n409), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n408), .A2(G190), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(G200), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n420), .A3(new_n414), .A4(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n276), .A2(G238), .A3(new_n268), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n269), .B2(new_n274), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  OAI211_X1 g0232(.A(G232), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n433));
  OAI211_X1 g0233(.A(G226), .B(new_n254), .C1(new_n328), .C2(new_n329), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n265), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n432), .B1(new_n431), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(G169), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n431), .A2(new_n437), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT13), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(G179), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(G169), .C1(new_n438), .C2(new_n439), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n284), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n392), .A2(G33), .A3(G77), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT11), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n419), .A2(G68), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n413), .A2(new_n213), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT12), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n452), .B2(KEYINPUT11), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n448), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(G200), .B1(new_n438), .B2(new_n439), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n443), .A2(G190), .A3(new_n444), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n429), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n322), .A2(new_n402), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT21), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n205), .B2(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n416), .A2(new_n418), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n413), .A2(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n250), .A2(G97), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n222), .A2(new_n224), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n283), .A2(new_n260), .B1(G20), .B2(new_n469), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n475), .A2(KEYINPUT20), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT20), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n471), .B(new_n472), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G169), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n271), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n276), .ZN(new_n488));
  INV_X1    g0288(.A(G270), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(G264), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n491));
  OAI211_X1 g0291(.A(G257), .B(new_n254), .C1(new_n328), .C2(new_n329), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n251), .A2(G303), .A3(new_n252), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n351), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT77), .A4(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n468), .B1(new_n480), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT78), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT78), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n468), .C1(new_n480), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n480), .A2(new_n498), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n362), .B(new_n490), .C1(new_n496), .C2(new_n497), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(KEYINPUT21), .B1(new_n479), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n498), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n479), .B1(new_n508), .B2(G200), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n312), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n487), .A2(G257), .A3(new_n276), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n484), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(new_n254), .C1(new_n328), .C2(new_n329), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n474), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n519), .B2(new_n265), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n393), .A2(new_n394), .A3(new_n404), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n202), .B1(new_n293), .B2(new_n294), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n404), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G97), .B(G107), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n525), .B1(new_n529), .B2(new_n392), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n284), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n302), .A2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n205), .A2(G33), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n302), .A2(new_n533), .A3(new_n260), .A4(new_n283), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(G97), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n531), .B(new_n536), .C1(new_n520), .C2(new_n388), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n337), .A2(G107), .A3(new_n339), .ZN(new_n538));
  AND2_X1   g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n528), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n404), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n524), .B1(new_n543), .B2(new_n225), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n449), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n536), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n520), .A2(G169), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(G179), .B(new_n513), .C1(new_n519), .C2(new_n265), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n522), .A2(new_n537), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n410), .A2(new_n302), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n222), .A2(new_n224), .A3(G33), .A4(G97), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n253), .A2(new_n392), .A3(G68), .ZN(new_n554));
  NAND3_X1  g0354(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n222), .A2(new_n224), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n540), .A2(new_n215), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n550), .B1(new_n559), .B2(new_n284), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n535), .A2(new_n410), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n271), .A2(new_n482), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n276), .B(G250), .C1(G1), .C2(new_n481), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G238), .B(new_n254), .C1(new_n328), .C2(new_n329), .ZN(new_n566));
  OAI211_X1 g0366(.A(G244), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n265), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n362), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n265), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n563), .A2(new_n564), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n281), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n562), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n534), .A2(new_n215), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n550), .B(new_n577), .C1(new_n559), .C2(new_n284), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n570), .A2(G190), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n549), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n487), .A2(G264), .A3(new_n276), .ZN(new_n584));
  INV_X1    g0384(.A(G294), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n250), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G250), .A2(G1698), .ZN(new_n587));
  INV_X1    g0387(.A(G257), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n589), .B2(new_n253), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n484), .B(new_n584), .C1(new_n590), .C2(new_n351), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n312), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT82), .B1(new_n591), .B2(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n388), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n413), .A2(new_n404), .ZN(new_n598));
  NOR2_X1   g0398(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n600), .A2(new_n602), .B1(G107), .B2(new_n535), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n206), .ZN(new_n606));
  NAND2_X1  g0406(.A1(KEYINPUT23), .A2(G107), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n404), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n607), .C1(new_n392), .C2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n222), .B(new_n224), .C1(new_n328), .C2(new_n329), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT22), .B1(new_n610), .B2(new_n215), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT22), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n253), .A2(new_n392), .A3(new_n612), .A4(G87), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n284), .B1(new_n614), .B2(KEYINPUT24), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT24), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n616), .B(new_n609), .C1(new_n611), .C2(new_n613), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n603), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n597), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n591), .A2(G169), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n588), .A2(G1698), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G250), .B2(G1698), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n622), .A2(new_n338), .B1(new_n250), .B2(new_n585), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n265), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(G179), .A3(new_n484), .A4(new_n584), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT80), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n620), .A2(KEYINPUT80), .A3(new_n625), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n618), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT81), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n618), .A2(new_n628), .A3(KEYINPUT81), .A4(new_n629), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n583), .A2(new_n619), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n467), .A2(new_n511), .A3(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n467), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n618), .A2(new_n626), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n503), .A2(new_n506), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT84), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n503), .A2(new_n640), .A3(new_n506), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n531), .A2(new_n536), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n520), .A2(new_n362), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n642), .B(new_n643), .C1(G169), .C2(new_n520), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n545), .A2(new_n546), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n645), .B(new_n521), .C1(new_n388), .C2(new_n520), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n644), .B(new_n646), .C1(new_n597), .C2(new_n618), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT83), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n569), .A2(new_n648), .A3(new_n265), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n569), .B2(new_n265), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n573), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n281), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n560), .A2(new_n561), .B1(new_n570), .B2(new_n362), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n572), .A2(KEYINPUT83), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n569), .A2(new_n648), .A3(new_n265), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n565), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n579), .B(new_n578), .C1(new_n657), .C2(new_n388), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n647), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n639), .A2(new_n641), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n659), .B2(new_n644), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT85), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n662), .C1(new_n659), .C2(new_n644), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n519), .A2(new_n265), .ZN(new_n667));
  INV_X1    g0467(.A(new_n513), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n669), .A2(new_n281), .B1(new_n531), .B2(new_n536), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n576), .A3(new_n581), .A4(new_n643), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n664), .A2(new_n666), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n661), .A2(new_n674), .A3(new_n654), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n636), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n386), .A2(new_n399), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n465), .A2(new_n424), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n461), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n380), .B(new_n342), .C1(new_n364), .C2(new_n365), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n371), .A2(new_n372), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n380), .B1(new_n683), .B2(new_n342), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n680), .A2(KEYINPUT87), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n319), .A2(new_n321), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT87), .B1(new_n680), .B2(new_n686), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n310), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n677), .A2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(G13), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n392), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n392), .A2(new_n698), .A3(new_n695), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n479), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n507), .A2(new_n510), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n507), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n632), .A2(new_n633), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n619), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n618), .A2(new_n702), .ZN(new_n710));
  INV_X1    g0510(.A(new_n702), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n709), .A2(new_n710), .B1(new_n630), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n507), .A2(new_n702), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n619), .A3(new_n708), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n618), .A2(new_n626), .A3(new_n711), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n209), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n205), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n557), .A2(G116), .ZN(new_n722));
  INV_X1    g0522(.A(new_n228), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n721), .A2(new_n722), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n498), .A2(G179), .ZN(new_n727));
  INV_X1    g0527(.A(new_n488), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(G264), .B1(new_n623), .B2(new_n265), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n520), .A2(new_n729), .A3(new_n570), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n570), .A2(new_n729), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n505), .A2(new_n732), .A3(KEYINPUT30), .A4(new_n520), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n592), .A2(G179), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n508), .A2(new_n734), .A3(new_n669), .A4(new_n651), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n702), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n702), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n503), .A2(new_n510), .A3(new_n506), .A4(new_n711), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n739), .B(new_n740), .C1(new_n634), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n675), .A2(new_n711), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(KEYINPUT88), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT88), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n675), .B2(new_n711), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n745), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n632), .A2(new_n503), .A3(new_n506), .A4(new_n633), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n660), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n578), .A2(new_n579), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n651), .A2(G200), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(new_n652), .B2(new_n653), .ZN(new_n755));
  INV_X1    g0555(.A(new_n644), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n662), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n654), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n702), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT29), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n744), .B1(new_n750), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n725), .B1(new_n762), .B2(G1), .ZN(G364));
  NOR2_X1   g0563(.A1(new_n225), .A2(new_n694), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT89), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n721), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n705), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n260), .B1(G20), .B2(new_n281), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n719), .A2(new_n253), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n481), .B2(new_n723), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n244), .B2(new_n481), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n209), .A2(new_n253), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT90), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G355), .B1(new_n469), .B2(new_n719), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n775), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n392), .A2(new_n362), .A3(new_n312), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  INV_X1    g0585(.A(G326), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n392), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n388), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n785), .A2(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n788), .A2(G20), .A3(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n253), .B1(new_n793), .B2(G303), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n225), .B1(new_n312), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n799), .A2(new_n362), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n794), .B1(new_n798), .B2(new_n585), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n799), .A2(new_n796), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n791), .B(new_n803), .C1(G329), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n784), .A2(new_n388), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT91), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(KEYINPUT91), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G322), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n787), .A2(G179), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT93), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n814), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT33), .B(G317), .Z(new_n819));
  OAI211_X1 g0619(.A(new_n805), .B(new_n812), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n785), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n800), .A2(G77), .B1(new_n821), .B2(G50), .ZN(new_n822));
  INV_X1    g0622(.A(G58), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n810), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT92), .Z(new_n825));
  NAND2_X1  g0625(.A1(new_n804), .A2(G159), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT32), .Z(new_n827));
  NOR2_X1   g0627(.A1(new_n792), .A2(new_n215), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G97), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n253), .C1(new_n798), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n789), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(G107), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n827), .B(new_n833), .C1(new_n213), .C2(new_n818), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n820), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n783), .B1(new_n835), .B2(new_n773), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n767), .B1(new_n772), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n767), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n705), .A2(G330), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(new_n706), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT94), .ZN(G396));
  NOR2_X1   g0642(.A1(new_n425), .A2(new_n702), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n421), .A2(new_n702), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n424), .B1(new_n428), .B2(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n747), .A2(new_n749), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n429), .A2(new_n711), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n675), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n846), .A2(new_n744), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT97), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n846), .A2(new_n849), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n767), .C1(new_n744), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n773), .A2(new_n768), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n767), .B1(new_n202), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n843), .A2(new_n845), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n810), .A2(new_n585), .B1(new_n830), .B2(new_n798), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT95), .Z(new_n859));
  AOI22_X1  g0659(.A1(G311), .A2(new_n804), .B1(new_n832), .B2(G87), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n338), .B1(new_n792), .B2(new_n404), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n821), .B2(G303), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(new_n469), .C2(new_n801), .ZN(new_n863));
  INV_X1    g0663(.A(new_n818), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(G283), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n800), .A2(G159), .B1(new_n821), .B2(G137), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n818), .B2(new_n297), .C1(new_n868), .C2(new_n810), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n832), .A2(G68), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n338), .B1(new_n793), .B2(G50), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n804), .A2(G132), .B1(G58), .B2(new_n797), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n866), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT96), .ZN(new_n878));
  INV_X1    g0678(.A(new_n773), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n856), .B1(new_n769), .B2(new_n857), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n854), .A2(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n765), .A2(new_n205), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n327), .B1(new_n332), .B2(new_n334), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(new_n391), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n325), .B1(new_n884), .B2(new_n336), .ZN(new_n885));
  INV_X1    g0685(.A(new_n700), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n400), .B1(new_n379), .B2(new_n380), .ZN(new_n889));
  AOI211_X1 g0689(.A(KEYINPUT18), .B(new_n376), .C1(new_n377), .C2(new_n378), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n390), .A2(new_n398), .A3(new_n325), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n700), .B(KEYINPUT100), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n342), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n374), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n376), .A2(new_n390), .B1(new_n885), .B2(new_n886), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n683), .A2(new_n885), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n891), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n374), .A2(new_n898), .B1(new_n902), .B2(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n401), .B2(new_n888), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n459), .A2(new_n711), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n448), .B2(new_n464), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT99), .ZN(new_n911));
  INV_X1    g0711(.A(new_n909), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n461), .A2(new_n465), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT99), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n909), .C1(new_n448), .C2(new_n464), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n742), .A2(new_n916), .A3(new_n857), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT40), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n895), .B1(new_n685), .B2(new_n400), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n342), .B1(new_n364), .B2(new_n365), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n893), .A3(new_n895), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n374), .A2(new_n898), .B1(new_n922), .B2(KEYINPUT37), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n892), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n919), .B1(new_n905), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n918), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n636), .A2(new_n742), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(G330), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n930), .A2(KEYINPUT102), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(KEYINPUT102), .B2(new_n930), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n663), .A2(KEYINPUT85), .B1(KEYINPUT26), .B2(new_n672), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(new_n666), .B1(new_n653), .B2(new_n652), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n847), .B1(new_n934), .B2(new_n661), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n916), .B1(new_n935), .B2(new_n843), .ZN(new_n936));
  INV_X1    g0736(.A(new_n906), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n891), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n377), .A2(new_n378), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n897), .B1(new_n939), .B2(new_n342), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT38), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n401), .B2(new_n888), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n936), .A2(new_n944), .B1(new_n685), .B2(new_n894), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n448), .A2(new_n460), .A3(new_n711), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT39), .B1(new_n938), .B2(new_n943), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT101), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  AND4_X1   g0750(.A1(new_n949), .A2(new_n905), .A3(new_n950), .A4(new_n924), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n921), .A2(KEYINPUT18), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n400), .A2(new_n952), .A3(new_n681), .ZN(new_n953));
  INV_X1    g0753(.A(new_n895), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n893), .A2(new_n895), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n371), .A2(new_n372), .B1(new_n398), .B2(new_n325), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT37), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n379), .B2(new_n897), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT39), .B1(new_n960), .B2(new_n892), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n949), .B1(new_n961), .B2(new_n905), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n948), .B1(new_n951), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n945), .B1(new_n947), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n467), .B1(KEYINPUT29), .B2(new_n760), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n691), .B1(new_n750), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n882), .B1(new_n932), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n932), .ZN(new_n969));
  OAI21_X1  g0769(.A(G77), .B1(new_n823), .B2(new_n213), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n970), .A2(new_n228), .B1(G50), .B2(new_n213), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(G1), .A3(new_n694), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT98), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n469), .B(new_n227), .C1(KEYINPUT35), .C2(new_n543), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(KEYINPUT35), .B2(new_n543), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT36), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n969), .A2(new_n978), .ZN(G367));
  OR2_X1    g0779(.A1(new_n235), .A2(new_n777), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n775), .B1(new_n719), .B2(new_n410), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n767), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n755), .B1(new_n578), .B2(new_n711), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n654), .A2(new_n578), .A3(new_n711), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n789), .A2(new_n830), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n785), .A2(new_n802), .B1(new_n798), .B2(new_n404), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(G317), .C2(new_n804), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n792), .A2(new_n469), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n253), .B(new_n990), .C1(G283), .C2(new_n800), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G303), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n585), .B2(new_n818), .C1(new_n993), .C2(new_n810), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT105), .ZN(new_n995));
  INV_X1    g0795(.A(new_n804), .ZN(new_n996));
  INV_X1    g0796(.A(G137), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(new_n823), .B2(new_n792), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n811), .A2(G150), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n995), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n864), .A2(G159), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n253), .B1(new_n798), .B2(new_n213), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n785), .A2(new_n868), .B1(new_n789), .B2(new_n202), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(G50), .C2(new_n800), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n994), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  OAI221_X1 g0807(.A(new_n982), .B1(new_n771), .B2(new_n985), .C1(new_n1007), .C2(new_n879), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n766), .A2(G1), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n756), .A2(new_n702), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n644), .B(new_n646), .C1(new_n645), .C2(new_n711), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n717), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT45), .Z(new_n1014));
  NOR3_X1   g0814(.A1(new_n717), .A2(KEYINPUT103), .A3(new_n1012), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT44), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT103), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n715), .A2(new_n716), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1012), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OR3_X1    g0820(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1016), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1014), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT104), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n713), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n715), .B1(new_n712), .B2(new_n714), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n707), .B(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n762), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1023), .A2(KEYINPUT104), .A3(new_n707), .A4(new_n712), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n762), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n720), .B(KEYINPUT41), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1009), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n715), .A2(new_n1019), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT42), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n644), .B1(new_n708), .B2(new_n1011), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1035), .A2(KEYINPUT42), .B1(new_n711), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(new_n1038), .B1(KEYINPUT43), .B2(new_n985), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n713), .A2(new_n1019), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1008), .B1(new_n1034), .B2(new_n1043), .ZN(G387));
  OR2_X1    g0844(.A1(new_n712), .A2(new_n771), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n776), .B1(new_n240), .B2(new_n481), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n781), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n722), .B2(new_n1047), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n287), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n287), .B2(G50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n722), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1048), .A2(new_n1052), .B1(new_n404), .B2(new_n719), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n838), .B1(new_n1053), .B2(new_n775), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n864), .A2(new_n324), .B1(G68), .B2(new_n800), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT107), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n986), .A2(new_n338), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n797), .A2(new_n410), .ZN(new_n1058));
  INV_X1    g0858(.A(G159), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(new_n785), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G50), .B2(new_n811), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n804), .A2(G150), .B1(G77), .B2(new_n793), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT106), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1056), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n253), .B1(new_n804), .B2(G326), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n798), .A2(new_n790), .B1(new_n585), .B2(new_n792), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n800), .A2(G303), .B1(new_n821), .B2(G322), .ZN(new_n1067));
  INV_X1    g0867(.A(G317), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n818), .B2(new_n802), .C1(new_n1068), .C2(new_n810), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1065), .B1(new_n469), .B2(new_n789), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1054), .B1(new_n1076), .B2(new_n773), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1027), .A2(new_n1009), .B1(new_n1045), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1028), .A2(new_n720), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n762), .A2(new_n1027), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  XNOR2_X1  g0881(.A(new_n1023), .B(new_n713), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1031), .B(new_n720), .C1(new_n1029), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1019), .A2(new_n770), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT108), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n810), .A2(new_n1059), .B1(new_n297), .B2(new_n785), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  OAI22_X1  g0887(.A1(new_n818), .A2(new_n303), .B1(new_n287), .B2(new_n801), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT109), .Z(new_n1089));
  OAI221_X1 g0889(.A(new_n253), .B1(new_n213), .B2(new_n792), .C1(new_n789), .C2(new_n215), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n996), .A2(new_n868), .B1(new_n798), .B2(new_n202), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT110), .Z(new_n1093));
  AOI21_X1  g0893(.A(new_n253), .B1(new_n832), .B2(G107), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n469), .B2(new_n798), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n804), .A2(G322), .B1(G283), .B2(new_n793), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT111), .Z(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G294), .C2(new_n800), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n810), .A2(new_n802), .B1(new_n1068), .B2(new_n785), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT52), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n993), .C2(new_n818), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT112), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n879), .B1(new_n1093), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n777), .A2(new_n247), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n775), .B(new_n1104), .C1(G97), .C2(new_n719), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1103), .A2(new_n767), .A3(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1082), .A2(new_n1009), .B1(new_n1085), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1083), .A2(new_n1107), .ZN(G390));
  INV_X1    g0908(.A(new_n843), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n849), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n947), .B1(new_n1110), .B2(new_n916), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n702), .B(new_n845), .C1(new_n752), .C2(new_n759), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n916), .B1(new_n1112), .B2(new_n843), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n947), .B1(new_n905), .B2(new_n924), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT113), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n963), .A2(new_n1111), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n742), .A2(new_n916), .A3(G330), .A4(new_n857), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n843), .B1(new_n675), .B2(new_n848), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n916), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n946), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n948), .C1(new_n962), .C2(new_n951), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT38), .B1(new_n955), .B2(new_n959), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n946), .B1(new_n943), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n752), .A2(new_n759), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n845), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n711), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1123), .B1(new_n1130), .B2(new_n1109), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT113), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1125), .A2(new_n1134), .A3(new_n1119), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1121), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1009), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n963), .A2(new_n769), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n855), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n810), .A2(new_n469), .B1(new_n202), .B2(new_n798), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT116), .Z(new_n1142));
  NOR2_X1   g0942(.A1(new_n801), .A2(new_n830), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G283), .A2(new_n821), .B1(new_n804), .B2(G294), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n338), .A3(new_n829), .A4(new_n873), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G107), .C2(new_n864), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n864), .A2(G137), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n821), .A2(G128), .B1(new_n832), .B2(G50), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n792), .A2(new_n297), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(new_n1059), .C2(new_n798), .ZN(new_n1151));
  INV_X1    g0951(.A(G125), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n253), .B1(new_n996), .B2(new_n1152), .C1(new_n801), .C2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1151), .B(new_n1154), .C1(G132), .C2(new_n811), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1142), .A2(new_n1146), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n838), .B1(new_n324), .B2(new_n1140), .C1(new_n1156), .C2(new_n879), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT117), .Z(new_n1158));
  OAI22_X1  g0958(.A1(new_n1136), .A2(new_n1137), .B1(new_n1139), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n720), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n467), .A2(new_n743), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n691), .B(new_n1161), .C1(new_n750), .C2(new_n965), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n743), .A2(KEYINPUT115), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n857), .B1(new_n743), .B2(KEYINPUT115), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1123), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1120), .A2(new_n843), .A3(new_n1112), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n742), .A2(G330), .A3(new_n857), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1123), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1119), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT114), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1110), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n1170), .B2(new_n1110), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1162), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1160), .B1(new_n1136), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1121), .A2(new_n1135), .A3(new_n1162), .A4(new_n1175), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1159), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G378));
  AOI21_X1  g0980(.A(new_n700), .B1(new_n301), .B2(new_n308), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n322), .A2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n311), .B(new_n1181), .C1(new_n319), .C2(new_n321), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n322), .A2(new_n1182), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n1184), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n768), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n838), .B1(G50), .B2(new_n1140), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n800), .A2(new_n410), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n253), .A2(G41), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n793), .B2(G77), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(new_n213), .C2(new_n798), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n789), .A2(new_n823), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n996), .A2(new_n790), .B1(new_n469), .B2(new_n785), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n830), .B2(new_n818), .C1(new_n404), .C2(new_n810), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  INV_X1    g1002(.A(G41), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G50), .B1(new_n250), .B2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1201), .A2(new_n1202), .B1(new_n1195), .B2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n801), .A2(new_n997), .B1(new_n792), .B2(new_n1153), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n811), .B2(G128), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n864), .A2(G132), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n785), .A2(new_n1152), .B1(new_n798), .B2(new_n297), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT118), .Z(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT59), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT119), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n804), .A2(G124), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n832), .C2(G159), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1212), .A2(KEYINPUT119), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1205), .B1(new_n1202), .B2(new_n1201), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1193), .B1(new_n1218), .B2(new_n773), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1192), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n678), .B1(new_n374), .B2(KEYINPUT18), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n887), .B1(new_n1221), .B2(new_n381), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n899), .A2(new_n958), .B1(new_n953), .B2(new_n954), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1222), .A2(new_n942), .B1(new_n1223), .B2(KEYINPUT38), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n917), .A3(KEYINPUT40), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(G330), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT120), .B1(new_n1226), .B2(new_n918), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n917), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n919), .B1(new_n944), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT120), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n929), .B1(new_n925), .B2(new_n917), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1227), .A2(new_n1232), .A3(new_n1191), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(KEYINPUT120), .C1(new_n918), .C2(new_n1226), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n964), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1233), .A2(new_n964), .A3(new_n1235), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1220), .B1(new_n1240), .B2(new_n1137), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1233), .A2(new_n964), .A3(new_n1235), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n964), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1178), .A2(new_n1162), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1238), .A2(KEYINPUT57), .A3(new_n1239), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1162), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1125), .A2(new_n1134), .A3(new_n1119), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1119), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(new_n1251), .B2(new_n1175), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n720), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1246), .B1(new_n1253), .B2(KEYINPUT121), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT121), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1255), .B(new_n720), .C1(new_n1247), .C2(new_n1252), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1241), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G375));
  NAND2_X1  g1058(.A1(new_n1175), .A2(new_n1009), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1259), .A2(KEYINPUT122), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n767), .B1(new_n213), .B2(new_n855), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n338), .B(new_n1198), .C1(G159), .C2(new_n793), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n804), .A2(G128), .B1(G50), .B2(new_n797), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n297), .C2(new_n801), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT123), .Z(new_n1265));
  AOI22_X1  g1065(.A1(new_n811), .A2(G137), .B1(G132), .B2(new_n821), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n818), .C2(new_n1153), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n338), .B1(new_n830), .B2(new_n792), .C1(new_n789), .C2(new_n202), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1058), .B1(new_n585), .B2(new_n785), .C1(new_n996), .C2(new_n993), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(G107), .C2(new_n800), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1270), .B1(new_n469), .B2(new_n818), .C1(new_n790), .C2(new_n810), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1261), .B1(new_n769), .B2(new_n916), .C1(new_n1272), .C2(new_n879), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1259), .A2(KEYINPUT122), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1260), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1162), .A2(new_n1175), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1033), .A3(new_n1176), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(G381));
  INV_X1    g1079(.A(G384), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1083), .A2(new_n1280), .A3(new_n1107), .A4(new_n1281), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(G387), .A2(new_n1282), .A3(G378), .A4(G381), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1257), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT124), .Z(G407));
  NAND2_X1  g1085(.A1(new_n1179), .A2(new_n701), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G407), .B(G213), .C1(G375), .C2(new_n1286), .ZN(G409));
  XNOR2_X1  g1087(.A(G387), .B(G390), .ZN(new_n1288));
  XOR2_X1   g1088(.A(G393), .B(G396), .Z(new_n1289));
  AND2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G213), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1293), .A2(G343), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1276), .A2(KEYINPUT60), .A3(new_n1176), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n720), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1275), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1280), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1275), .A2(new_n1299), .A3(G384), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n1179), .B(new_n1241), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1244), .A2(new_n1033), .A3(new_n1245), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1179), .B1(new_n1306), .B2(new_n1241), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1309), .B(new_n1179), .C1(new_n1306), .C2(new_n1241), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1295), .B(new_n1304), .C1(new_n1305), .C2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT62), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1257), .A2(G378), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1295), .A4(new_n1304), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1295), .B1(new_n1305), .B2(new_n1311), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1294), .A2(G2897), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1301), .A2(new_n1302), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1320), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1313), .B(new_n1318), .C1(new_n1324), .C2(KEYINPUT127), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1294), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1323), .ZN(new_n1328));
  OAI211_X1 g1128(.A(KEYINPUT127), .B(new_n1326), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1292), .B1(new_n1325), .B2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1312), .A2(new_n1333), .A3(KEYINPUT63), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT63), .B1(new_n1312), .B2(new_n1333), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1332), .B(new_n1324), .C1(new_n1334), .C2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1331), .A2(new_n1336), .ZN(G405));
  NOR2_X1   g1137(.A1(new_n1257), .A2(G378), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1338), .A2(new_n1305), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(new_n1304), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1332), .ZN(G402));
endmodule


