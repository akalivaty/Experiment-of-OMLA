//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G77), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT66), .B(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n202), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT64), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n208), .A2(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n215), .B1(new_n214), .B2(new_n213), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT0), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(new_n225), .A2(new_n226), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n233), .B1(new_n226), .B2(new_n225), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n223), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G226), .B(G232), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G97), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G68), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n247), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT25), .B1(new_n256), .B2(G107), .ZN(new_n257));
  OR3_X1    g0057(.A1(new_n256), .A2(KEYINPUT25), .A3(G107), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n230), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G107), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n257), .B(new_n258), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  XOR2_X1   g0065(.A(new_n265), .B(KEYINPUT84), .Z(new_n266));
  INV_X1    g0066(.A(KEYINPUT23), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(new_n231), .B2(G107), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(KEYINPUT23), .A3(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G116), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(G20), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(new_n231), .A4(G87), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT22), .ZN(new_n279));
  INV_X1    g0079(.A(G87), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n280), .A2(KEYINPUT22), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT68), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n276), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT68), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n279), .B1(new_n288), .B2(KEYINPUT83), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT68), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT68), .B1(new_n275), .B2(new_n277), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT83), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n273), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT24), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n261), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n278), .A2(KEYINPUT22), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n292), .B2(new_n293), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n288), .A2(KEYINPUT83), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n272), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n266), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT5), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G41), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G1), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n306), .A2(G274), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G41), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(G1), .A3(G13), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n307), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n305), .ZN(new_n314));
  INV_X1    g0114(.A(G264), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n310), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT3), .B(G33), .ZN(new_n317));
  INV_X1    g0117(.A(G250), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n317), .B(new_n320), .C1(G257), .C2(new_n319), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G294), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n312), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G169), .B2(new_n324), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT85), .B1(new_n303), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n265), .B(KEYINPUT84), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n260), .B1(new_n301), .B2(KEYINPUT24), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n295), .A2(new_n296), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT85), .ZN(new_n333));
  INV_X1    g0133(.A(new_n327), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(G190), .B2(new_n324), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n328), .A2(new_n335), .B1(new_n303), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n286), .A2(new_n287), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(G222), .A3(new_n319), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(G1698), .ZN(new_n342));
  INV_X1    g0142(.A(G223), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n341), .B1(new_n207), .B2(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n312), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G274), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n312), .A2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n210), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n203), .A2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G20), .A2(G33), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT8), .B(G58), .Z(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n231), .A2(G33), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n355), .B1(new_n356), .B2(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n260), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n255), .A2(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n261), .A2(new_n364), .ZN(new_n365));
  MUX2_X1   g0165(.A(new_n256), .B(new_n365), .S(G50), .Z(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n351), .B1(new_n344), .B2(new_n345), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(G169), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n354), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n353), .A2(G200), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(G190), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n367), .B(KEYINPUT9), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT70), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT70), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n377), .A3(KEYINPUT10), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT10), .B1(new_n373), .B2(KEYINPUT69), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(new_n371), .A4(new_n372), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n370), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G238), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n349), .B1(new_n350), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(G232), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n386));
  OAI211_X1 g0186(.A(G226), .B(new_n319), .C1(new_n290), .C2(new_n291), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G97), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n385), .B1(new_n389), .B2(new_n345), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI211_X1 g0192(.A(KEYINPUT13), .B(new_n385), .C1(new_n389), .C2(new_n345), .ZN(new_n393));
  OAI21_X1  g0193(.A(G200), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n256), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n249), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT12), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n357), .A2(G50), .ZN(new_n398));
  INV_X1    g0198(.A(G77), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n398), .B1(new_n231), .B2(G68), .C1(new_n399), .C2(new_n361), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n397), .B(new_n401), .C1(new_n249), .C2(new_n365), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT11), .B1(new_n400), .B2(new_n260), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n394), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT71), .B1(new_n390), .B2(new_n391), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n391), .B2(new_n390), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n390), .A2(new_n408), .A3(new_n391), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n405), .B1(G190), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT71), .ZN(new_n413));
  OAI21_X1  g0213(.A(G179), .B1(new_n413), .B2(new_n409), .ZN(new_n414));
  OAI21_X1  g0214(.A(G169), .B1(new_n392), .B2(new_n393), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(G169), .C1(new_n392), .C2(new_n393), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n404), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n412), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n210), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n317), .B(new_n422), .C1(G223), .C2(G1698), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT75), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n312), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n349), .B1(new_n350), .B2(new_n220), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G179), .ZN(new_n429));
  INV_X1    g0229(.A(G169), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(new_n428), .ZN(new_n431));
  XNOR2_X1  g0231(.A(G58), .B(G68), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(G20), .B1(G159), .B2(new_n357), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(G20), .B1(new_n275), .B2(new_n277), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT7), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n433), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n260), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n275), .A2(new_n277), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT73), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT73), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n436), .A2(new_n447), .A3(KEYINPUT7), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n286), .A2(new_n231), .A3(new_n287), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n446), .A2(new_n448), .B1(new_n449), .B2(new_n435), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n433), .B1(new_n450), .B2(new_n249), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n443), .B1(new_n451), .B2(new_n442), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT74), .B1(new_n359), .B2(new_n364), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n453), .A2(new_n395), .A3(new_n260), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n359), .A2(KEYINPUT74), .A3(new_n364), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n454), .A2(new_n455), .B1(new_n395), .B2(new_n360), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n431), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT18), .B(new_n431), .C1(new_n452), .C2(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G190), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n426), .A2(new_n463), .A3(new_n427), .ZN(new_n464));
  INV_X1    g0264(.A(new_n428), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G200), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n290), .A2(new_n291), .A3(G20), .ZN(new_n467));
  NOR4_X1   g0267(.A1(new_n317), .A2(KEYINPUT73), .A3(new_n439), .A4(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n447), .B1(new_n436), .B2(KEYINPUT7), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n467), .A2(new_n434), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G68), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT16), .B1(new_n471), .B2(new_n433), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n456), .B(new_n466), .C1(new_n472), .C2(new_n443), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n451), .A2(new_n442), .ZN(new_n477));
  INV_X1    g0277(.A(new_n433), .ZN(new_n478));
  INV_X1    g0278(.A(new_n440), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n437), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n261), .B1(new_n480), .B2(KEYINPUT16), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n457), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n466), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n360), .A2(new_n358), .B1(new_n207), .B2(new_n231), .ZN(new_n485));
  XOR2_X1   g0285(.A(KEYINPUT15), .B(G87), .Z(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n361), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n260), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI221_X1 g0289(.A(new_n489), .B1(new_n399), .B2(new_n365), .C1(new_n208), .C2(new_n256), .ZN(new_n490));
  INV_X1    g0290(.A(new_n349), .ZN(new_n491));
  INV_X1    g0291(.A(new_n350), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n209), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n340), .A2(G232), .A3(new_n319), .ZN(new_n495));
  OAI221_X1 g0295(.A(new_n495), .B1(new_n264), .B2(new_n340), .C1(new_n342), .C2(new_n384), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(new_n345), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n497), .B2(G190), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n336), .B2(new_n497), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n497), .A2(G169), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n325), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n490), .A3(new_n501), .ZN(new_n502));
  AND4_X1   g0302(.A1(new_n462), .A2(new_n484), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n383), .A2(new_n421), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n256), .A2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(new_n263), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n264), .A2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n510), .B2(new_n246), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n512), .A2(new_n231), .B1(new_n399), .B2(new_n358), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n470), .B2(G107), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n508), .B1(new_n514), .B2(new_n261), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT77), .ZN(new_n516));
  AND2_X1   g0316(.A1(KEYINPUT4), .A2(G244), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n319), .B(new_n517), .C1(new_n290), .C2(new_n291), .ZN(new_n518));
  OAI211_X1 g0318(.A(G250), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(new_n319), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n520), .A2(new_n521), .B1(G33), .B2(G283), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n345), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(new_n312), .C1(new_n313), .C2(new_n305), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(G179), .A3(new_n310), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n525), .ZN(new_n527));
  INV_X1    g0327(.A(new_n310), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n523), .C2(new_n345), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n526), .B1(new_n529), .B2(new_n430), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n446), .A2(new_n448), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n449), .A2(new_n435), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n264), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n260), .B1(new_n533), .B2(new_n513), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n508), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n516), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(G190), .ZN(new_n538));
  INV_X1    g0338(.A(new_n508), .ZN(new_n539));
  INV_X1    g0339(.A(new_n513), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n450), .B2(new_n264), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n260), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n538), .B(new_n542), .C1(new_n336), .C2(new_n529), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n259), .A2(new_n230), .B1(G20), .B2(new_n211), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(G33), .B2(G283), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(G33), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n551), .B(KEYINPUT20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n395), .A2(new_n211), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n263), .B2(new_n211), .ZN(new_n554));
  OAI21_X1  g0354(.A(G169), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n310), .B1(new_n314), .B2(new_n212), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n317), .A2(G257), .A3(new_n319), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT81), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n286), .A2(G303), .A3(new_n287), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n317), .A2(G264), .A3(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n317), .A2(KEYINPUT81), .A3(G257), .A4(new_n319), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n563), .B2(new_n345), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n546), .B1(new_n555), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(G190), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n552), .A2(new_n554), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n568), .C1(new_n336), .C2(new_n564), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n564), .B(G179), .C1(new_n552), .C2(new_n554), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n546), .B(new_n571), .C1(new_n555), .C2(new_n564), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n275), .A2(new_n277), .A3(G238), .A4(new_n319), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n271), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n345), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT78), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n308), .B2(G1), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n255), .A2(KEYINPUT78), .A3(G45), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n312), .A2(new_n579), .A3(G250), .A4(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(KEYINPUT79), .B1(G274), .B2(new_n309), .ZN(new_n582));
  INV_X1    g0382(.A(new_n230), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n318), .B1(new_n583), .B2(new_n311), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT79), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n580), .A4(new_n579), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n577), .A2(new_n582), .A3(new_n325), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n231), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n280), .A2(new_n549), .A3(new_n264), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n275), .A2(new_n277), .A3(new_n231), .A4(G68), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n361), .B2(new_n549), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n260), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n486), .A2(new_n261), .A3(new_n256), .A4(new_n262), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n487), .A2(new_n395), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(KEYINPUT80), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n587), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n595), .A2(new_n260), .B1(new_n395), .B2(new_n487), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT80), .B1(new_n601), .B2(new_n597), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n577), .A2(new_n586), .A3(new_n582), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n430), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(G200), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n507), .A2(G87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n604), .B2(G190), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n603), .A2(new_n606), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n573), .A2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n339), .A2(new_n505), .A3(new_n545), .A4(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n379), .A2(new_n382), .ZN(new_n615));
  INV_X1    g0415(.A(new_n502), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n419), .B2(new_n420), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n476), .A2(new_n483), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n617), .A2(new_n412), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n460), .A2(new_n461), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n370), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n338), .B(new_n329), .C1(new_n331), .C2(new_n330), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n581), .A2(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n309), .A2(G274), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n586), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n345), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT86), .B1(new_n576), .B2(new_n345), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n430), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(G200), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n603), .A2(new_n633), .B1(new_n634), .B2(new_n610), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n537), .A2(new_n625), .A3(new_n543), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n601), .A2(new_n597), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT80), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n587), .A3(new_n599), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT86), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n577), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n345), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(G169), .B1(new_n645), .B2(new_n629), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n336), .B1(new_n645), .B2(new_n629), .ZN(new_n647));
  INV_X1    g0447(.A(new_n609), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n577), .A2(new_n582), .A3(G190), .A4(new_n586), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n641), .A2(new_n646), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n303), .B2(new_n338), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT87), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n537), .A4(new_n543), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n303), .A2(new_n327), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n566), .A2(new_n570), .A3(new_n572), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n637), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n603), .A2(new_n633), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n634), .A2(new_n610), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n530), .A2(new_n659), .A3(new_n660), .A4(new_n515), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n603), .B2(new_n633), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n641), .A2(new_n646), .A3(KEYINPUT88), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n661), .A2(KEYINPUT26), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g0465(.A(KEYINPUT77), .B(new_n539), .C1(new_n541), .C2(new_n260), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n535), .B1(new_n534), .B2(new_n508), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n530), .A3(new_n611), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(KEYINPUT26), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n658), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n624), .B1(new_n504), .B2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n255), .A2(new_n231), .A3(G13), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n678));
  INV_X1    g0478(.A(G213), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n339), .A2(new_n656), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n655), .B2(new_n684), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n568), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n656), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n573), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n332), .A2(new_n683), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n339), .A2(new_n692), .B1(new_n655), .B2(new_n683), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n687), .B1(new_n691), .B2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n224), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n590), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n228), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT29), .B1(new_n671), .B2(new_n684), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n656), .B1(new_n328), .B2(new_n335), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n636), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT90), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n664), .B2(new_n663), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT88), .B1(new_n641), .B2(new_n646), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n603), .A2(new_n633), .A3(new_n662), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n661), .A2(KEYINPUT26), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT26), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n668), .A2(new_n712), .A3(new_n530), .A4(new_n611), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n684), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n684), .C1(new_n704), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n702), .B1(new_n719), .B2(KEYINPUT29), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n564), .A2(G179), .A3(new_n324), .A4(new_n604), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n527), .B1(new_n523), .B2(new_n345), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR3_X1    g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n722), .B2(new_n725), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n564), .A2(G179), .A3(new_n324), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n310), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n632), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n731), .B2(new_n683), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n339), .A2(new_n545), .A3(new_n613), .A4(new_n684), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n721), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n720), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n701), .B1(new_n737), .B2(G1), .ZN(G364));
  AND2_X1   g0538(.A1(new_n231), .A2(G13), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n255), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n696), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n691), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n690), .A2(G330), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n690), .A2(G20), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n230), .B1(G20), .B2(new_n430), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n231), .A2(new_n325), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(G190), .A3(new_n336), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n231), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n336), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n752), .A2(G58), .B1(new_n756), .B2(G107), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n325), .A2(new_n336), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n231), .A2(new_n463), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n754), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n757), .B1(new_n202), .B2(new_n760), .C1(new_n280), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n753), .A2(new_n325), .A3(new_n336), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G159), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n463), .A2(G179), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n231), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n549), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n758), .A2(new_n753), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n750), .A2(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n340), .B1(new_n249), .B2(new_n770), .C1(new_n207), .C2(new_n772), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n762), .A2(new_n766), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n764), .A2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT33), .B(G317), .Z(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n776), .B2(new_n772), .C1(new_n770), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n340), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n768), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n751), .A2(new_n782), .B1(new_n755), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n760), .A2(new_n785), .B1(new_n761), .B2(new_n786), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n778), .A2(new_n781), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n749), .B1(new_n774), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n779), .A2(new_n695), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G355), .B1(new_n211), .B2(new_n695), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n253), .A2(new_n308), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n695), .A2(new_n317), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n228), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n747), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n749), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n743), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n789), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT92), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n744), .A2(new_n745), .B1(new_n748), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT93), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n490), .A2(new_n683), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n499), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n502), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n616), .A2(new_n684), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n672), .B2(new_n683), .ZN(new_n809));
  INV_X1    g0609(.A(new_n808), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n671), .A2(new_n684), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n736), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n742), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n749), .A2(new_n746), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n743), .B1(new_n399), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n749), .ZN(new_n818));
  INV_X1    g0618(.A(new_n770), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n752), .A2(G143), .B1(new_n819), .B2(G150), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G159), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n760), .C1(new_n822), .C2(new_n772), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n317), .B1(new_n761), .B2(new_n202), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n763), .A2(new_n828), .B1(new_n755), .B2(new_n249), .ZN(new_n829));
  INV_X1    g0629(.A(new_n768), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n827), .B(new_n829), .C1(G58), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n825), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n776), .A2(new_n763), .B1(new_n770), .B2(new_n783), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n760), .A2(new_n786), .B1(new_n761), .B2(new_n264), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n833), .A2(new_n834), .A3(new_n769), .A4(new_n340), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n755), .A2(new_n280), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G294), .B2(new_n752), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n835), .B(new_n837), .C1(new_n211), .C2(new_n772), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n817), .B1(new_n818), .B2(new_n839), .C1(new_n810), .C2(new_n747), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n815), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(new_n512), .ZN(new_n842));
  OAI211_X1 g0642(.A(G116), .B(new_n232), .C1(new_n842), .C2(KEYINPUT35), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(KEYINPUT35), .B2(new_n842), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n229), .B(new_n208), .C1(new_n219), .C2(new_n249), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n255), .B(G13), .C1(new_n846), .C2(new_n248), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n481), .B1(KEYINPUT16), .B2(new_n480), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n456), .ZN(new_n852));
  INV_X1    g0652(.A(new_n681), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n431), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n850), .B1(new_n854), .B2(new_n473), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n458), .A2(new_n473), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT95), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n857), .B(new_n853), .C1(new_n452), .C2(new_n457), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT95), .B1(new_n482), .B2(new_n681), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n855), .B1(new_n860), .B2(new_n850), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n852), .A2(new_n853), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n484), .B2(new_n462), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n849), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT96), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n858), .ZN(new_n866));
  INV_X1    g0666(.A(new_n856), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(new_n850), .ZN(new_n868));
  INV_X1    g0668(.A(new_n855), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n862), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n620), .B2(new_n618), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n864), .A2(new_n865), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT96), .A4(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n734), .A2(new_n735), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n416), .A2(new_n418), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n325), .B1(new_n407), .B2(new_n410), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n420), .B(new_n683), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT94), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT94), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n419), .A2(new_n883), .A3(new_n420), .A4(new_n683), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n420), .A2(new_n683), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n882), .A2(new_n884), .B1(new_n421), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n878), .A2(new_n886), .A3(new_n808), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n877), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n866), .A2(new_n867), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n868), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n866), .B1(new_n484), .B2(new_n462), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n849), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n895), .B2(new_n873), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n888), .A2(new_n889), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n813), .A2(new_n504), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n897), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n504), .A2(new_n878), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n729), .A2(G169), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n542), .B1(new_n905), .B2(new_n526), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n712), .B1(new_n906), .B2(new_n635), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n537), .A2(new_n612), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n712), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(new_n710), .C1(new_n636), .C2(new_n703), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n717), .B1(new_n910), .B2(new_n684), .ZN(new_n911));
  INV_X1    g0711(.A(new_n718), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT29), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n702), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n505), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT97), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n720), .A2(KEYINPUT97), .A3(new_n505), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n623), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n904), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n886), .B1(new_n811), .B2(new_n807), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n877), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n895), .A2(new_n924), .A3(new_n873), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n419), .A2(new_n420), .A3(new_n684), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n922), .B1(new_n462), .B2(new_n853), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT98), .Z(new_n930));
  NAND2_X1  g0730(.A1(new_n920), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n255), .B2(new_n739), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n920), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n848), .B1(new_n932), .B2(new_n933), .ZN(G367));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n542), .A2(new_n684), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n530), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT100), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n544), .A2(new_n936), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n687), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT45), .Z(new_n943));
  OR3_X1    g0743(.A1(new_n687), .A2(KEYINPUT102), .A3(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT102), .B1(new_n687), .B2(new_n941), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  OAI211_X1 g0748(.A(KEYINPUT102), .B(new_n948), .C1(new_n687), .C2(new_n941), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n943), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n693), .A2(new_n691), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n656), .A2(new_n684), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n686), .B1(new_n693), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n691), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n737), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n950), .A2(new_n951), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT103), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n736), .B(new_n720), .C1(new_n953), .C2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n696), .B(KEYINPUT41), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n935), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n953), .A2(new_n960), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n737), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(KEYINPUT104), .A3(new_n962), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n740), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n941), .A2(new_n686), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n328), .A2(new_n335), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n537), .B1(new_n940), .B2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n969), .A2(KEYINPUT42), .B1(new_n971), .B2(new_n684), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(KEYINPUT42), .B2(new_n969), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n635), .B1(new_n648), .B2(new_n684), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n707), .A2(new_n708), .A3(new_n609), .A4(new_n683), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n973), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n974), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n951), .A2(new_n941), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n978), .A2(new_n796), .ZN(new_n984));
  INV_X1    g0784(.A(new_n793), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n243), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n797), .B1(new_n224), .B2(new_n487), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n742), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n761), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(G116), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n444), .B1(new_n780), .B2(new_n770), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n755), .A2(new_n549), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n751), .A2(new_n786), .B1(new_n763), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n760), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n996), .C1(G311), .C2(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n768), .A2(new_n264), .B1(new_n772), .B2(new_n783), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT105), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n993), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n768), .A2(new_n249), .B1(new_n751), .B2(new_n356), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT106), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(G143), .B2(new_n997), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT107), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n989), .A2(G58), .B1(new_n756), .B2(new_n208), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n821), .B2(new_n763), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n779), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n202), .A2(new_n772), .B1(new_n770), .B2(new_n822), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT108), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1006), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1005), .A2(KEYINPUT107), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1001), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT47), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n818), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n988), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n968), .A2(new_n983), .B1(new_n984), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT109), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n240), .A2(G45), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n359), .A2(new_n202), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1025));
  XOR2_X1   g0825(.A(new_n1024), .B(new_n1025), .Z(new_n1026));
  OAI211_X1 g0826(.A(new_n698), .B(new_n308), .C1(new_n249), .C2(new_n399), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1023), .B(new_n793), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n340), .A2(new_n224), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(G107), .B2(new_n224), .C1(new_n698), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1030), .A2(KEYINPUT111), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n797), .B1(new_n1030), .B2(KEYINPUT111), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n994), .A2(new_n444), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n989), .A2(new_n208), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n356), .C2(new_n763), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n360), .A2(new_n770), .B1(new_n202), .B2(new_n751), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n760), .A2(new_n822), .B1(new_n772), .B2(new_n249), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n487), .A2(new_n768), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n444), .B1(new_n763), .B2(new_n785), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n830), .A2(G283), .B1(new_n989), .B2(G294), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n772), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G322), .A2(new_n997), .B1(new_n1042), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n776), .B2(new_n770), .C1(new_n995), .C2(new_n751), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT112), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT49), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1040), .B(new_n1049), .C1(G116), .C2(new_n756), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n742), .B1(new_n1031), .B2(new_n1032), .C1(new_n1052), .C2(new_n818), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT113), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n693), .B2(new_n796), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n956), .B2(new_n741), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n697), .B1(new_n737), .B2(new_n956), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n737), .B2(new_n956), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(G393));
  AOI21_X1  g0859(.A(new_n697), .B1(new_n952), .B2(new_n957), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n965), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n952), .A2(new_n740), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n940), .A2(new_n796), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n247), .A2(new_n985), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n797), .B1(new_n549), .B2(new_n224), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n742), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n752), .A2(G159), .B1(new_n997), .B2(G150), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G143), .A2(new_n764), .B1(new_n989), .B2(G68), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1067), .A2(KEYINPUT51), .B1(new_n1068), .B2(KEYINPUT114), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n360), .A2(new_n772), .B1(new_n202), .B2(new_n770), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n768), .A2(new_n399), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1071), .A2(new_n1072), .A3(new_n444), .A4(new_n836), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1068), .A2(KEYINPUT114), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n782), .A2(new_n763), .B1(new_n761), .B2(new_n783), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT115), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n770), .A2(new_n786), .B1(new_n755), .B2(new_n264), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G294), .B2(new_n1042), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n340), .B1(G116), .B2(new_n830), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n751), .A2(new_n776), .B1(new_n760), .B2(new_n995), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI21_X1  g0883(.A(new_n1075), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1066), .B1(new_n1084), .B2(new_n749), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1062), .B1(new_n1063), .B2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1061), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  AOI21_X1  g0888(.A(KEYINPUT97), .B1(new_n720), .B2(new_n505), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT29), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n716), .B2(new_n718), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1091), .A2(new_n916), .A3(new_n702), .A4(new_n504), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n624), .B(new_n900), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n811), .A2(new_n807), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n882), .A2(new_n884), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n421), .A2(new_n885), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n736), .A3(new_n810), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT116), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n808), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n736), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n736), .A2(new_n810), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n886), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1104), .A2(new_n1098), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n716), .A2(new_n718), .A3(new_n807), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n806), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1094), .A2(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1093), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n928), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n923), .B(new_n925), .C1(new_n921), .C2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1107), .A2(new_n806), .A3(new_n1097), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1112), .B1(new_n895), .B2(new_n873), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n736), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT116), .B1(new_n1101), .B2(new_n736), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1113), .A2(new_n1116), .A3(new_n1098), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1111), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1105), .A2(new_n1094), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n919), .A2(new_n1128), .A3(new_n900), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT117), .B1(new_n1129), .B2(new_n1124), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1113), .A2(new_n1116), .A3(new_n1098), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1120), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1093), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1128), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n697), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n927), .A2(new_n746), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n816), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n742), .B1(new_n359), .B2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n549), .A2(new_n772), .B1(new_n770), .B2(new_n264), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n761), .A2(new_n280), .B1(new_n755), .B2(new_n249), .ZN(new_n1143));
  OR4_X1    g0943(.A1(new_n340), .A2(new_n1142), .A3(new_n1143), .A4(new_n1072), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G283), .A2(new_n997), .B1(new_n764), .B2(G294), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n211), .B2(new_n751), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n761), .A2(new_n356), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G128), .A2(new_n997), .B1(new_n756), .B2(G50), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT54), .B(G143), .Z(new_n1150));
  AOI22_X1  g0950(.A1(G125), .A2(new_n764), .B1(new_n1042), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n752), .A2(G132), .B1(new_n819), .B2(G137), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n340), .C1(new_n822), .C2(new_n768), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1144), .A2(new_n1146), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1141), .B1(new_n1155), .B2(new_n749), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1133), .A2(new_n741), .B1(new_n1139), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1138), .A2(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n615), .A2(new_n622), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT55), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n367), .A2(new_n853), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n383), .A2(KEYINPUT55), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1165), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1161), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(new_n1160), .A3(new_n1167), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1172), .A3(KEYINPUT121), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n897), .A3(G330), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1173), .B1(new_n897), .B2(G330), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n929), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n898), .A2(KEYINPUT121), .A3(new_n1172), .A4(new_n1170), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n929), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n1174), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1093), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(KEYINPUT122), .B(new_n1093), .C1(new_n1130), .C2(new_n1136), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1159), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1129), .A2(new_n1124), .A3(KEYINPUT117), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1135), .B1(new_n1110), .B2(new_n1133), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1134), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT122), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(KEYINPUT57), .A3(new_n1191), .A4(new_n1181), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1186), .A2(new_n1192), .A3(new_n696), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1170), .A2(new_n1172), .A3(new_n746), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n742), .B1(G50), .B2(new_n1140), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n317), .A2(G41), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n751), .A2(new_n264), .B1(new_n755), .B2(new_n219), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1034), .A2(new_n1196), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G68), .C2(new_n830), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G116), .A2(new_n997), .B1(new_n764), .B2(G283), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G97), .A2(new_n819), .B1(new_n1042), .B2(new_n486), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT58), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1198), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n997), .A2(G125), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n828), .B2(new_n770), .C1(new_n821), .C2(new_n772), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n752), .A2(G128), .B1(new_n989), .B2(new_n1150), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT119), .Z(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G150), .C2(new_n830), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1207), .B1(new_n822), .B2(new_n755), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1206), .B1(new_n1205), .B2(new_n1204), .C1(new_n1214), .C2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1195), .B1(new_n1217), .B2(new_n749), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1181), .A2(new_n741), .B1(new_n1194), .B2(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1193), .A2(KEYINPUT123), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT123), .B1(new_n1193), .B2(new_n1219), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1093), .A2(new_n1109), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1111), .A2(new_n962), .A3(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1097), .A2(new_n747), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT124), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(KEYINPUT124), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n760), .A2(new_n780), .B1(new_n770), .B2(new_n211), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n772), .A2(new_n264), .B1(new_n755), .B2(new_n399), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1038), .A4(new_n340), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G303), .A2(new_n764), .B1(new_n989), .B2(G97), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n783), .C2(new_n751), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n751), .A2(new_n821), .B1(new_n760), .B2(new_n828), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n444), .B(new_n1235), .C1(G58), .C2(new_n756), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G128), .A2(new_n764), .B1(new_n989), .B2(G159), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G150), .A2(new_n1042), .B1(new_n819), .B2(new_n1150), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n830), .A2(G50), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n818), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n743), .B(new_n1241), .C1(new_n249), .C2(new_n816), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT125), .Z(new_n1243));
  NOR3_X1   g1043(.A1(new_n1228), .A2(new_n1229), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1128), .B2(new_n741), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1225), .A2(new_n1245), .ZN(G381));
  NOR3_X1   g1046(.A1(new_n1220), .A2(new_n1221), .A3(G378), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1056), .A2(new_n802), .A3(new_n1058), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1021), .A2(new_n1247), .A3(new_n1249), .ZN(G407));
  NAND2_X1  g1050(.A1(new_n1193), .A2(new_n1219), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G378), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1193), .A2(KEYINPUT123), .A3(new_n1219), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1061), .A2(new_n1086), .B1(new_n1258), .B2(new_n1248), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1248), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1020), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1087), .B2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1019), .B(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1224), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n696), .A3(new_n1129), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1245), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(G384), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n682), .A2(G213), .A3(G2897), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1271), .B(new_n1272), .Z(new_n1273));
  AOI21_X1  g1073(.A(new_n1254), .B1(new_n1193), .B2(new_n1219), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1175), .A2(new_n1176), .A3(new_n929), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1179), .B1(new_n1178), .B2(new_n1174), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT126), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1177), .A2(new_n1180), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n741), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1194), .A2(new_n1218), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1138), .A3(new_n1157), .A4(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1184), .A2(new_n963), .A3(new_n1185), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1282), .A2(new_n1283), .B1(new_n679), .B2(G343), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1273), .B1(new_n1274), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1271), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1274), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1265), .B(new_n1285), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1251), .A2(G378), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1284), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1271), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1264), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1285), .A2(new_n1265), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n1297), .A3(new_n1263), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(G405));
  XOR2_X1   g1100(.A(new_n1271), .B(KEYINPUT127), .Z(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1256), .A2(new_n1290), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1256), .B2(new_n1290), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1264), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1301), .B1(new_n1247), .B2(new_n1274), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1256), .A2(new_n1290), .A3(new_n1302), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1263), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(G402));
endmodule


