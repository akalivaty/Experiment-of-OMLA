//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(G101), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n464), .A2(new_n466), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(G2105), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n462), .A3(new_n485), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n481), .B1(new_n486), .B2(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT69), .Z(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NOR2_X1   g067(.A1(new_n463), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G102), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(new_n463), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n475), .B2(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(new_n462), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n462), .A2(G138), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n475), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n462), .A2(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n468), .B2(new_n469), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n500), .A2(new_n499), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT67), .B1(new_n473), .B2(new_n474), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n498), .B1(new_n506), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n514), .A2(new_n516), .A3(new_n522), .A4(new_n524), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n521), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR3_X1    g112(.A1(new_n535), .A2(new_n534), .A3(new_n536), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n533), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n526), .A2(new_n540), .B1(new_n541), .B2(new_n529), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI221_X1 g124(.A(new_n547), .B1(new_n548), .B2(new_n526), .C1(new_n549), .C2(new_n529), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AOI22_X1  g126(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n520), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n526), .A2(new_n554), .B1(new_n555), .B2(new_n529), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n517), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n525), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G53), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n571), .B2(G53), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n569), .B1(new_n570), .B2(new_n529), .C1(new_n573), .C2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND2_X1  g152(.A1(new_n571), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(new_n529), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G87), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n514), .A2(new_n516), .A3(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n520), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n518), .A2(new_n525), .A3(G86), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n522), .A2(new_n524), .A3(G48), .A4(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G305));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n526), .A2(new_n590), .B1(new_n591), .B2(new_n529), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n520), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n580), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n517), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n571), .A2(G54), .B1(new_n603), .B2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT74), .ZN(G284));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(new_n486), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G123), .ZN(new_n620));
  INV_X1    g195(.A(new_n489), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n462), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n620), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n508), .A2(new_n509), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n493), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT75), .Z(G156));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT77), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT78), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2084), .B(G2090), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT80), .Z(new_n662));
  NOR3_X1   g237(.A1(new_n654), .A2(new_n658), .A3(new_n656), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n654), .A2(new_n658), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n665), .B(new_n656), .C1(new_n660), .C2(new_n654), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT81), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n678), .A2(KEYINPUT20), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n681), .B(new_n683), .C1(KEYINPUT20), .C2(new_n678), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1991), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G19), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n558), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G1341), .Z(new_n694));
  NOR2_X1   g269(.A1(G4), .A2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT84), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n605), .B2(new_n691), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1348), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G168), .A2(G16), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G16), .B2(G21), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  INV_X1    g280(.A(G28), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n625), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G5), .A2(G16), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G171), .B2(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G1961), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n705), .A2(new_n711), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n704), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2078), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n712), .A2(G27), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  INV_X1    g298(.A(G126), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n484), .A2(new_n724), .B1(new_n495), .B2(new_n463), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n725), .A2(G2105), .B1(G102), .B2(new_n493), .ZN(new_n726));
  OAI21_X1  g301(.A(KEYINPUT4), .B1(new_n484), .B2(new_n502), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n510), .B2(KEYINPUT70), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n504), .A2(new_n505), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(G29), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n699), .B(new_n720), .C1(new_n721), .C2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G299), .B2(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n691), .A2(G20), .ZN(new_n735));
  MUX2_X1   g310(.A(new_n733), .B(new_n734), .S(new_n735), .Z(new_n736));
  INV_X1    g311(.A(G1956), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n619), .A2(G129), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n621), .A2(G141), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT26), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n746), .A2(new_n747), .B1(G105), .B2(new_n493), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n742), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n739), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n731), .A2(new_n721), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n738), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n712), .A2(G33), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n493), .A2(G103), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n489), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT86), .Z(new_n762));
  AOI22_X1  g337(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(new_n462), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT87), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n757), .B1(new_n767), .B2(new_n712), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2072), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n732), .A2(new_n756), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n771));
  INV_X1    g346(.A(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G29), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n491), .B2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n773), .B1(new_n775), .B2(new_n771), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n752), .A2(new_n753), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n712), .B1(KEYINPUT24), .B2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(KEYINPUT24), .B2(G34), .ZN(new_n781));
  INV_X1    g356(.A(G160), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT88), .Z(new_n784));
  OAI221_X1 g359(.A(new_n779), .B1(G1961), .B2(new_n715), .C1(G2084), .C2(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT92), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(KEYINPUT92), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n718), .A2(new_n719), .B1(G2084), .B2(new_n784), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n712), .A2(G26), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT85), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  INV_X1    g368(.A(G140), .ZN(new_n794));
  OAI221_X1 g369(.A(new_n792), .B1(new_n486), .B2(new_n793), .C1(new_n794), .C2(new_n489), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(G29), .ZN(new_n796));
  MUX2_X1   g371(.A(new_n789), .B(new_n796), .S(KEYINPUT28), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n770), .A2(new_n778), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n691), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n691), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1971), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G23), .ZN(new_n807));
  INV_X1    g382(.A(G288), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G6), .B(G305), .S(G16), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n806), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G24), .B(G290), .S(G16), .Z(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1986), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n619), .A2(G119), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n621), .A2(G131), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n462), .A2(G107), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(G29), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n818), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT83), .Z(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n817), .B2(new_n816), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n802), .A2(new_n803), .B1(new_n833), .B2(new_n834), .ZN(G311));
  XNOR2_X1  g410(.A(new_n832), .B(KEYINPUT36), .ZN(new_n836));
  INV_X1    g411(.A(new_n803), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n800), .A2(new_n801), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(G150));
  NOR2_X1   g414(.A1(new_n605), .A2(new_n613), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n571), .A2(G55), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT96), .B(G93), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OAI221_X1 g420(.A(new_n843), .B1(new_n529), .B2(new_n844), .C1(new_n520), .C2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n557), .B(new_n846), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n846), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  NAND2_X1  g428(.A1(new_n619), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n621), .A2(G142), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n462), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n795), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n750), .B(new_n825), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n767), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n767), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  INV_X1    g440(.A(new_n859), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT97), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G164), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n625), .B(G160), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n491), .Z(new_n874));
  NAND3_X1  g449(.A1(new_n864), .A2(new_n867), .A3(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n874), .B1(new_n872), .B2(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI211_X1 g456(.A(KEYINPUT98), .B(new_n874), .C1(new_n872), .C2(new_n875), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT40), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n878), .B(new_n885), .C1(new_n881), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(G303), .B(G288), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n890), .B(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n847), .B(new_n615), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n605), .B(G299), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(KEYINPUT41), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n896), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n894), .B2(new_n895), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(KEYINPUT100), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(KEYINPUT100), .ZN(new_n904));
  OAI21_X1  g479(.A(G868), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n846), .A2(new_n609), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n906), .ZN(G331));
  XNOR2_X1  g483(.A(G301), .B(G168), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n847), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n910), .A2(new_n897), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n893), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n890), .B(new_n891), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n916), .A3(new_n877), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n913), .A2(new_n916), .A3(new_n919), .A4(new_n877), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(KEYINPUT44), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n922), .A3(new_n920), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n925), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G164), .B2(G1384), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G40), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n472), .A2(new_n930), .A3(new_n478), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n750), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n795), .B(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n825), .B(new_n828), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n932), .ZN(new_n940));
  NOR2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT102), .ZN(new_n943));
  NAND2_X1  g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT106), .B(G8), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n504), .A2(new_n505), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n511), .A2(new_n949), .A3(new_n727), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n950), .B2(new_n726), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n951), .B2(new_n931), .ZN(new_n952));
  INV_X1    g527(.A(G1981), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n586), .A2(new_n953), .A3(new_n587), .A4(new_n588), .ZN(new_n954));
  INV_X1    g529(.A(G86), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n588), .B1(new_n529), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G1981), .B1(new_n956), .B2(new_n585), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n961), .B(KEYINPUT49), .C1(new_n954), .C2(new_n957), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n954), .A2(new_n957), .A3(KEYINPUT49), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI211_X1 g539(.A(G1976), .B(G288), .C1(new_n964), .C2(new_n952), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n954), .B(KEYINPUT108), .Z(new_n966));
  OAI21_X1  g541(.A(new_n952), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n730), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n928), .A2(new_n970), .A3(G40), .A4(G160), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT103), .B(G1971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n730), .A2(new_n975), .A3(new_n969), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT104), .B(G2090), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n976), .A3(new_n931), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n968), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT55), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n973), .A2(KEYINPUT105), .A3(new_n978), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n931), .A2(new_n730), .A3(new_n969), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n808), .A2(G1976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n947), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n958), .A2(new_n959), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n963), .B1(new_n991), .B2(new_n961), .ZN(new_n992));
  INV_X1    g567(.A(new_n962), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n952), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(G288), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n952), .A2(new_n988), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n990), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n967), .B1(new_n986), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n979), .A2(new_n947), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n983), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n964), .A2(new_n952), .B1(new_n989), .B2(KEYINPUT52), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(KEYINPUT109), .A3(new_n997), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n986), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n971), .B2(new_n702), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n974), .A2(new_n976), .A3(new_n931), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2084), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n971), .A2(KEYINPUT110), .A3(new_n702), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n948), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G168), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1000), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT63), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT109), .B1(new_n1005), .B2(new_n997), .ZN(new_n1018));
  AND4_X1   g593(.A1(KEYINPUT109), .A2(new_n990), .A3(new_n994), .A4(new_n997), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n948), .B1(new_n973), .B2(new_n978), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n1018), .A2(new_n1019), .B1(new_n984), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n971), .A2(new_n702), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1011), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1013), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n947), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(G286), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1022), .A2(new_n1029), .A3(KEYINPUT111), .A4(new_n986), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1016), .A2(new_n1017), .A3(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1015), .A2(new_n1017), .A3(new_n998), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n981), .A2(new_n985), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n983), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n986), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n999), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n1037));
  INV_X1    g612(.A(G1348), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1010), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n987), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n951), .A2(KEYINPUT114), .A3(new_n931), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n935), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1043), .A3(KEYINPUT60), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n606), .A2(KEYINPUT119), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n605), .B(KEYINPUT119), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(new_n1039), .A3(new_n1043), .A4(KEYINPUT60), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1046), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n971), .A2(G1996), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT58), .B(G1341), .Z(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n558), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(KEYINPUT59), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1060), .B1(new_n1058), .B2(KEYINPUT59), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n558), .B(new_n1062), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1052), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n730), .A2(new_n969), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n930), .B1(new_n1066), .B2(new_n927), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(G160), .A3(new_n970), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1070), .A2(KEYINPUT112), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n573), .A2(new_n575), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n569), .B1(new_n570), .B2(new_n529), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(KEYINPUT112), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1075), .B(KEYINPUT113), .Z(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(G299), .A2(new_n1071), .A3(new_n1076), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1010), .A2(new_n737), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1069), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1069), .B2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1065), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1084), .A2(new_n1085), .B1(new_n1086), .B2(KEYINPUT118), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1069), .A2(new_n1081), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1080), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1069), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT61), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1064), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n606), .A3(new_n1047), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1090), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1037), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1052), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1092), .A2(KEYINPUT61), .B1(new_n1102), .B2(new_n1093), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1084), .A2(new_n1094), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1099), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(KEYINPUT120), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n971), .B2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1010), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n721), .A2(KEYINPUT53), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n470), .A2(new_n471), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(KEYINPUT124), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n462), .B1(new_n1115), .B2(KEYINPUT124), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n478), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1067), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1110), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1120), .A2(G171), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1067), .A2(new_n1114), .A3(G160), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1110), .A2(new_n1122), .A3(new_n1112), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(G171), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n985), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT105), .B1(new_n973), .B2(new_n978), .ZN(new_n1127));
  NOR4_X1   g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n968), .A4(new_n983), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT125), .B1(new_n1128), .B2(new_n1021), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n986), .A2(new_n1130), .A3(new_n1002), .A4(new_n1007), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1110), .A2(G301), .A3(new_n1122), .A4(new_n1112), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT54), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1120), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1110), .A2(KEYINPUT126), .A3(new_n1119), .A4(new_n1112), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1133), .B(new_n1136), .C1(new_n1140), .C2(G301), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT127), .B1(new_n1142), .B2(new_n1135), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n971), .A2(KEYINPUT110), .A3(new_n702), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1147), .B2(new_n968), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1027), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G168), .A2(new_n948), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1150), .A2(KEYINPUT51), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1014), .B2(KEYINPUT122), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1028), .A2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1152), .A2(KEYINPUT51), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1027), .A2(new_n1150), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1132), .B(new_n1144), .C1(new_n1158), .C2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1036), .B1(new_n1108), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT62), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1027), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1150), .B1(new_n1167), .B2(new_n1145), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1168), .B2(new_n1149), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1164), .B(new_n1159), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1124), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1163), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n946), .B1(new_n1162), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n940), .A2(KEYINPUT46), .A3(new_n933), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT46), .B1(new_n940), .B2(new_n933), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n932), .B1(new_n751), .B2(new_n936), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT47), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n942), .A2(new_n932), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1179), .A2(KEYINPUT48), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(KEYINPUT48), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n939), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n937), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n825), .A2(new_n827), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1183), .A2(new_n1184), .B1(G2067), .B2(new_n795), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1178), .B(new_n1182), .C1(new_n940), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1173), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g762(.A1(new_n651), .A2(G319), .ZN(new_n1189));
  OR2_X1    g763(.A1(G227), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g764(.A1(G229), .A2(new_n1190), .ZN(new_n1191));
  AND4_X1   g765(.A1(new_n883), .A2(new_n924), .A3(new_n923), .A4(new_n1191), .ZN(G308));
  NAND4_X1  g766(.A1(new_n883), .A2(new_n924), .A3(new_n923), .A4(new_n1191), .ZN(G225));
endmodule


