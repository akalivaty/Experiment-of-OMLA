

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790;

  AND2_X1 U373 ( .A1(n408), .A2(n407), .ZN(n389) );
  XNOR2_X1 U374 ( .A(n598), .B(KEYINPUT101), .ZN(n478) );
  AND2_X1 U375 ( .A1(n392), .A2(n430), .ZN(n598) );
  XNOR2_X1 U376 ( .A(n557), .B(n385), .ZN(n392) );
  XNOR2_X2 U377 ( .A(n349), .B(n386), .ZN(n477) );
  NAND2_X2 U378 ( .A1(n458), .A2(n457), .ZN(n349) );
  NAND2_X2 U379 ( .A1(n350), .A2(n360), .ZN(n429) );
  AND2_X2 U380 ( .A1(n362), .A2(n357), .ZN(n350) );
  NOR2_X1 U381 ( .A1(n697), .A2(n699), .ZN(n438) );
  XOR2_X1 U382 ( .A(n630), .B(n479), .Z(n351) );
  XNOR2_X1 U383 ( .A(n433), .B(n447), .ZN(n679) );
  AND2_X1 U384 ( .A1(n404), .A2(KEYINPUT48), .ZN(n352) );
  AND2_X2 U385 ( .A1(n679), .A2(KEYINPUT34), .ZN(n370) );
  XNOR2_X2 U386 ( .A(n448), .B(n372), .ZN(n747) );
  BUF_X2 U387 ( .A(n586), .Z(n657) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n580) );
  AND2_X1 U389 ( .A1(n717), .A2(n716), .ZN(n720) );
  AND2_X1 U390 ( .A1(n358), .A2(n646), .ZN(n357) );
  AND2_X1 U391 ( .A1(n401), .A2(n426), .ZN(n724) );
  NAND2_X1 U392 ( .A1(n400), .A2(n686), .ZN(n366) );
  NAND2_X1 U393 ( .A1(n369), .A2(n622), .ZN(n368) );
  NAND2_X1 U394 ( .A1(n376), .A2(n397), .ZN(n687) );
  AND2_X1 U395 ( .A1(n617), .A2(n354), .ZN(n353) );
  NAND2_X1 U396 ( .A1(n393), .A2(n594), .ZN(n433) );
  INV_X1 U397 ( .A(n617), .ZN(n355) );
  INV_X1 U398 ( .A(n656), .ZN(n430) );
  OR2_X1 U399 ( .A1(n510), .A2(n513), .ZN(n509) );
  XNOR2_X1 U400 ( .A(n489), .B(n551), .ZN(n660) );
  OR2_X1 U401 ( .A1(n713), .A2(G902), .ZN(n464) );
  OR2_X1 U402 ( .A1(n693), .A2(n517), .ZN(n490) );
  NOR2_X1 U403 ( .A1(G902), .A2(n747), .ZN(n557) );
  XNOR2_X1 U404 ( .A(n356), .B(n474), .ZN(n693) );
  XNOR2_X1 U405 ( .A(n767), .B(n475), .ZN(n356) );
  XNOR2_X1 U406 ( .A(n560), .B(n518), .ZN(n767) );
  XNOR2_X1 U407 ( .A(n476), .B(n531), .ZN(n475) );
  XNOR2_X1 U408 ( .A(n519), .B(n530), .ZN(n560) );
  XNOR2_X1 U409 ( .A(n364), .B(G116), .ZN(n519) );
  INV_X1 U410 ( .A(n556), .ZN(n449) );
  XOR2_X1 U411 ( .A(G146), .B(G140), .Z(n553) );
  NAND2_X1 U412 ( .A1(n355), .A2(KEYINPUT77), .ZN(n455) );
  INV_X1 U413 ( .A(n671), .ZN(n354) );
  NAND2_X1 U414 ( .A1(n440), .A2(n355), .ZN(n456) );
  NAND2_X1 U415 ( .A1(n389), .A2(n404), .ZN(n363) );
  NAND2_X1 U416 ( .A1(n352), .A2(n389), .ZN(n362) );
  OR2_X1 U417 ( .A1(n410), .A2(n488), .ZN(n358) );
  NAND2_X1 U418 ( .A1(n363), .A2(n361), .ZN(n360) );
  AND2_X1 U419 ( .A1(n410), .A2(n488), .ZN(n361) );
  XNOR2_X2 U420 ( .A(G113), .B(KEYINPUT93), .ZN(n364) );
  XNOR2_X2 U421 ( .A(n365), .B(KEYINPUT35), .ZN(n788) );
  NAND2_X2 U422 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X2 U423 ( .A1(n370), .A2(n368), .ZN(n367) );
  NAND2_X1 U424 ( .A1(n599), .A2(KEYINPUT34), .ZN(n369) );
  NOR2_X1 U425 ( .A1(n787), .A2(n409), .ZN(n405) );
  NOR2_X1 U426 ( .A1(n698), .A2(n500), .ZN(n499) );
  INV_X1 U427 ( .A(G234), .ZN(n500) );
  XNOR2_X1 U428 ( .A(n644), .B(n603), .ZN(n672) );
  INV_X1 U429 ( .A(KEYINPUT38), .ZN(n603) );
  NAND2_X1 U430 ( .A1(n660), .A2(n659), .ZN(n656) );
  XNOR2_X1 U431 ( .A(n432), .B(KEYINPUT0), .ZN(n600) );
  NOR2_X1 U432 ( .A1(n729), .A2(KEYINPUT47), .ZN(n628) );
  NAND2_X1 U433 ( .A1(n490), .A2(n516), .ZN(n437) );
  NAND2_X1 U434 ( .A1(n698), .A2(n373), .ZN(n516) );
  NAND2_X1 U435 ( .A1(n351), .A2(n375), .ZN(n411) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n488) );
  NOR2_X1 U437 ( .A1(n420), .A2(n506), .ZN(n422) );
  INV_X1 U438 ( .A(n722), .ZN(n506) );
  NOR2_X1 U439 ( .A1(n602), .A2(n627), .ZN(n420) );
  NOR2_X1 U440 ( .A1(n740), .A2(n724), .ZN(n602) );
  OR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n534) );
  INV_X1 U442 ( .A(n437), .ZN(n515) );
  NAND2_X1 U443 ( .A1(n693), .A2(n380), .ZN(n514) );
  INV_X1 U444 ( .A(KEYINPUT19), .ZN(n513) );
  INV_X1 U445 ( .A(KEYINPUT1), .ZN(n431) );
  XOR2_X1 U446 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n559) );
  XNOR2_X1 U447 ( .A(n481), .B(G146), .ZN(n538) );
  INV_X1 U448 ( .A(G125), .ZN(n481) );
  XNOR2_X1 U449 ( .A(n495), .B(G101), .ZN(n562) );
  INV_X1 U450 ( .A(KEYINPUT67), .ZN(n495) );
  INV_X1 U451 ( .A(KEYINPUT87), .ZN(n428) );
  XNOR2_X1 U452 ( .A(n502), .B(n501), .ZN(n631) );
  INV_X1 U453 ( .A(KEYINPUT69), .ZN(n501) );
  INV_X1 U454 ( .A(KEYINPUT33), .ZN(n447) );
  XNOR2_X1 U455 ( .A(n663), .B(KEYINPUT6), .ZN(n635) );
  NOR2_X1 U456 ( .A1(n758), .A2(G902), .ZN(n489) );
  XNOR2_X1 U457 ( .A(KEYINPUT12), .B(KEYINPUT103), .ZN(n468) );
  XNOR2_X1 U458 ( .A(G113), .B(G131), .ZN(n581) );
  XNOR2_X1 U459 ( .A(n538), .B(n484), .ZN(n774) );
  XNOR2_X1 U460 ( .A(G140), .B(KEYINPUT10), .ZN(n484) );
  XNOR2_X1 U461 ( .A(G143), .B(G122), .ZN(n577) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(G104), .Z(n578) );
  XNOR2_X1 U463 ( .A(n470), .B(KEYINPUT104), .ZN(n469) );
  NAND2_X1 U464 ( .A1(n580), .A2(G214), .ZN(n470) );
  AND2_X1 U465 ( .A1(n657), .A2(n426), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n472), .B(n471), .ZN(n596) );
  XNOR2_X1 U467 ( .A(n584), .B(G475), .ZN(n471) );
  OR2_X1 U468 ( .A1(n751), .A2(G902), .ZN(n472) );
  INV_X1 U469 ( .A(n635), .ZN(n594) );
  BUF_X1 U470 ( .A(n660), .Z(n483) );
  XNOR2_X1 U471 ( .A(n473), .B(n387), .ZN(n592) );
  NOR2_X1 U472 ( .A1(n600), .A2(n504), .ZN(n473) );
  OR2_X1 U473 ( .A1(n673), .A2(n505), .ZN(n504) );
  INV_X1 U474 ( .A(G953), .ZN(n778) );
  NOR2_X1 U475 ( .A1(G952), .A2(n778), .ZN(n760) );
  INV_X1 U476 ( .A(KEYINPUT46), .ZN(n409) );
  INV_X1 U477 ( .A(KEYINPUT74), .ZN(n479) );
  INV_X1 U478 ( .A(KEYINPUT44), .ZN(n441) );
  INV_X1 U479 ( .A(KEYINPUT92), .ZN(n434) );
  XNOR2_X1 U480 ( .A(G902), .B(KEYINPUT15), .ZN(n533) );
  XNOR2_X1 U481 ( .A(n537), .B(n536), .ZN(n659) );
  XOR2_X1 U482 ( .A(KEYINPUT68), .B(G137), .Z(n556) );
  XNOR2_X1 U483 ( .A(n532), .B(n379), .ZN(n476) );
  NOR2_X1 U484 ( .A1(n745), .A2(n645), .ZN(n646) );
  NAND2_X1 U485 ( .A1(G237), .A2(G234), .ZN(n520) );
  NAND2_X1 U486 ( .A1(n430), .A2(n450), .ZN(n443) );
  INV_X1 U487 ( .A(n596), .ZN(n585) );
  NAND2_X1 U488 ( .A1(n515), .A2(n514), .ZN(n644) );
  NAND2_X1 U489 ( .A1(n507), .A2(n511), .ZN(n620) );
  NOR2_X1 U490 ( .A1(n512), .A2(n381), .ZN(n511) );
  INV_X1 U491 ( .A(n659), .ZN(n505) );
  XNOR2_X1 U492 ( .A(n503), .B(n425), .ZN(n424) );
  XNOR2_X1 U493 ( .A(G122), .B(KEYINPUT16), .ZN(n518) );
  XNOR2_X1 U494 ( .A(G128), .B(G119), .ZN(n539) );
  INV_X1 U495 ( .A(G143), .ZN(n528) );
  XNOR2_X1 U496 ( .A(G116), .B(G122), .ZN(n565) );
  XOR2_X1 U497 ( .A(G134), .B(G107), .Z(n566) );
  XOR2_X1 U498 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n568) );
  XOR2_X1 U499 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n543) );
  XNOR2_X1 U500 ( .A(n494), .B(n768), .ZN(n555) );
  XNOR2_X1 U501 ( .A(n562), .B(KEYINPUT71), .ZN(n494) );
  NOR2_X1 U502 ( .A1(n631), .A2(n426), .ZN(n609) );
  NAND2_X1 U503 ( .A1(n398), .A2(n371), .ZN(n397) );
  BUF_X1 U504 ( .A(n644), .Z(n482) );
  NAND2_X1 U505 ( .A1(n620), .A2(n619), .ZN(n729) );
  XNOR2_X1 U506 ( .A(n493), .B(G104), .ZN(n768) );
  XNOR2_X1 U507 ( .A(G107), .B(G110), .ZN(n493) );
  INV_X1 U508 ( .A(KEYINPUT65), .ZN(n487) );
  XNOR2_X1 U509 ( .A(n469), .B(n467), .ZN(n582) );
  XNOR2_X1 U510 ( .A(n581), .B(n468), .ZN(n467) );
  INV_X1 U511 ( .A(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U512 ( .A(n451), .B(KEYINPUT32), .ZN(n417) );
  INV_X1 U513 ( .A(KEYINPUT66), .ZN(n396) );
  XNOR2_X1 U514 ( .A(n403), .B(n402), .ZN(n401) );
  INV_X1 U515 ( .A(KEYINPUT102), .ZN(n402) );
  NAND2_X1 U516 ( .A1(n592), .A2(n657), .ZN(n593) );
  XNOR2_X1 U517 ( .A(n749), .B(n748), .ZN(n750) );
  AND2_X1 U518 ( .A1(n491), .A2(n604), .ZN(n371) );
  XOR2_X1 U519 ( .A(n555), .B(n554), .Z(n372) );
  AND2_X1 U520 ( .A1(G210), .A2(n534), .ZN(n373) );
  AND2_X1 U521 ( .A1(n728), .A2(n417), .ZN(n374) );
  AND2_X1 U522 ( .A1(n626), .A2(n733), .ZN(n375) );
  AND2_X1 U523 ( .A1(n399), .A2(n466), .ZN(n376) );
  AND2_X1 U524 ( .A1(n659), .A2(n614), .ZN(n377) );
  XNOR2_X1 U525 ( .A(G134), .B(G131), .ZN(n378) );
  XNOR2_X1 U526 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n379) );
  AND2_X1 U527 ( .A1(n699), .A2(n517), .ZN(n380) );
  NOR2_X1 U528 ( .A1(n671), .A2(n513), .ZN(n381) );
  AND2_X1 U529 ( .A1(n461), .A2(n462), .ZN(n382) );
  XOR2_X1 U530 ( .A(KEYINPUT53), .B(n692), .Z(G75) );
  NAND2_X1 U531 ( .A1(n671), .A2(n513), .ZN(n384) );
  XOR2_X1 U532 ( .A(KEYINPUT70), .B(G469), .Z(n385) );
  XOR2_X1 U533 ( .A(n618), .B(KEYINPUT39), .Z(n386) );
  XOR2_X1 U534 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n387) );
  INV_X1 U535 ( .A(KEYINPUT75), .ZN(n450) );
  XNOR2_X1 U536 ( .A(n533), .B(n434), .ZN(n698) );
  XOR2_X1 U537 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n388) );
  INV_X1 U538 ( .A(n756), .ZN(n390) );
  INV_X1 U539 ( .A(n390), .ZN(n391) );
  XNOR2_X1 U540 ( .A(n392), .B(n431), .ZN(n586) );
  AND2_X1 U541 ( .A1(n497), .A2(n392), .ZN(n619) );
  NOR2_X1 U542 ( .A1(n411), .A2(n785), .ZN(n410) );
  NAND2_X1 U543 ( .A1(n787), .A2(n409), .ZN(n407) );
  XNOR2_X1 U544 ( .A(n546), .B(n547), .ZN(n758) );
  NAND2_X1 U545 ( .A1(n393), .A2(n663), .ZN(n666) );
  OR2_X2 U546 ( .A1(n442), .A2(n444), .ZN(n393) );
  NAND2_X1 U547 ( .A1(n592), .A2(n395), .ZN(n394) );
  XNOR2_X1 U548 ( .A(n394), .B(n396), .ZN(n480) );
  INV_X1 U549 ( .A(n674), .ZN(n398) );
  XNOR2_X2 U550 ( .A(n453), .B(KEYINPUT110), .ZN(n674) );
  NAND2_X1 U551 ( .A1(n674), .A2(n492), .ZN(n399) );
  NOR2_X1 U552 ( .A1(n599), .A2(KEYINPUT34), .ZN(n400) );
  OR2_X1 U553 ( .A1(n599), .A2(n478), .ZN(n403) );
  NAND2_X1 U554 ( .A1(n406), .A2(n405), .ZN(n404) );
  INV_X1 U555 ( .A(n790), .ZN(n406) );
  NAND2_X1 U556 ( .A1(n790), .A2(n409), .ZN(n408) );
  NAND2_X1 U557 ( .A1(n414), .A2(n412), .ZN(n423) );
  NAND2_X1 U558 ( .A1(n413), .A2(n374), .ZN(n412) );
  NOR2_X1 U559 ( .A1(n788), .A2(n441), .ZN(n413) );
  NAND2_X1 U560 ( .A1(n415), .A2(n441), .ZN(n414) );
  NAND2_X1 U561 ( .A1(n416), .A2(n374), .ZN(n415) );
  INV_X1 U562 ( .A(n788), .ZN(n416) );
  XNOR2_X1 U563 ( .A(n417), .B(G119), .ZN(n789) );
  XNOR2_X2 U564 ( .A(n418), .B(n496), .ZN(n790) );
  NAND2_X1 U565 ( .A1(n477), .A2(n737), .ZN(n418) );
  XNOR2_X2 U566 ( .A(n421), .B(n388), .ZN(n697) );
  NAND2_X1 U567 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U568 ( .A(n454), .B(n424), .ZN(n713) );
  INV_X1 U569 ( .A(n560), .ZN(n425) );
  INV_X1 U570 ( .A(n663), .ZN(n426) );
  NAND2_X1 U571 ( .A1(n427), .A2(KEYINPUT2), .ZN(n647) );
  INV_X1 U572 ( .A(n429), .ZN(n427) );
  XNOR2_X1 U573 ( .A(n429), .B(n428), .ZN(n696) );
  NAND2_X1 U574 ( .A1(n620), .A2(n535), .ZN(n432) );
  NAND2_X1 U575 ( .A1(n446), .A2(n445), .ZN(n444) );
  NAND2_X1 U576 ( .A1(n435), .A2(n701), .ZN(n702) );
  NAND2_X1 U577 ( .A1(n438), .A2(n439), .ZN(n435) );
  NAND2_X1 U578 ( .A1(n586), .A2(KEYINPUT75), .ZN(n446) );
  NAND2_X1 U579 ( .A1(n508), .A2(n436), .ZN(n507) );
  NAND2_X1 U580 ( .A1(n437), .A2(n384), .ZN(n436) );
  INV_X1 U581 ( .A(n696), .ZN(n439) );
  XNOR2_X1 U582 ( .A(n563), .B(n564), .ZN(n503) );
  NOR2_X1 U583 ( .A1(n478), .A2(n616), .ZN(n440) );
  NOR2_X1 U584 ( .A1(n586), .A2(n443), .ZN(n442) );
  NAND2_X1 U585 ( .A1(n656), .A2(KEYINPUT75), .ZN(n445) );
  XNOR2_X1 U586 ( .A(n448), .B(n775), .ZN(n780) );
  XNOR2_X2 U587 ( .A(n454), .B(n449), .ZN(n448) );
  NAND2_X1 U588 ( .A1(n452), .A2(n592), .ZN(n451) );
  XNOR2_X1 U589 ( .A(n591), .B(KEYINPUT79), .ZN(n452) );
  NAND2_X1 U590 ( .A1(n672), .A2(n671), .ZN(n453) );
  XNOR2_X2 U591 ( .A(n465), .B(n378), .ZN(n454) );
  NAND2_X1 U592 ( .A1(n478), .A2(n463), .ZN(n461) );
  NAND2_X1 U593 ( .A1(n616), .A2(n463), .ZN(n462) );
  NAND2_X1 U594 ( .A1(n456), .A2(n455), .ZN(n458) );
  NAND2_X1 U595 ( .A1(n457), .A2(n382), .ZN(n623) );
  NAND2_X1 U596 ( .A1(n459), .A2(n460), .ZN(n457) );
  NOR2_X1 U597 ( .A1(n478), .A2(n463), .ZN(n459) );
  INV_X1 U598 ( .A(n616), .ZN(n460) );
  INV_X1 U599 ( .A(KEYINPUT77), .ZN(n463) );
  XNOR2_X2 U600 ( .A(n464), .B(G472), .ZN(n663) );
  XNOR2_X1 U601 ( .A(n465), .B(n555), .ZN(n474) );
  XNOR2_X2 U602 ( .A(n575), .B(KEYINPUT4), .ZN(n465) );
  INV_X1 U603 ( .A(n673), .ZN(n491) );
  NAND2_X1 U604 ( .A1(n673), .A2(n492), .ZN(n466) );
  NAND2_X1 U605 ( .A1(n477), .A2(n739), .ZN(n744) );
  XNOR2_X1 U606 ( .A(n752), .B(n753), .ZN(n754) );
  XNOR2_X1 U607 ( .A(n704), .B(n705), .ZN(n706) );
  XNOR2_X1 U608 ( .A(n708), .B(n709), .ZN(n710) );
  NAND2_X1 U609 ( .A1(n480), .A2(n587), .ZN(n728) );
  XNOR2_X2 U610 ( .A(n610), .B(n611), .ZN(n787) );
  INV_X1 U611 ( .A(n660), .ZN(n587) );
  XNOR2_X2 U612 ( .A(n529), .B(n528), .ZN(n575) );
  NAND2_X1 U613 ( .A1(n571), .A2(G221), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n542), .B(n543), .ZN(n571) );
  AND2_X2 U615 ( .A1(n486), .A2(n485), .ZN(n756) );
  INV_X1 U616 ( .A(n703), .ZN(n485) );
  XNOR2_X1 U617 ( .A(n702), .B(n487), .ZN(n486) );
  NAND2_X1 U618 ( .A1(n687), .A2(n619), .ZN(n610) );
  INV_X1 U619 ( .A(n604), .ZN(n492) );
  XNOR2_X1 U620 ( .A(n609), .B(KEYINPUT28), .ZN(n497) );
  INV_X1 U621 ( .A(n698), .ZN(n699) );
  NAND2_X1 U622 ( .A1(n548), .A2(G217), .ZN(n549) );
  XNOR2_X1 U623 ( .A(n499), .B(n498), .ZN(n548) );
  INV_X1 U624 ( .A(KEYINPUT20), .ZN(n498) );
  NAND2_X1 U625 ( .A1(n377), .A2(n587), .ZN(n502) );
  NAND2_X1 U626 ( .A1(n663), .A2(n671), .ZN(n613) );
  NAND2_X1 U627 ( .A1(n515), .A2(n509), .ZN(n508) );
  INV_X1 U628 ( .A(n514), .ZN(n510) );
  NOR2_X1 U629 ( .A1(n514), .A2(n384), .ZN(n512) );
  INV_X1 U630 ( .A(n373), .ZN(n517) );
  XNOR2_X1 U631 ( .A(n653), .B(KEYINPUT82), .ZN(n654) );
  BUF_X1 U632 ( .A(n697), .Z(n761) );
  XNOR2_X1 U633 ( .A(n562), .B(n561), .ZN(n563) );
  INV_X1 U634 ( .A(KEYINPUT30), .ZN(n612) );
  INV_X1 U635 ( .A(n679), .ZN(n686) );
  INV_X1 U636 ( .A(KEYINPUT72), .ZN(n618) );
  XNOR2_X1 U637 ( .A(n520), .B(KEYINPUT14), .ZN(n523) );
  NAND2_X1 U638 ( .A1(G952), .A2(n523), .ZN(n685) );
  NOR2_X1 U639 ( .A1(n685), .A2(G953), .ZN(n521) );
  XOR2_X1 U640 ( .A(n521), .B(KEYINPUT94), .Z(n608) );
  INV_X1 U641 ( .A(n608), .ZN(n526) );
  NOR2_X1 U642 ( .A1(G898), .A2(n778), .ZN(n522) );
  XNOR2_X1 U643 ( .A(KEYINPUT95), .B(n522), .ZN(n771) );
  NAND2_X1 U644 ( .A1(G902), .A2(n523), .ZN(n605) );
  NOR2_X1 U645 ( .A1(n771), .A2(n605), .ZN(n524) );
  XNOR2_X1 U646 ( .A(n524), .B(KEYINPUT96), .ZN(n525) );
  NOR2_X1 U647 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U648 ( .A(KEYINPUT97), .B(n527), .ZN(n535) );
  XNOR2_X2 U649 ( .A(G128), .B(KEYINPUT81), .ZN(n529) );
  XNOR2_X1 U650 ( .A(G119), .B(KEYINPUT3), .ZN(n530) );
  XNOR2_X1 U651 ( .A(n538), .B(KEYINPUT17), .ZN(n531) );
  NAND2_X1 U652 ( .A1(G224), .A2(n778), .ZN(n532) );
  NAND2_X1 U653 ( .A1(G214), .A2(n534), .ZN(n671) );
  XNOR2_X1 U654 ( .A(n600), .B(KEYINPUT98), .ZN(n599) );
  XOR2_X1 U655 ( .A(KEYINPUT21), .B(KEYINPUT100), .Z(n537) );
  NAND2_X1 U656 ( .A1(n548), .A2(G221), .ZN(n536) );
  XOR2_X1 U657 ( .A(KEYINPUT24), .B(G110), .Z(n540) );
  XNOR2_X1 U658 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U659 ( .A(n774), .B(n541), .ZN(n547) );
  XOR2_X1 U660 ( .A(n556), .B(KEYINPUT23), .Z(n545) );
  NAND2_X1 U661 ( .A1(G234), .A2(n778), .ZN(n542) );
  XNOR2_X1 U662 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U663 ( .A(KEYINPUT99), .B(KEYINPUT25), .Z(n550) );
  XNOR2_X1 U664 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U665 ( .A1(G227), .A2(n778), .ZN(n552) );
  XNOR2_X1 U666 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U667 ( .A1(n580), .A2(G210), .ZN(n558) );
  XNOR2_X1 U668 ( .A(n559), .B(n558), .ZN(n564) );
  XOR2_X1 U669 ( .A(G146), .B(G137), .Z(n561) );
  XNOR2_X1 U670 ( .A(n566), .B(n565), .ZN(n570) );
  XNOR2_X1 U671 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n567) );
  XNOR2_X1 U672 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U673 ( .A(n570), .B(n569), .Z(n573) );
  NAND2_X1 U674 ( .A1(G217), .A2(n571), .ZN(n572) );
  XNOR2_X1 U675 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U676 ( .A(n575), .B(n574), .ZN(n709) );
  NOR2_X1 U677 ( .A1(G902), .A2(n709), .ZN(n576) );
  XNOR2_X1 U678 ( .A(n576), .B(G478), .ZN(n597) );
  XNOR2_X1 U679 ( .A(KEYINPUT105), .B(KEYINPUT13), .ZN(n584) );
  XNOR2_X1 U680 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U681 ( .A(n774), .B(n579), .ZN(n583) );
  XNOR2_X1 U682 ( .A(n583), .B(n582), .ZN(n751) );
  NOR2_X1 U683 ( .A1(n597), .A2(n585), .ZN(n622) );
  NAND2_X1 U684 ( .A1(n597), .A2(n585), .ZN(n673) );
  NOR2_X1 U685 ( .A1(n483), .A2(n657), .ZN(n588) );
  XNOR2_X1 U686 ( .A(n588), .B(KEYINPUT108), .ZN(n590) );
  XOR2_X1 U687 ( .A(n594), .B(KEYINPUT80), .Z(n589) );
  NAND2_X1 U688 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U689 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U690 ( .A1(n595), .A2(n483), .ZN(n722) );
  NAND2_X1 U691 ( .A1(n596), .A2(n597), .ZN(n632) );
  INV_X1 U692 ( .A(n632), .ZN(n737) );
  NOR2_X1 U693 ( .A1(n597), .A2(n596), .ZN(n739) );
  NOR2_X1 U694 ( .A1(n737), .A2(n739), .ZN(n675) );
  XOR2_X1 U695 ( .A(KEYINPUT83), .B(n675), .Z(n627) );
  NOR2_X1 U696 ( .A1(n600), .A2(n666), .ZN(n601) );
  XOR2_X1 U697 ( .A(KEYINPUT31), .B(n601), .Z(n740) );
  XOR2_X1 U698 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n611) );
  XNOR2_X1 U699 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n604) );
  NOR2_X1 U700 ( .A1(G900), .A2(n605), .ZN(n606) );
  NAND2_X1 U701 ( .A1(G953), .A2(n606), .ZN(n607) );
  NAND2_X1 U702 ( .A1(n608), .A2(n607), .ZN(n614) );
  INV_X1 U703 ( .A(n672), .ZN(n617) );
  XNOR2_X1 U704 ( .A(n613), .B(n612), .ZN(n615) );
  NAND2_X1 U705 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U706 ( .A1(n729), .A2(n675), .ZN(n621) );
  NAND2_X1 U707 ( .A1(KEYINPUT47), .A2(n621), .ZN(n626) );
  INV_X1 U708 ( .A(n622), .ZN(n624) );
  NOR2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n482), .A2(n625), .ZN(n733) );
  INV_X1 U711 ( .A(n627), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n633), .A2(n671), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n640) );
  AND2_X1 U716 ( .A1(n482), .A2(n640), .ZN(n636) );
  XNOR2_X1 U717 ( .A(KEYINPUT36), .B(n636), .ZN(n638) );
  INV_X1 U718 ( .A(n657), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT113), .ZN(n785) );
  NAND2_X1 U721 ( .A1(n657), .A2(n640), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n641), .B(KEYINPUT109), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(KEYINPUT43), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n482), .A2(n643), .ZN(n745) );
  INV_X1 U725 ( .A(n744), .ZN(n645) );
  XNOR2_X1 U726 ( .A(KEYINPUT88), .B(n647), .ZN(n648) );
  NOR2_X1 U727 ( .A1(n761), .A2(n648), .ZN(n703) );
  INV_X1 U728 ( .A(KEYINPUT2), .ZN(n650) );
  AND2_X1 U729 ( .A1(n650), .A2(n697), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT85), .ZN(n652) );
  BUF_X1 U731 ( .A(n696), .Z(n777) );
  NAND2_X1 U732 ( .A1(n650), .A2(n777), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U734 ( .A1(n703), .A2(n654), .ZN(n655) );
  NOR2_X1 U735 ( .A1(G953), .A2(n655), .ZN(n691) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(KEYINPUT50), .ZN(n665) );
  NOR2_X1 U738 ( .A1(n483), .A2(n659), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT49), .B(n661), .Z(n662) );
  NOR2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n669) );
  XOR2_X1 U743 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n668) );
  XNOR2_X1 U744 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n670), .A2(n687), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n673), .A2(n353), .ZN(n677) );
  NOR2_X1 U747 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U749 ( .A(KEYINPUT121), .B(n678), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n680), .A2(n686), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U752 ( .A(KEYINPUT52), .B(n683), .Z(n684) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n689) );
  AND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U757 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n695) );
  XNOR2_X1 U758 ( .A(n693), .B(KEYINPUT89), .ZN(n694) );
  XNOR2_X1 U759 ( .A(n695), .B(n694), .ZN(n705) );
  XOR2_X1 U760 ( .A(n699), .B(KEYINPUT86), .Z(n700) );
  NAND2_X1 U761 ( .A1(n700), .A2(KEYINPUT2), .ZN(n701) );
  NAND2_X1 U762 ( .A1(n756), .A2(G210), .ZN(n704) );
  NOR2_X2 U763 ( .A1(n706), .A2(n760), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n707), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U765 ( .A1(n756), .A2(G478), .ZN(n708) );
  NOR2_X2 U766 ( .A1(n710), .A2(n760), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT122), .ZN(G63) );
  INV_X1 U768 ( .A(n760), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n756), .A2(G472), .ZN(n715) );
  XOR2_X1 U770 ( .A(KEYINPUT62), .B(KEYINPUT90), .Z(n712) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U772 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U773 ( .A(KEYINPUT63), .B(KEYINPUT114), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n718), .B(KEYINPUT91), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(G57) );
  XOR2_X1 U776 ( .A(G101), .B(KEYINPUT115), .Z(n721) );
  XNOR2_X1 U777 ( .A(n722), .B(n721), .ZN(G3) );
  NAND2_X1 U778 ( .A1(n737), .A2(n724), .ZN(n723) );
  XNOR2_X1 U779 ( .A(G104), .B(n723), .ZN(G6) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n726) );
  NAND2_X1 U781 ( .A1(n724), .A2(n739), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U783 ( .A(G107), .B(n727), .ZN(G9) );
  XNOR2_X1 U784 ( .A(n728), .B(G110), .ZN(G12) );
  XOR2_X1 U785 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n731) );
  INV_X1 U786 ( .A(n729), .ZN(n734) );
  NAND2_X1 U787 ( .A1(n734), .A2(n739), .ZN(n730) );
  XNOR2_X1 U788 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U789 ( .A(G128), .B(n732), .ZN(G30) );
  XNOR2_X1 U790 ( .A(G143), .B(n733), .ZN(G45) );
  XOR2_X1 U791 ( .A(G146), .B(KEYINPUT117), .Z(n736) );
  NAND2_X1 U792 ( .A1(n734), .A2(n737), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(G48) );
  NAND2_X1 U794 ( .A1(n740), .A2(n737), .ZN(n738) );
  XNOR2_X1 U795 ( .A(n738), .B(G113), .ZN(G15) );
  NAND2_X1 U796 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U797 ( .A(n741), .B(KEYINPUT118), .ZN(n742) );
  XNOR2_X1 U798 ( .A(G116), .B(n742), .ZN(G18) );
  XOR2_X1 U799 ( .A(G134), .B(KEYINPUT119), .Z(n743) );
  XNOR2_X1 U800 ( .A(n744), .B(n743), .ZN(G36) );
  XOR2_X1 U801 ( .A(G140), .B(n745), .Z(G42) );
  NAND2_X1 U802 ( .A1(n391), .A2(G469), .ZN(n749) );
  XOR2_X1 U803 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n746) );
  XNOR2_X1 U804 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U805 ( .A1(n760), .A2(n750), .ZN(G54) );
  XOR2_X1 U806 ( .A(n751), .B(KEYINPUT59), .Z(n753) );
  NAND2_X1 U807 ( .A1(n756), .A2(G475), .ZN(n752) );
  NOR2_X2 U808 ( .A1(n754), .A2(n760), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U810 ( .A1(G217), .A2(n391), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U812 ( .A1(n760), .A2(n759), .ZN(G66) );
  NOR2_X1 U813 ( .A1(G953), .A2(n761), .ZN(n762) );
  XNOR2_X1 U814 ( .A(n762), .B(KEYINPUT123), .ZN(n766) );
  NAND2_X1 U815 ( .A1(G953), .A2(G224), .ZN(n763) );
  XNOR2_X1 U816 ( .A(KEYINPUT61), .B(n763), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n764), .A2(G898), .ZN(n765) );
  NAND2_X1 U818 ( .A1(n766), .A2(n765), .ZN(n773) );
  XNOR2_X1 U819 ( .A(n767), .B(G101), .ZN(n769) );
  XNOR2_X1 U820 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U821 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U822 ( .A(n773), .B(n772), .Z(G69) );
  XNOR2_X1 U823 ( .A(n774), .B(KEYINPUT124), .ZN(n775) );
  XOR2_X1 U824 ( .A(KEYINPUT125), .B(n780), .Z(n776) );
  XNOR2_X1 U825 ( .A(n777), .B(n776), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n779), .A2(n778), .ZN(n784) );
  XNOR2_X1 U827 ( .A(G227), .B(n780), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U829 ( .A1(n782), .A2(G953), .ZN(n783) );
  NAND2_X1 U830 ( .A1(n784), .A2(n783), .ZN(G72) );
  XNOR2_X1 U831 ( .A(G125), .B(n785), .ZN(n786) );
  XNOR2_X1 U832 ( .A(n786), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U833 ( .A(n787), .B(G137), .Z(G39) );
  XOR2_X1 U834 ( .A(n788), .B(G122), .Z(G24) );
  XNOR2_X1 U835 ( .A(n789), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U836 ( .A(n790), .B(G131), .Z(G33) );
endmodule

