//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT72), .B(G902), .Z(new_n193));
  AOI211_X1 g007(.A(new_n187), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT21), .B(G898), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G902), .ZN(new_n197));
  XNOR2_X1  g011(.A(G113), .B(G122), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT16), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(KEYINPUT16), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n202), .B(G146), .C1(KEYINPUT16), .C2(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(G237), .A2(G953), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(G143), .A3(G214), .ZN(new_n212));
  AOI21_X1  g026(.A(G143), .B1(new_n211), .B2(G214), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT17), .A3(G131), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n212), .A2(new_n213), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n210), .B(new_n215), .C1(KEYINPUT17), .C2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(KEYINPUT18), .A3(G131), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n216), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n201), .B(new_n206), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n200), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n207), .A3(new_n208), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n200), .B(new_n224), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n197), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G475), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT20), .ZN(new_n232));
  XOR2_X1   g046(.A(new_n201), .B(KEYINPUT19), .Z(new_n233));
  OAI211_X1 g047(.A(new_n218), .B(new_n208), .C1(G146), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n224), .ZN(new_n235));
  INV_X1    g049(.A(new_n200), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n228), .ZN(new_n238));
  NOR2_X1   g052(.A1(G475), .A2(G902), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  AOI211_X1 g055(.A(KEYINPUT20), .B(new_n241), .C1(new_n237), .C2(new_n228), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n231), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G122), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT14), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT94), .Z(new_n247));
  INV_X1    g061(.A(G122), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G116), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n245), .B2(KEYINPUT14), .ZN(new_n250));
  OAI21_X1  g064(.A(G107), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n249), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G107), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G128), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G134), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n255), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(KEYINPUT93), .A2(new_n253), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n251), .B(new_n262), .C1(KEYINPUT93), .C2(new_n253), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT9), .B(G234), .Z(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT78), .ZN(new_n265));
  INV_X1    g079(.A(G217), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n265), .A2(new_n266), .A3(G953), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT13), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n257), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n255), .A2(new_n268), .ZN(new_n271));
  OAI21_X1  g085(.A(G134), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n273), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n252), .B(G107), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n274), .A2(new_n261), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n263), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n267), .B1(new_n263), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n193), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G478), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(KEYINPUT15), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n263), .A2(new_n277), .ZN(new_n285));
  INV_X1    g099(.A(new_n267), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n278), .ZN(new_n288));
  INV_X1    g102(.A(new_n283), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n193), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(KEYINPUT95), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT95), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n288), .B2(new_n193), .ZN(new_n293));
  INV_X1    g107(.A(new_n193), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n283), .C1(new_n287), .C2(new_n278), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n196), .B(new_n243), .C1(new_n291), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n244), .B2(G119), .ZN(new_n300));
  INV_X1    g114(.A(G119), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT68), .A3(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n244), .A2(G119), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G113), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n308), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n310), .A2(new_n300), .A3(new_n302), .A4(new_n303), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(new_n199), .B2(G107), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n316), .A2(new_n199), .A3(G107), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n318), .A2(G104), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G101), .ZN(new_n322));
  INV_X1    g136(.A(G101), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n323), .B(new_n315), .C1(new_n317), .C2(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n316), .B1(new_n199), .B2(G107), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n318), .A2(KEYINPUT79), .A3(KEYINPUT3), .A4(G104), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n328), .B2(new_n315), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n312), .B(new_n322), .C1(new_n325), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n199), .A2(G107), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n318), .A2(G104), .ZN(new_n332));
  OAI21_X1  g146(.A(G101), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n244), .A2(G119), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n305), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n304), .B2(new_n336), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n311), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G122), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT87), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n330), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n206), .A2(G143), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n254), .A2(G146), .ZN(new_n348));
  AND2_X1   g162(.A1(KEYINPUT0), .A2(G128), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G143), .B(G146), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G128), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT88), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n348), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n206), .A2(G143), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n356), .A2(new_n256), .B1(KEYINPUT1), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT1), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n347), .A2(new_n348), .A3(new_n359), .A4(G128), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n203), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT88), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n353), .A2(new_n362), .A3(G125), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n355), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G224), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n364), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n340), .A2(new_n368), .A3(new_n342), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n346), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT89), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n346), .A2(new_n367), .A3(new_n372), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n345), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT7), .B1(new_n365), .B2(G953), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n364), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n355), .A2(new_n361), .A3(new_n363), .A4(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n342), .B(KEYINPUT8), .Z(new_n381));
  NAND2_X1  g195(.A1(new_n338), .A2(new_n311), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n324), .A2(new_n333), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n339), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n375), .B1(new_n387), .B2(KEYINPUT90), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n380), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G902), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n374), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G210), .B1(G237), .B2(G902), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n374), .A2(new_n391), .A3(new_n393), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(KEYINPUT91), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n298), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n266), .B1(new_n193), .B2(G234), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n201), .A2(new_n206), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n301), .A2(G128), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n301), .A2(G128), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(KEYINPUT23), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(G110), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n411));
  XNOR2_X1  g225(.A(G119), .B(G128), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT24), .B(G110), .Z(new_n413));
  OAI22_X1  g227(.A1(new_n410), .A2(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n208), .B(new_n405), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G110), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n418), .B2(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n412), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n209), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT77), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT22), .B(G137), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n416), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n416), .B2(new_n423), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT25), .A3(new_n193), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT25), .B1(new_n430), .B2(new_n193), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n404), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n404), .A2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT65), .ZN(new_n438));
  INV_X1    g252(.A(G137), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(G134), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n260), .A2(KEYINPUT65), .A3(G137), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n260), .A2(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(G134), .ZN(new_n446));
  NOR2_X1   g260(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(new_n443), .ZN(new_n449));
  OAI21_X1  g263(.A(G131), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n439), .A2(G134), .ZN(new_n451));
  AOI22_X1  g265(.A1(KEYINPUT65), .A2(new_n451), .B1(new_n446), .B2(new_n443), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n442), .B1(new_n444), .B2(new_n447), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n217), .A4(new_n440), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n353), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n446), .A2(KEYINPUT66), .ZN(new_n457));
  INV_X1    g271(.A(new_n451), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n439), .A3(G134), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n358), .A2(new_n360), .B1(new_n461), .B2(G131), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n455), .A2(new_n456), .B1(new_n462), .B2(new_n454), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT67), .B1(new_n463), .B2(KEYINPUT30), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT69), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n350), .B(new_n465), .C1(new_n351), .C2(new_n352), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n455), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n454), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n358), .A2(new_n360), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n461), .A2(G131), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n473), .A2(new_n454), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n353), .B1(new_n450), .B2(new_n454), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n471), .B(new_n472), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n464), .A2(new_n312), .A3(new_n470), .A4(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n312), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n450), .A2(new_n454), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n467), .A2(new_n466), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n469), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n190), .A2(new_n187), .A3(G210), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT26), .B(G101), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n478), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT31), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n482), .A2(KEYINPUT28), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n468), .A2(new_n491), .A3(new_n479), .A4(new_n469), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n312), .B1(new_n475), .B2(new_n476), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n487), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n478), .A2(new_n498), .A3(new_n482), .A4(new_n487), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(G472), .A2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n487), .A2(KEYINPUT29), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n479), .B1(new_n468), .B2(new_n469), .ZN(new_n509));
  AOI211_X1 g323(.A(new_n508), .B(new_n509), .C1(new_n490), .C2(new_n492), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT73), .B1(new_n510), .B2(new_n294), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n490), .B2(new_n492), .ZN(new_n512));
  INV_X1    g326(.A(new_n508), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n193), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n495), .A2(new_n487), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n482), .A2(new_n496), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n478), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT29), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G472), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n501), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n437), .B1(new_n507), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G110), .B(G140), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n187), .A2(G227), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n473), .A2(KEYINPUT10), .A3(new_n324), .A4(new_n333), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n322), .A2(new_n467), .A3(new_n466), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n325), .A2(new_n329), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(G128), .B1(new_n347), .B2(new_n348), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n348), .A2(new_n359), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT81), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n357), .A2(KEYINPUT1), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT81), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(new_n351), .C2(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n360), .A2(KEYINPUT80), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n351), .A2(new_n540), .A3(new_n359), .A4(G128), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n535), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT10), .B1(new_n542), .B2(new_n334), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n532), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT82), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n480), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n334), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT10), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n320), .A2(G101), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n466), .A3(new_n467), .A4(new_n322), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n549), .A2(new_n480), .A3(new_n552), .A4(new_n529), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT82), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n528), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n549), .A2(new_n552), .A3(new_n529), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n480), .B1(new_n556), .B2(KEYINPUT83), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT83), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n549), .A2(new_n558), .A3(new_n552), .A4(new_n529), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT84), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT83), .B1(new_n532), .B2(new_n543), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n561), .A2(new_n559), .A3(KEYINPUT84), .A4(new_n455), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n555), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n383), .A2(new_n358), .A3(new_n360), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n480), .B1(new_n547), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT12), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n545), .B1(new_n544), .B2(new_n480), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n553), .A2(KEYINPUT82), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n528), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n564), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G469), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT85), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT85), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n561), .A2(new_n559), .A3(new_n455), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT84), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n562), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(new_n555), .B1(new_n570), .B2(new_n528), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n575), .B(G469), .C1(new_n580), .C2(G902), .ZN(new_n581));
  INV_X1    g395(.A(new_n528), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n546), .A2(new_n554), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n555), .A2(new_n567), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n573), .B(new_n193), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n574), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n588));
  OAI21_X1  g402(.A(G221), .B1(new_n265), .B2(G902), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n403), .B(new_n525), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n589), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT86), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n395), .A2(new_n396), .ZN(new_n598));
  INV_X1    g412(.A(new_n196), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n401), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n294), .A2(new_n282), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n279), .A2(KEYINPUT33), .A3(new_n280), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n287), .B2(new_n278), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n281), .A2(new_n282), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n243), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n504), .A2(new_n506), .ZN(new_n610));
  INV_X1    g424(.A(new_n437), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n500), .A2(new_n193), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n597), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n242), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n240), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n238), .A2(KEYINPUT96), .A3(new_n232), .A4(new_n239), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n622), .A2(new_n291), .A3(new_n296), .A4(new_n231), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n600), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n597), .A2(new_n614), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n416), .A2(new_n423), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n427), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n435), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n434), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n504), .A2(new_n632), .A3(new_n613), .A4(new_n506), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n403), .B(new_n633), .C1(new_n590), .C2(new_n591), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  INV_X1    g451(.A(G900), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n192), .B1(new_n194), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n623), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n402), .B1(new_n395), .B2(new_n396), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n632), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n507), .B2(new_n524), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n642), .B(new_n644), .C1(new_n590), .C2(new_n591), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XOR2_X1   g460(.A(new_n639), .B(KEYINPUT39), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n597), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n400), .A2(KEYINPUT38), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n397), .A2(new_n652), .A3(new_n399), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n296), .A2(new_n291), .A3(new_n243), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n401), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n519), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n197), .B1(new_n657), .B2(new_n509), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n496), .B1(new_n478), .B2(new_n482), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n507), .A2(new_n523), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n656), .A2(new_n632), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n649), .A2(new_n650), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  INV_X1    g479(.A(new_n639), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n607), .A2(new_n243), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n641), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n644), .B(new_n669), .C1(new_n590), .C2(new_n591), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  OAI21_X1  g485(.A(new_n193), .B1(new_n584), .B2(new_n585), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G469), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n673), .A2(new_n589), .A3(new_n586), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n609), .A2(new_n525), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND3_X1  g491(.A1(new_n624), .A2(new_n525), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND4_X1  g493(.A1(new_n644), .A2(new_n674), .A3(new_n297), .A4(new_n641), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  INV_X1    g495(.A(new_n600), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n489), .B(new_n499), .C1(new_n512), .C2(new_n487), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n501), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n436), .A2(new_n613), .A3(new_n434), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n674), .A2(new_n682), .A3(new_n685), .A4(new_n655), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  AND4_X1   g501(.A1(new_n613), .A2(new_n632), .A3(new_n667), .A4(new_n684), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n674), .A3(new_n641), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  INV_X1    g504(.A(new_n589), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n402), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n397), .B2(new_n399), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n580), .B2(G902), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n586), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT98), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n586), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n694), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n522), .A2(new_n523), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT32), .B1(new_n500), .B2(new_n501), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n611), .B(new_n667), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT42), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n586), .A2(new_n695), .A3(new_n698), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n698), .B1(new_n586), .B2(new_n695), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n667), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(KEYINPUT42), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n525), .A3(new_n694), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n217), .ZN(G33));
  NAND4_X1  g526(.A1(new_n707), .A2(new_n525), .A3(new_n640), .A4(new_n694), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT99), .B(G134), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G36));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n580), .A2(KEYINPUT45), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n580), .A2(KEYINPUT45), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n573), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n573), .A2(new_n197), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n721), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n725), .B(KEYINPUT46), .C1(new_n573), .C2(new_n197), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n586), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(new_n589), .ZN(new_n728));
  INV_X1    g542(.A(new_n607), .ZN(new_n729));
  OR3_X1    g543(.A1(new_n729), .A2(KEYINPUT43), .A3(new_n243), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n729), .B2(new_n243), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n730), .A2(new_n632), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n610), .A2(new_n613), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n402), .B1(new_n397), .B2(new_n399), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n728), .A2(new_n647), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  NAND2_X1  g554(.A1(new_n728), .A2(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n727), .A2(new_n589), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n507), .A2(new_n524), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n737), .A2(new_n746), .A3(new_n708), .A4(new_n611), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  NOR4_X1   g563(.A1(new_n437), .A2(new_n243), .A3(new_n729), .A4(new_n693), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT101), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n673), .A2(new_n586), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n751), .B1(KEYINPUT49), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(KEYINPUT49), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT102), .ZN(new_n756));
  INV_X1    g570(.A(new_n654), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n756), .A3(new_n662), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT107), .B(KEYINPUT51), .ZN(new_n759));
  INV_X1    g573(.A(new_n674), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n737), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n730), .A2(new_n192), .A3(new_n731), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT110), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(KEYINPUT110), .A3(new_n762), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n613), .A2(new_n684), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n632), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT111), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n771), .B(new_n768), .C1(new_n764), .C2(new_n765), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n762), .A2(new_n685), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n654), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n674), .B2(new_n402), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n760), .A2(KEYINPUT109), .A3(new_n401), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n775), .B(KEYINPUT50), .C1(new_n778), .C2(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n761), .A2(new_n611), .A3(new_n192), .A4(new_n662), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n607), .A2(new_n243), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT113), .B1(new_n773), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n774), .A2(new_n737), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n752), .A2(new_n691), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT108), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n745), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n773), .A2(new_n789), .A3(KEYINPUT113), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n759), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n741), .A2(new_n744), .A3(new_n792), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT115), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n741), .A2(new_n800), .A3(new_n744), .A4(new_n792), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n801), .A3(new_n791), .ZN(new_n802));
  INV_X1    g616(.A(new_n789), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n766), .A2(new_n769), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n771), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n769), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT114), .B1(new_n773), .B2(new_n789), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n802), .A2(new_n809), .A3(new_n810), .A4(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n674), .A2(new_n641), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n188), .B1(new_n774), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n611), .B1(new_n701), .B2(new_n702), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n766), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n608), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n784), .B(KEYINPUT112), .Z(new_n820));
  AOI211_X1 g634(.A(new_n813), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n797), .A2(new_n811), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n680), .A2(new_n675), .A3(new_n678), .A4(new_n686), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n711), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n707), .A2(new_n688), .A3(new_n694), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n713), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n746), .A2(new_n632), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n595), .B2(new_n596), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n284), .A2(new_n290), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n639), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(new_n231), .A3(new_n622), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n736), .A2(KEYINPUT104), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT104), .B1(new_n736), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n827), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  OAI221_X1 g650(.A(new_n403), .B1(new_n525), .B2(new_n633), .C1(new_n590), .C2(new_n591), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n830), .B(new_n231), .C1(new_n240), .C2(new_n242), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n196), .B1(new_n608), .B2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n401), .A2(new_n839), .A3(new_n399), .A4(new_n397), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n614), .B(new_n840), .C1(new_n590), .C2(new_n591), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n837), .A2(KEYINPUT103), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT103), .B1(new_n837), .B2(new_n841), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n825), .B(new_n836), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n689), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n829), .B2(new_n642), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n589), .A2(new_n641), .A3(new_n666), .A4(new_n655), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n707), .A3(new_n643), .A4(new_n661), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n670), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n645), .A2(new_n670), .A3(new_n689), .A4(new_n849), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n823), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n844), .A2(new_n853), .A3(new_n823), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT54), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n829), .A2(new_n835), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n713), .A2(new_n826), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT53), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n592), .A2(new_n634), .A3(new_n841), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n837), .A2(KEYINPUT103), .A3(new_n841), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n675), .A2(new_n680), .A3(new_n678), .A4(new_n686), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n704), .A2(new_n710), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT106), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT106), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n824), .B2(new_n711), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n852), .A3(new_n871), .A4(new_n850), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n854), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n857), .A2(KEYINPUT105), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT105), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n876), .B(KEYINPUT54), .C1(new_n855), .C2(new_n856), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n822), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n758), .B1(new_n878), .B2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n854), .A2(new_n872), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n193), .A2(new_n393), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n346), .A2(new_n369), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n367), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n883), .A2(new_n887), .B1(G952), .B2(new_n187), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n883), .B2(KEYINPUT117), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n881), .A2(KEYINPUT117), .A3(new_n882), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n886), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n888), .B1(new_n893), .B2(new_n895), .ZN(G51));
  NOR2_X1   g710(.A1(new_n187), .A2(G952), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n874), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n881), .A2(new_n900), .A3(KEYINPUT54), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n723), .B(KEYINPUT57), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n584), .B2(new_n585), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n193), .B1(new_n854), .B2(new_n872), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n722), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n897), .B1(new_n904), .B2(new_n906), .ZN(G54));
  AND3_X1   g721(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n238), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n238), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n897), .ZN(G60));
  OR2_X1    g725(.A1(new_n602), .A2(new_n604), .ZN(new_n912));
  XOR2_X1   g726(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n282), .A2(new_n197), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n899), .A2(new_n901), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT121), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n899), .A2(new_n919), .A3(new_n901), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n875), .A2(new_n877), .A3(new_n915), .ZN(new_n922));
  INV_X1    g736(.A(new_n912), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n897), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n921), .A2(new_n924), .ZN(G63));
  XOR2_X1   g739(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n266), .A2(new_n197), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n430), .B1(new_n881), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n897), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n881), .A2(new_n630), .A3(new_n929), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n931), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n926), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  INV_X1    g753(.A(new_n195), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n187), .B1(new_n940), .B2(G224), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n824), .B1(new_n863), .B2(new_n864), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n943), .B2(new_n187), .ZN(new_n944));
  INV_X1    g758(.A(G898), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n884), .B1(new_n945), .B2(G953), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G69));
  AND2_X1   g761(.A1(new_n748), .A2(new_n739), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n846), .A2(new_n670), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n664), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n952));
  INV_X1    g766(.A(new_n525), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n608), .A2(new_n838), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n648), .A2(new_n953), .A3(new_n737), .A4(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n948), .A2(new_n951), .A3(new_n952), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n187), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n464), .A2(new_n470), .A3(new_n477), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n233), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n815), .A2(new_n641), .A3(new_n655), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n728), .B(new_n647), .C1(new_n738), .C2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n867), .A2(new_n713), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n748), .A3(new_n949), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n969), .A2(new_n748), .A3(new_n972), .A4(new_n949), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n964), .B1(new_n974), .B2(G953), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n963), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n963), .A2(new_n975), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n974), .B2(new_n943), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n478), .A3(new_n519), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n958), .B2(new_n943), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n897), .B1(new_n988), .B2(new_n659), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n520), .A2(new_n985), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n659), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n855), .B2(new_n856), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n987), .A2(new_n989), .A3(new_n992), .ZN(G57));
endmodule


