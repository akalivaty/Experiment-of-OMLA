//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n217), .B2(new_n218), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n208), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(new_n207), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(KEYINPUT18), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n208), .B(new_n220), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n226), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(G197gat), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT11), .B(G169gat), .Z(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(KEYINPUT12), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n228), .A2(new_n240), .A3(new_n229), .A4(new_n232), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n244));
  AND2_X1   g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G155gat), .ZN(new_n248));
  INV_X1    g047(.A(G162gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(KEYINPUT78), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G141gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G148gat), .ZN(new_n255));
  INV_X1    g054(.A(G148gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G141gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT79), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(G155gat), .B2(G162gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n257), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n253), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(G141gat), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n255), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n251), .B1(new_n250), .B2(KEYINPUT2), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT81), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n256), .A2(G141gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n254), .A2(G148gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n262), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n260), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n258), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n247), .A2(new_n252), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n268), .A2(new_n269), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n271), .A2(KEYINPUT3), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g088(.A(G127gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(G134gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G127gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(G134gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT70), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n286), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n294), .A2(new_n295), .A3(new_n288), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n292), .A2(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n276), .A2(new_n277), .B1(new_n268), .B2(new_n269), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n282), .A2(new_n305), .ZN(new_n306));
  AND4_X1   g105(.A1(KEYINPUT4), .A2(new_n302), .A3(new_n278), .A4(new_n280), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT4), .B1(new_n303), .B2(new_n302), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n306), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT83), .ZN(new_n313));
  INV_X1    g112(.A(new_n311), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n307), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(new_n316), .A3(new_n306), .A4(new_n310), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n319));
  INV_X1    g118(.A(new_n302), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n271), .A2(new_n281), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n302), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n314), .ZN(new_n324));
  AND4_X1   g123(.A1(KEYINPUT82), .A2(new_n319), .A3(KEYINPUT5), .A4(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n310), .B1(new_n315), .B2(new_n306), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT82), .B1(new_n326), .B2(new_n324), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n318), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT0), .ZN(new_n330));
  XNOR2_X1  g129(.A(G57gat), .B(G85gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(KEYINPUT6), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n313), .B2(new_n317), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n327), .B2(new_n325), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n319), .A2(KEYINPUT5), .A3(new_n324), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n324), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n332), .B1(new_n343), .B2(new_n318), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n334), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348));
  AND2_X1   g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n347), .A2(new_n348), .B1(new_n349), .B2(KEYINPUT22), .ZN(new_n350));
  NOR2_X1   g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G197gat), .ZN(new_n355));
  INV_X1    g154(.A(G204gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358));
  NAND2_X1  g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n357), .A2(new_n346), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  INV_X1    g160(.A(G218gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT76), .A3(new_n359), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371));
  INV_X1    g170(.A(G169gat), .ZN(new_n372));
  INV_X1    g171(.A(G176gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT26), .ZN(new_n374));
  NAND2_X1  g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n371), .B(new_n374), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n378), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n382), .B(KEYINPUT69), .C1(new_n378), .C2(new_n377), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n385));
  OR2_X1    g184(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(KEYINPUT28), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G183gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT27), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT27), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G183gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n385), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n387), .ZN(new_n395));
  NOR2_X1   g194(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT27), .B(G183gat), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT68), .A4(KEYINPUT28), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n391), .B1(new_n389), .B2(KEYINPUT66), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(KEYINPUT64), .A3(KEYINPUT27), .A4(G183gat), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n401), .B(new_n403), .C1(KEYINPUT64), .C2(G183gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n397), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n384), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n371), .A2(KEYINPUT24), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(G183gat), .A3(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n386), .A2(new_n387), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT64), .B(G183gat), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n378), .A2(KEYINPUT23), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(G169gat), .B2(G176gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n375), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n420), .A3(KEYINPUT25), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT25), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n409), .A2(new_n411), .B1(new_n389), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n424), .B2(new_n419), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT77), .B1(new_n408), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n394), .A2(new_n399), .ZN(new_n428));
  INV_X1    g227(.A(new_n406), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n404), .B2(new_n397), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n381), .B(new_n383), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n421), .A2(new_n425), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n370), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n431), .A2(new_n433), .A3(new_n368), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n367), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(new_n434), .A3(new_n368), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n369), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n366), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(new_n441), .A3(new_n445), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT30), .A3(new_n448), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n345), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n303), .B2(new_n304), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT85), .B1(new_n456), .B2(new_n367), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n278), .A2(new_n304), .A3(new_n280), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n366), .ZN(new_n462));
  INV_X1    g261(.A(G228gat), .ZN(new_n463));
  INV_X1    g262(.A(G233gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n459), .B1(new_n354), .B2(new_n365), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n304), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n271), .A2(new_n467), .A3(new_n281), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n457), .A2(new_n462), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G22gat), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n367), .B1(new_n458), .B2(new_n459), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n360), .A2(new_n359), .A3(new_n363), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n459), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n303), .B1(new_n304), .B2(new_n474), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n471), .A2(new_n475), .B1(new_n463), .B2(new_n464), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n469), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n470), .B1(new_n469), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n455), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n468), .B(new_n465), .C1(new_n471), .C2(new_n461), .ZN(new_n480));
  INV_X1    g279(.A(new_n462), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G22gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n469), .A2(new_n470), .A3(new_n476), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT31), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G50gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n455), .B(new_n488), .C1(new_n477), .C2(new_n478), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT72), .B1(new_n408), .B2(new_n426), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n431), .A2(new_n494), .A3(new_n433), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(new_n320), .ZN(new_n496));
  NAND2_X1  g295(.A1(G227gat), .A2(G233gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n439), .A2(KEYINPUT72), .A3(new_n302), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT33), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT73), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(KEYINPUT73), .A3(new_n501), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G43gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G71gat), .B(G99gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n500), .B2(KEYINPUT32), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n500), .B(KEYINPUT32), .C1(new_n501), .C2(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT75), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n498), .B1(new_n496), .B2(new_n499), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n497), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n514), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n514), .B(new_n517), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n492), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n345), .A2(KEYINPUT84), .A3(new_n451), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n454), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT88), .B1(new_n338), .B2(new_n344), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n328), .A2(new_n333), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n337), .A4(new_n336), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n530), .A3(new_n334), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n510), .A2(new_n521), .A3(new_n511), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n521), .B1(new_n510), .B2(new_n511), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n532), .A2(new_n492), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n451), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n526), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n341), .A2(new_n342), .B1(new_n313), .B2(new_n317), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n336), .B(new_n337), .C1(new_n540), .C2(new_n332), .ZN(new_n541));
  AOI221_X4 g340(.A(new_n453), .B1(new_n450), .B2(new_n449), .C1(new_n541), .C2(new_n334), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT84), .B1(new_n345), .B2(new_n451), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n492), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n451), .A2(new_n344), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n311), .B1(new_n306), .B2(new_n309), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n332), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n321), .A2(new_n311), .A3(new_n322), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT87), .A3(KEYINPUT39), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT87), .B1(new_n550), .B2(KEYINPUT39), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n546), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT40), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n492), .B1(new_n545), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT90), .B1(new_n442), .B2(KEYINPUT37), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n437), .A2(new_n559), .A3(new_n560), .A4(new_n441), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n442), .A2(KEYINPUT37), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n446), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n560), .B1(new_n437), .B2(new_n441), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT91), .B1(new_n566), .B2(new_n445), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT38), .ZN(new_n569));
  INV_X1    g368(.A(new_n448), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n445), .A2(KEYINPUT38), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n435), .A2(new_n436), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT89), .B1(new_n572), .B2(new_n366), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n438), .A2(new_n440), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n366), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n435), .A2(new_n367), .A3(new_n436), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n560), .B1(new_n576), .B2(KEYINPUT89), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n571), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n570), .B1(new_n578), .B2(new_n562), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n569), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n557), .B1(new_n580), .B2(new_n531), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT36), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n521), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n521), .B1(new_n512), .B2(KEYINPUT75), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n585), .B2(KEYINPUT36), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n544), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n243), .B1(new_n539), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n596), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n595), .B(new_n602), .Z(new_n603));
  AND2_X1   g402(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n605));
  OAI21_X1  g404(.A(G57gat), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT95), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(G57gat), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n607), .B(new_n609), .C1(G57gat), .C2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(G71gat), .ZN(new_n612));
  INV_X1    g411(.A(G78gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n611), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n614), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n610), .A2(G57gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n610), .A2(G57gat), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT9), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n620), .B(new_n623), .C1(new_n619), .C2(new_n615), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  MUX2_X1   g424(.A(new_n600), .B(new_n603), .S(new_n625), .Z(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n626), .A2(new_n631), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT100), .Z(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n638), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(KEYINPUT99), .A3(new_n638), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n625), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G127gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n208), .B1(new_n625), .B2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G155gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n600), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n224), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(G232gat), .A2(G233gat), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n600), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G190gat), .B(G218gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(KEYINPUT41), .ZN(new_n667));
  XNOR2_X1  g466(.A(G134gat), .B(G162gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n645), .A2(new_n659), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n588), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n345), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT101), .B(G1gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  NOR2_X1   g478(.A1(new_n676), .A2(new_n451), .ZN(new_n680));
  NAND2_X1  g479(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n203), .A2(new_n206), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n206), .B2(new_n680), .ZN(new_n684));
  MUX2_X1   g483(.A(new_n683), .B(new_n684), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g484(.A(G15gat), .B1(new_n676), .B2(new_n586), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n532), .A2(new_n533), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n686), .B1(new_n676), .B2(new_n689), .ZN(G1326gat));
  INV_X1    g489(.A(new_n492), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  XNOR2_X1  g493(.A(new_n659), .B(KEYINPUT102), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n242), .A3(new_n645), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI211_X1 g496(.A(KEYINPUT44), .B(new_n673), .C1(new_n539), .C2(new_n587), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT35), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n542), .A2(new_n543), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n523), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n587), .B1(new_n702), .B2(new_n537), .ZN(new_n703));
  INV_X1    g502(.A(new_n673), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n699), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n697), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n544), .A2(new_n581), .A3(new_n586), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n537), .B1(new_n525), .B2(KEYINPUT35), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT44), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n703), .A2(new_n699), .A3(new_n704), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n697), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n345), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n704), .A2(new_n658), .A3(new_n657), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n588), .A2(new_n645), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n345), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n213), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n717), .A2(new_n724), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n720), .A2(G36gat), .A3(new_n451), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI211_X1 g532(.A(KEYINPUT105), .B(new_n726), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  INV_X1    g533(.A(new_n716), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n209), .B1(new_n735), .B2(new_n535), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n696), .B1(new_n711), .B2(new_n712), .ZN(new_n739));
  INV_X1    g538(.A(new_n586), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n688), .A2(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT47), .B1(new_n720), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT107), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G43gat), .B1(new_n706), .B2(new_n586), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747));
  INV_X1    g546(.A(new_n744), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n721), .A2(new_n751), .A3(new_n742), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n720), .B2(new_n743), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n707), .A2(new_n740), .A3(new_n715), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(G43gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n756), .B2(KEYINPUT47), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n750), .B(KEYINPUT108), .C1(new_n756), .C2(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1330gat));
  NOR2_X1   g560(.A1(new_n691), .A2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n720), .B2(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(KEYINPUT109), .B2(new_n720), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G50gat), .B1(new_n706), .B2(new_n691), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n735), .A2(new_n492), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(G50gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g570(.A(new_n242), .B1(new_n539), .B2(new_n587), .ZN(new_n772));
  INV_X1    g571(.A(new_n644), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT99), .B1(new_n635), .B2(new_n638), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n773), .A2(new_n774), .B1(new_n635), .B2(new_n639), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(new_n659), .A3(new_n673), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n345), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT110), .B(G57gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1332gat));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n777), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n535), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT49), .B(G64gat), .Z(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(G1333gat));
  NOR2_X1   g585(.A1(new_n586), .A2(new_n612), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n782), .A2(KEYINPUT112), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n687), .A3(new_n776), .ZN(new_n793));
  AOI21_X1  g592(.A(G71gat), .B1(new_n793), .B2(KEYINPUT113), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(KEYINPUT113), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT50), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n492), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g601(.A1(new_n772), .A2(new_n719), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT114), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n719), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n775), .A2(new_n592), .A3(new_n722), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n645), .A2(new_n659), .A3(new_n242), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n713), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n722), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G85gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT115), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n818), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1336gat));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n821), .A3(new_n807), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n803), .A2(KEYINPUT116), .A3(new_n804), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n645), .A2(G92gat), .A3(new_n451), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n593), .B1(new_n813), .B2(new_n535), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n808), .A2(new_n824), .ZN(new_n828));
  XNOR2_X1  g627(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(G1337gat));
  NOR3_X1   g630(.A1(new_n645), .A2(G99gat), .A3(new_n688), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n808), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n740), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G99gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1338gat));
  NOR3_X1   g635(.A1(new_n645), .A2(G106gat), .A3(new_n691), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n822), .A2(new_n823), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(G106gat), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n813), .B2(new_n492), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT53), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n808), .A2(new_n837), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(G1339gat));
  NOR2_X1   g643(.A1(new_n674), .A2(new_n242), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT118), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n674), .B2(new_n242), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n630), .A2(new_n631), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n633), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n638), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n632), .B2(KEYINPUT54), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n643), .A2(new_n644), .B1(new_n855), .B2(KEYINPUT55), .ZN(new_n856));
  INV_X1    g655(.A(new_n855), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n242), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n225), .A2(new_n226), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n230), .A2(new_n231), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n237), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n241), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n775), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n704), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n856), .A2(new_n859), .A3(new_n704), .A4(new_n865), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n695), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n722), .A3(new_n451), .A4(new_n534), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n285), .A3(new_n243), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n345), .B1(new_n849), .B2(new_n870), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n523), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n451), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n242), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(new_n285), .ZN(G1340gat));
  NOR3_X1   g677(.A1(new_n872), .A2(new_n283), .A3(new_n645), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n775), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n283), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n876), .A2(new_n290), .A3(new_n659), .ZN(new_n882));
  OAI21_X1  g681(.A(G127gat), .B1(new_n872), .B2(new_n695), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1342gat));
  NOR2_X1   g683(.A1(new_n673), .A2(new_n535), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n875), .A2(new_n293), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n872), .B2(new_n673), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n887), .B(new_n888), .C1(new_n890), .C2(new_n891), .ZN(G1343gat));
  NOR2_X1   g691(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n857), .A2(KEYINPUT122), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n858), .B1(new_n855), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n856), .B(new_n242), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n775), .A2(new_n899), .A3(new_n865), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT121), .B1(new_n645), .B2(new_n864), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n673), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n659), .B1(new_n903), .B2(new_n868), .ZN(new_n904));
  INV_X1    g703(.A(new_n849), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n492), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n586), .A2(new_n722), .A3(new_n451), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT120), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n691), .B1(new_n849), .B2(new_n870), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n907), .A2(new_n242), .A3(new_n909), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G141gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n740), .A2(new_n691), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n243), .A2(G141gat), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n874), .A2(new_n451), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n894), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n893), .B(new_n919), .C1(new_n913), .C2(G141gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(G1344gat));
  AND3_X1   g722(.A1(new_n874), .A2(new_n451), .A3(new_n915), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n775), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n265), .A3(new_n266), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n910), .A2(new_n911), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n911), .B(new_n492), .C1(new_n904), .C2(new_n845), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n909), .A2(new_n775), .ZN(new_n931));
  OAI211_X1 g730(.A(KEYINPUT59), .B(G148gat), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n907), .A2(new_n909), .A3(new_n912), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n645), .A2(KEYINPUT59), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n927), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(G155gat), .B1(new_n933), .B2(new_n695), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n248), .A3(new_n659), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n933), .B2(new_n673), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n874), .A2(new_n249), .A3(new_n885), .A4(new_n915), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n722), .A2(new_n451), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n849), .B2(new_n870), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n523), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(G169gat), .B1(new_n946), .B2(new_n242), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n944), .A2(new_n534), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n243), .A2(new_n372), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(G1348gat));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n373), .A3(new_n775), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n948), .A2(new_n775), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n373), .ZN(G1349gat));
  INV_X1    g752(.A(new_n414), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n659), .B(KEYINPUT102), .Z(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n659), .A2(new_n398), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT124), .B1(new_n945), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g759(.A(new_n423), .B1(new_n948), .B2(new_n704), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n673), .A2(new_n413), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT125), .B1(new_n945), .B2(new_n968), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n945), .A2(KEYINPUT125), .A3(new_n968), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n962), .A2(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n965), .A2(new_n971), .ZN(G1351gat));
  XOR2_X1   g771(.A(KEYINPUT127), .B(G197gat), .Z(new_n973));
  NOR2_X1   g772(.A1(new_n740), .A2(new_n943), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n928), .A2(new_n929), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n973), .B1(new_n975), .B2(new_n243), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n910), .A2(new_n974), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n243), .A2(new_n973), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR3_X1   g778(.A1(new_n977), .A2(G204gat), .A3(new_n645), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n975), .B2(new_n645), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1353gat));
  INV_X1    g782(.A(new_n977), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n361), .A3(new_n659), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n928), .A2(new_n659), .A3(new_n929), .A4(new_n974), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n975), .B2(new_n673), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n984), .A2(new_n362), .A3(new_n704), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


