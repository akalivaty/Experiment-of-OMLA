//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT78), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(G134), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(G137), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n198), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n199), .A2(new_n200), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT11), .B1(new_n205), .B2(new_n202), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT65), .A2(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT65), .A2(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n202), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n198), .ZN(new_n212));
  INV_X1    g026(.A(new_n203), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G134), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G137), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n208), .B(new_n212), .C1(new_n215), .C2(new_n198), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(KEYINPUT3), .A3(G104), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n218), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(G107), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n219), .A2(KEYINPUT3), .A3(G104), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(new_n219), .B2(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(KEYINPUT0), .B2(G128), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT0), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT64), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n234), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n239), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n231), .A2(new_n218), .A3(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n233), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT66), .B(G128), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(G143), .B2(new_n240), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n244), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n236), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n219), .A2(G104), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n226), .B1(new_n228), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n225), .B2(new_n226), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n262), .A3(KEYINPUT10), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n226), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n264));
  INV_X1    g078(.A(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT1), .B1(new_n242), .B2(G146), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n267), .A2(G128), .B1(new_n241), .B2(new_n243), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n257), .A2(new_n241), .A3(new_n243), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT79), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n246), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n258), .B1(new_n272), .B2(new_n236), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT79), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n262), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT10), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n252), .B(new_n263), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT10), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n262), .A2(new_n273), .A3(new_n274), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n262), .B2(new_n273), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n217), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(new_n217), .C1(new_n278), .C2(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n271), .A2(new_n275), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n277), .A3(new_n279), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n252), .A2(new_n263), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n217), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n289), .A2(new_n291), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n292), .B1(KEYINPUT80), .B2(new_n282), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(KEYINPUT81), .A3(new_n294), .A4(new_n291), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n197), .B1(new_n288), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n256), .A2(new_n258), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n266), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n290), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n217), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT83), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT12), .ZN(new_n308));
  INV_X1    g122(.A(new_n304), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(new_n294), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n304), .A2(new_n311), .A3(new_n217), .A4(new_n305), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n300), .A2(new_n197), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n191), .B(new_n189), .C1(new_n301), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT86), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n300), .A2(new_n197), .A3(new_n313), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n285), .A2(new_n287), .B1(new_n297), .B2(new_n299), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(new_n197), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n191), .A4(new_n189), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n300), .A2(new_n313), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n197), .B1(new_n323), .B2(KEYINPUT84), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n300), .A2(new_n325), .A3(new_n313), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n196), .B1(new_n297), .B2(new_n299), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n324), .A2(new_n326), .B1(new_n288), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G469), .B1(new_n328), .B2(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n190), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT32), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n211), .B1(G134), .B2(new_n202), .ZN(new_n333));
  AOI22_X1  g147(.A1(G131), .A2(new_n333), .B1(new_n256), .B2(new_n258), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n334), .A2(new_n216), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n249), .B1(new_n207), .B2(new_n216), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n217), .A2(new_n250), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n216), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(KEYINPUT30), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G119), .ZN(new_n341));
  OR2_X1    g155(.A1(KEYINPUT67), .A2(G116), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT67), .A2(G116), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G116), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G119), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT68), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n343), .ZN(new_n348));
  NOR2_X1   g162(.A1(KEYINPUT67), .A2(G116), .ZN(new_n349));
  OAI21_X1  g163(.A(G119), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n351));
  INV_X1    g165(.A(new_n346), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT2), .B(G113), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n347), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n352), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n356), .A2(new_n354), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n337), .A2(new_n340), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n360));
  INV_X1    g174(.A(new_n358), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n338), .A2(new_n361), .A3(new_n339), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n363));
  NOR2_X1   g177(.A1(G237), .A2(G953), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G210), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n363), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G101), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n360), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT71), .A2(KEYINPUT31), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT71), .A2(KEYINPUT31), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(new_n360), .A3(new_n368), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n335), .A2(new_n336), .A3(new_n358), .ZN(new_n376));
  INV_X1    g190(.A(new_n368), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT70), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n337), .A2(new_n340), .A3(new_n358), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n373), .A3(new_n374), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n371), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n358), .B1(new_n335), .B2(new_n336), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(new_n362), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT72), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n384), .A2(new_n385), .B1(new_n382), .B2(new_n362), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n362), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT28), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT72), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n375), .A2(new_n381), .B1(new_n390), .B2(new_n377), .ZN(new_n391));
  NOR2_X1   g205(.A1(G472), .A2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n331), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(new_n385), .A3(KEYINPUT28), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n362), .A2(new_n382), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n384), .A2(new_n385), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n377), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n380), .A2(new_n371), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n380), .A2(new_n371), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT32), .A3(new_n392), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n386), .A2(new_n389), .A3(new_n368), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n362), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n405), .B2(new_n377), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n388), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n388), .A2(KEYINPUT73), .A3(new_n396), .A4(new_n408), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n189), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G472), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n394), .A2(new_n403), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G125), .B(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n417));
  INV_X1    g231(.A(G125), .ZN(new_n418));
  OR3_X1    g232(.A1(new_n418), .A2(KEYINPUT16), .A3(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n240), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(G146), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT74), .B1(new_n341), .B2(G128), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n246), .A3(G119), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n246), .A2(G119), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n425), .B(new_n427), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n428), .B1(new_n253), .B2(G119), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT24), .B(G110), .Z(new_n433));
  AOI22_X1  g247(.A1(new_n431), .A2(G110), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT75), .Z(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT76), .B(G110), .ZN(new_n437));
  OAI22_X1  g251(.A1(new_n431), .A2(new_n437), .B1(new_n432), .B2(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n416), .A2(new_n240), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n422), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT77), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT22), .B(G137), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n442), .A3(new_n446), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n189), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT25), .A4(new_n189), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G217), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G234), .B2(new_n189), .ZN(new_n456));
  INV_X1    g270(.A(new_n448), .ZN(new_n457));
  INV_X1    g271(.A(new_n449), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n456), .A2(G902), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n454), .A2(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n415), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n246), .A2(G143), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n253), .B2(G143), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT13), .ZN(new_n465));
  INV_X1    g279(.A(new_n463), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(G134), .C1(KEYINPUT13), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n214), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n345), .A2(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT98), .ZN(new_n470));
  OAI21_X1  g284(.A(G122), .B1(new_n348), .B2(new_n349), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n219), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n472), .A2(new_n219), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n467), .B(new_n468), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT99), .B1(new_n471), .B2(KEYINPUT14), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(KEYINPUT14), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n470), .A3(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n471), .A2(KEYINPUT99), .A3(KEYINPUT14), .ZN(new_n480));
  OAI21_X1  g294(.A(G107), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n464), .B(new_n214), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n188), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n485), .A2(new_n455), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n476), .A2(new_n483), .A3(new_n486), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n490), .B1(KEYINPUT15), .B2(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n222), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT95), .Z(new_n499));
  AND3_X1   g313(.A1(new_n364), .A2(G143), .A3(G214), .ZN(new_n500));
  AOI21_X1  g314(.A(G143), .B1(new_n364), .B2(G214), .ZN(new_n501));
  OAI21_X1  g315(.A(G131), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n503));
  OR3_X1    g317(.A1(new_n502), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT93), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n416), .A2(new_n240), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  NAND2_X1  g321(.A1(KEYINPUT18), .A2(G131), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n439), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n208), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n502), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n502), .A2(new_n512), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n422), .A4(new_n421), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n499), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n498), .B1(new_n515), .B2(new_n510), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n189), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n518), .A2(KEYINPUT97), .ZN(new_n519));
  OAI21_X1  g333(.A(G475), .B1(new_n518), .B2(KEYINPUT97), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n496), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(G234), .A2(G237), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n523), .A2(G902), .A3(G953), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT21), .B(G898), .Z(new_n526));
  OR2_X1    g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n523), .A2(G952), .A3(new_n192), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G475), .A2(G902), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n511), .A2(new_n502), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT94), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n511), .A2(new_n535), .A3(new_n502), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n416), .B(KEYINPUT19), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n240), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n534), .A2(new_n422), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n498), .B1(new_n539), .B2(new_n510), .ZN(new_n540));
  OAI221_X1 g354(.A(new_n531), .B1(new_n532), .B2(KEYINPUT20), .C1(new_n540), .C2(new_n516), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n531), .B1(new_n540), .B2(new_n516), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n540), .A2(new_n516), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(KEYINPUT96), .ZN(new_n545));
  AND4_X1   g359(.A1(new_n522), .A2(new_n530), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G214), .B1(G237), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n249), .A2(G125), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n249), .A2(new_n554), .A3(G125), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n249), .B2(G125), .ZN(new_n557));
  AOI211_X1 g371(.A(KEYINPUT89), .B(new_n418), .C1(new_n239), .C2(new_n248), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT90), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n192), .A2(G224), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n302), .A2(new_n563), .A3(new_n418), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT91), .B1(new_n259), .B2(G125), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n560), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT5), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n347), .B2(new_n353), .ZN(new_n571));
  OAI21_X1  g385(.A(G113), .B1(new_n352), .B2(KEYINPUT5), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n357), .B(new_n262), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT87), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n344), .A2(KEYINPUT68), .A3(new_n346), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT5), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n572), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n357), .A4(new_n262), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G122), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n233), .A2(new_n251), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n358), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n575), .A2(new_n581), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT88), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n573), .A2(new_n574), .B1(new_n583), .B2(new_n358), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(new_n581), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT6), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n575), .A2(new_n581), .A3(new_n584), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT6), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n569), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n566), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n557), .A2(new_n558), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n564), .A2(KEYINPUT92), .A3(new_n565), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n560), .A2(KEYINPUT7), .A3(new_n562), .A4(new_n566), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n580), .A2(new_n357), .A3(new_n266), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n582), .B(KEYINPUT8), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n579), .B1(new_n356), .B2(new_n570), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(new_n357), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n606), .B(new_n607), .C1(new_n266), .C2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n604), .A2(new_n605), .A3(new_n585), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n189), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n550), .B1(new_n597), .B2(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n567), .A2(new_n568), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n595), .B1(new_n594), .B2(new_n585), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n591), .A2(KEYINPUT6), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n611), .A2(new_n189), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n549), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n548), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n330), .A2(new_n462), .A3(new_n546), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n322), .A2(new_n329), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n619), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n547), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT101), .B(new_n548), .C1(new_n613), .C2(new_n619), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n190), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n391), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(G472), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(KEYINPUT100), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(KEYINPUT100), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n391), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n461), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n488), .A2(new_n489), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n488), .A2(KEYINPUT33), .A3(new_n489), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(G478), .A3(new_n189), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n491), .A2(new_n492), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n545), .B(new_n541), .C1(new_n519), .C2(new_n520), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n527), .B2(new_n529), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(new_n496), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n530), .B(KEYINPUT103), .Z(new_n654));
  NAND3_X1  g468(.A1(new_n542), .A2(KEYINPUT102), .A3(new_n543), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n656));
  OAI21_X1  g470(.A(new_n655), .B1(new_n542), .B2(new_n656), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n653), .A2(new_n521), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n639), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n447), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n443), .B(new_n662), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n454), .A2(new_n456), .B1(new_n460), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n636), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n330), .A3(new_n546), .A4(new_n620), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n454), .A2(new_n456), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n663), .A2(new_n460), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n415), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n529), .B1(new_n525), .B2(G900), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n653), .A2(new_n521), .A3(new_n657), .A4(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n630), .A2(new_n669), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n330), .A2(new_n676), .A3(new_n673), .A4(new_n628), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  INV_X1    g495(.A(new_n330), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n674), .B(KEYINPUT39), .Z(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n378), .A2(new_n374), .A3(new_n379), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n387), .A2(new_n377), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(KEYINPUT105), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n189), .B1(new_n689), .B2(KEYINPUT105), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n394), .A2(new_n403), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n625), .B(KEYINPUT38), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n647), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n653), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n547), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n664), .A2(new_n686), .A3(new_n693), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n684), .B2(new_n685), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  NOR2_X1   g516(.A1(new_n648), .A2(new_n675), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n330), .A2(new_n628), .A3(new_n673), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT107), .B(G146), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G48));
  AOI21_X1  g520(.A(new_n191), .B1(new_n319), .B2(new_n189), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n190), .B(new_n707), .C1(new_n316), .C2(new_n321), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n462), .A3(new_n649), .A4(new_n628), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n462), .A3(new_n628), .A4(new_n658), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AOI21_X1  g529(.A(new_n707), .B1(new_n316), .B2(new_n321), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n628), .A2(new_n629), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n546), .A2(new_n415), .A3(new_n672), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n708), .A2(new_n628), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n673), .A2(new_n546), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  INV_X1    g539(.A(new_n654), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n496), .A2(new_n647), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n391), .B2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n375), .A2(new_n381), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n388), .A2(new_n396), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n377), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n393), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n461), .A2(new_n727), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n708), .A2(new_n734), .A3(new_n628), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  INV_X1    g550(.A(new_n728), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(new_n664), .A3(new_n732), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n703), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n721), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n418), .ZN(G27));
  NAND3_X1  g555(.A1(new_n613), .A2(new_n619), .A3(new_n547), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n330), .A2(new_n462), .A3(new_n703), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n190), .B(new_n742), .C1(new_n322), .C2(new_n329), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n462), .A4(new_n703), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND3_X1  g568(.A1(new_n747), .A2(new_n462), .A3(new_n676), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NAND2_X1  g570(.A1(new_n324), .A2(new_n326), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n288), .A2(new_n327), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n191), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n328), .A2(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(KEYINPUT111), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n761), .A2(new_n762), .B1(G469), .B2(G902), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(KEYINPUT46), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(new_n770), .A3(new_n322), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n629), .ZN(new_n773));
  INV_X1    g587(.A(new_n646), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(KEYINPUT43), .A3(new_n647), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n696), .A2(KEYINPUT112), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n696), .A2(KEYINPUT112), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n646), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n778), .B2(KEYINPUT43), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n664), .B1(new_n633), .B2(new_n635), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT44), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(KEYINPUT44), .A3(new_n780), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n742), .B(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n773), .A2(new_n683), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT114), .B(G137), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G39));
  NOR2_X1   g601(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n772), .B2(new_n629), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n637), .A2(new_n703), .A3(new_n743), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n415), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  INV_X1    g609(.A(G952), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n192), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n528), .A2(new_n716), .A3(new_n629), .A4(new_n743), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n637), .A2(new_n693), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n647), .A3(new_n646), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n637), .A2(new_n737), .A3(new_n732), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n779), .A2(new_n528), .A3(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n796), .B(G953), .C1(new_n803), .C2(new_n717), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n779), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT118), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n462), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n801), .B(new_n804), .C1(new_n807), .C2(KEYINPUT48), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(KEYINPUT48), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n800), .A2(new_n696), .A3(new_n774), .ZN(new_n811));
  NOR2_X1   g625(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n694), .A2(new_n547), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n803), .A2(new_n708), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n815));
  NAND4_X1  g629(.A1(new_n813), .A2(new_n779), .A3(new_n528), .A4(new_n802), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n716), .A2(new_n629), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n811), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n806), .A2(new_n738), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT51), .ZN(new_n821));
  INV_X1    g635(.A(new_n716), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n788), .A2(new_n790), .B1(new_n629), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n803), .A2(new_n783), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n810), .B1(new_n826), .B2(KEYINPUT120), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(KEYINPUT120), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n822), .A2(new_n629), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n788), .A2(new_n790), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(KEYINPUT116), .ZN(new_n833));
  OR3_X1    g647(.A1(new_n788), .A2(KEYINPUT116), .A3(new_n790), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n819), .A2(new_n820), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT119), .Z(new_n837));
  OAI21_X1  g651(.A(new_n830), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n709), .A2(new_n735), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n720), .B2(new_n723), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n496), .A2(new_n521), .A3(new_n657), .A4(new_n675), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n415), .A2(new_n672), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n739), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n747), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n696), .A2(new_n496), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n654), .B1(new_n846), .B2(new_n648), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n638), .A2(new_n330), .A3(new_n620), .A4(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n666), .A2(new_n848), .A3(new_n621), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n714), .A2(new_n841), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n740), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n693), .A2(new_n664), .A3(new_n674), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n330), .A2(new_n852), .A3(new_n628), .A4(new_n697), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n704), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n680), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  INV_X1    g670(.A(new_n755), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n750), .B2(new_n752), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n740), .B1(new_n677), .B2(new_n679), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n854), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n850), .A2(new_n856), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT53), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n704), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(KEYINPUT115), .B(new_n740), .C1(new_n677), .C2(new_n679), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n860), .B1(new_n867), .B2(new_n853), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n850), .A2(new_n869), .A3(new_n858), .A4(new_n861), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n863), .B(KEYINPUT54), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n841), .A2(new_n714), .A3(new_n849), .ZN(new_n872));
  AND4_X1   g686(.A1(KEYINPUT53), .A2(new_n749), .A3(new_n755), .A4(new_n845), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n872), .A2(new_n861), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n853), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n865), .A2(new_n875), .A3(new_n866), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(new_n860), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n862), .A2(new_n869), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n797), .B1(new_n839), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n694), .A2(new_n778), .A3(new_n190), .A4(new_n548), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(new_n884), .A3(new_n799), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n886), .ZN(G75));
  AOI21_X1  g701(.A(new_n189), .B1(new_n877), .B2(new_n878), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(G210), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n592), .A2(new_n569), .A3(new_n596), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n617), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n889), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n889), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n192), .A2(G952), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G51));
  AND2_X1   g713(.A1(new_n862), .A2(new_n869), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n872), .A2(new_n873), .A3(new_n861), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n859), .A2(new_n864), .ZN(new_n902));
  INV_X1    g716(.A(new_n866), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n704), .A4(new_n853), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n901), .B1(new_n904), .B2(KEYINPUT52), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n880), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n764), .B(KEYINPUT57), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n319), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n888), .A2(new_n762), .A3(new_n761), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n898), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND2_X1  g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT122), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n888), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n544), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n544), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n898), .ZN(G60));
  XNOR2_X1  g732(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n492), .A2(new_n189), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n881), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n642), .A2(new_n643), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n871), .B2(new_n880), .ZN(new_n927));
  INV_X1    g741(.A(new_n925), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT124), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n921), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n898), .B1(new_n907), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n926), .A2(new_n929), .A3(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(new_n877), .A2(new_n878), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n459), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n898), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n933), .A2(new_n663), .A3(new_n936), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n940), .A4(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(G66));
  AOI21_X1  g760(.A(new_n192), .B1(new_n526), .B2(G224), .ZN(new_n947));
  INV_X1    g761(.A(new_n872), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n192), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n592), .B(new_n596), .C1(G898), .C2(new_n192), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n949), .B(new_n950), .Z(G69));
  NAND2_X1  g765(.A1(new_n337), .A2(new_n340), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n537), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(G900), .B(G953), .C1(new_n954), .C2(G227), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(G227), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n867), .A2(new_n701), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n867), .A2(KEYINPUT62), .A3(new_n701), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n785), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n742), .B1(new_n648), .B2(new_n846), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n684), .A2(new_n462), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n794), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n953), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n773), .A2(new_n683), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n462), .A2(new_n628), .A3(new_n697), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n858), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n785), .B1(new_n791), .B2(new_n793), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(new_n867), .ZN(new_n972));
  AOI21_X1  g786(.A(G953), .B1(new_n972), .B2(new_n954), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n956), .B1(new_n966), .B2(new_n973), .ZN(G72));
  AOI21_X1  g788(.A(new_n377), .B1(new_n379), .B2(new_n362), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n948), .B(new_n965), .C1(new_n959), .C2(new_n960), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n975), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n970), .A2(new_n971), .A3(new_n872), .A4(new_n867), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT125), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n984), .A3(new_n978), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n405), .A2(new_n368), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n868), .A2(new_n870), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(KEYINPUT53), .B2(new_n862), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n405), .A2(new_n377), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n687), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n978), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n898), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n980), .A2(new_n987), .A3(new_n996), .ZN(G57));
endmodule


