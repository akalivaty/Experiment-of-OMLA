//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI211_X1 g050(.A(KEYINPUT69), .B(new_n466), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n465), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n480), .B(new_n482), .C1(G124), .C2(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n469), .B2(new_n470), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(KEYINPUT70), .B(new_n487), .C1(new_n469), .C2(new_n470), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n466), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n496), .A2(new_n498), .A3(new_n499), .A4(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n483), .A2(new_n502), .A3(KEYINPUT4), .A4(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n469), .B2(new_n470), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n492), .A2(new_n501), .A3(new_n505), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n511), .A2(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n511), .B2(new_n512), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(new_n518), .B2(G50), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n515), .A2(new_n516), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n527), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(new_n521), .A2(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n520), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n521), .A2(new_n527), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n528), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n538), .A2(new_n539), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n520), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n541), .A2(new_n551), .B1(new_n528), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT75), .Z(G188));
  AOI22_X1  g136(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n520), .B1(new_n563), .B2(new_n541), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n528), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n518), .A2(G53), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n564), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  NOR2_X1   g147(.A1(new_n522), .A2(new_n520), .ZN(new_n573));
  INV_X1    g148(.A(G88), .ZN(new_n574));
  INV_X1    g149(.A(G50), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n541), .A2(new_n574), .B1(new_n528), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT77), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n519), .B(new_n578), .C1(new_n520), .C2(new_n522), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(G303));
  NAND2_X1  g155(.A1(new_n517), .A2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n518), .A2(G49), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n517), .A2(G86), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n515), .B2(new_n516), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n518), .A2(G48), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n520), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n541), .A2(new_n594), .B1(new_n528), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n518), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n521), .A2(new_n527), .A3(G92), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n605));
  OAI221_X1 g180(.A(new_n601), .B1(new_n520), .B2(new_n602), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT79), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n600), .B1(new_n610), .B2(new_n611), .ZN(G284));
  XNOR2_X1  g187(.A(G284), .B(KEYINPUT80), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n570), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n570), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n607), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n483), .A2(new_n467), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT81), .B(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n465), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n466), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n632), .C2(new_n484), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT82), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n642), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(new_n650), .A3(G14), .ZN(G401));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT83), .ZN(new_n653));
  NOR2_X1   g228(.A1(G2072), .A2(G2078), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n442), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n655), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n655), .B(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n657), .C1(new_n653), .C2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n653), .A2(new_n661), .A3(new_n656), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n669), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n669), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G24), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n597), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n485), .A2(G119), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n465), .A2(G131), .ZN(new_n694));
  OR2_X1    g269(.A1(G95), .A2(G2105), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n695), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(new_n691), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT87), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  AOI21_X1  g276(.A(new_n690), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n687), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n687), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n687), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n687), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G6), .A2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G305), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n719), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n702), .B1(new_n701), .B2(new_n700), .C1(new_n720), .C2(KEYINPUT34), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(KEYINPUT34), .B2(new_n720), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT36), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n687), .A2(G5), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G171), .B2(new_n687), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G1961), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n691), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(new_n727), .ZN(new_n730));
  INV_X1    g305(.A(G160), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n691), .A2(G32), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  INV_X1    g312(.A(G129), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n737), .C1(new_n738), .C2(new_n484), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT97), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n691), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT98), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n726), .B1(G2084), .B2(new_n733), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT101), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n691), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT89), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n485), .A2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n465), .A2(G140), .ZN(new_n750));
  OR2_X1    g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n691), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT90), .B(G2067), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n687), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n554), .B2(new_n687), .ZN(new_n759));
  INV_X1    g334(.A(G1341), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n687), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n607), .B2(new_n687), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n757), .B(new_n761), .C1(new_n763), .C2(G1348), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G1348), .B2(new_n763), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT91), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n691), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n483), .A2(G127), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n466), .B1(new_n770), .B2(KEYINPUT92), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT92), .B2(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n773));
  NAND2_X1  g348(.A1(G103), .A2(G2104), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G2105), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n465), .A2(G139), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n767), .B1(new_n778), .B2(new_n691), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT93), .B(G2072), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n691), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n691), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT29), .B(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT31), .B(G11), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT100), .B(G28), .Z(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT30), .B2(new_n787), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n789), .C1(new_n633), .C2(new_n691), .ZN(new_n790));
  NOR2_X1   g365(.A1(G168), .A2(new_n687), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n687), .B2(G21), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT99), .B(G1966), .Z(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n781), .A2(new_n785), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n725), .A2(G1961), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n691), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n691), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n687), .A2(G20), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT23), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n570), .B2(new_n687), .ZN(new_n804));
  INV_X1    g379(.A(G1956), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n796), .A2(new_n797), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n733), .A2(G2084), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT96), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n807), .B(new_n809), .C1(new_n743), .C2(new_n742), .ZN(new_n810));
  AND4_X1   g385(.A1(new_n723), .A2(new_n745), .A3(new_n766), .A4(new_n810), .ZN(G311));
  NAND4_X1  g386(.A1(new_n723), .A2(new_n745), .A3(new_n766), .A4(new_n810), .ZN(G150));
  NAND2_X1  g387(.A1(new_n607), .A2(G559), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  INV_X1    g389(.A(G55), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n541), .A2(new_n814), .B1(new_n528), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n521), .A2(G67), .ZN(new_n817));
  AND2_X1   g392(.A1(G80), .A2(G543), .ZN(new_n818));
  OAI21_X1  g393(.A(G651), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n819), .B2(KEYINPUT102), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT102), .B2(new_n819), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n550), .A2(new_n553), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT103), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n554), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n821), .A2(new_n823), .A3(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n813), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  AOI21_X1  g409(.A(G860), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n821), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G145));
  INV_X1    g415(.A(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n466), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n484), .A2(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G142), .B2(new_n465), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n624), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n698), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n778), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G164), .ZN(new_n851));
  INV_X1    g426(.A(new_n740), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n754), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n754), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n848), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(G162), .B(new_n633), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G160), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n853), .A2(new_n754), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n854), .A3(new_n847), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n848), .A2(KEYINPUT107), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n855), .B2(new_n856), .ZN(new_n865));
  INV_X1    g440(.A(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n855), .A2(new_n856), .A3(new_n864), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n862), .B(new_n863), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g445(.A(new_n619), .B(new_n830), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n606), .A2(new_n570), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT108), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n606), .A2(new_n570), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n606), .A2(new_n875), .A3(new_n570), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n877), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n871), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n597), .B(new_n716), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n704), .B(new_n523), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n883), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n821), .A2(new_n609), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n895));
  XNOR2_X1  g470(.A(G168), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G301), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n828), .A3(new_n829), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n896), .A2(G301), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(G301), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n830), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n897), .A2(KEYINPUT110), .A3(new_n828), .A4(new_n829), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n879), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n901), .A3(new_n877), .ZN(new_n906));
  INV_X1    g481(.A(new_n887), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(G37), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT111), .B1(new_n910), .B2(G37), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT43), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n898), .A2(new_n901), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n879), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n881), .B1(new_n903), .B2(new_n904), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n887), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(new_n863), .A3(new_n908), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT112), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n923), .A3(new_n863), .A4(new_n908), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n916), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n915), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n916), .B1(new_n913), .B2(new_n914), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT127), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT113), .B(G1384), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT45), .B1(new_n509), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G40), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n475), .A2(new_n936), .A3(new_n476), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n753), .B(G2067), .Z(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n852), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n740), .A2(G1996), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n697), .B(new_n701), .Z(new_n944));
  OR2_X1    g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n597), .B(G1986), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT70), .B1(new_n483), .B2(new_n487), .ZN(new_n951));
  INV_X1    g526(.A(new_n491), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(KEYINPUT114), .B(new_n949), .C1(new_n950), .C2(new_n953), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT45), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n937), .B1(new_n959), .B2(new_n954), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n793), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n471), .A2(new_n472), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT69), .B1(new_n964), .B2(new_n466), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n473), .A2(new_n474), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n965), .A2(new_n966), .A3(G40), .A4(new_n468), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(KEYINPUT50), .B2(new_n954), .ZN(new_n968));
  INV_X1    g543(.A(G2084), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(G168), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G8), .ZN(new_n972));
  AOI21_X1  g547(.A(G168), .B1(new_n961), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT51), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n975), .A3(G8), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT62), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n577), .A2(new_n579), .A3(KEYINPUT55), .A4(G8), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n577), .A2(G8), .A3(new_n579), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n962), .B1(new_n956), .B2(new_n957), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n937), .B1(KEYINPUT50), .B2(new_n954), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT118), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n957), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT114), .B1(new_n509), .B2(new_n949), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT50), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n954), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n967), .B1(new_n995), .B2(new_n962), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G2090), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n954), .A2(new_n959), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n937), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n713), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n988), .B1(new_n1005), .B2(G8), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1001), .A2(new_n800), .A3(new_n937), .A4(new_n1002), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1961), .B1(new_n963), .B2(new_n968), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n958), .A2(new_n960), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(KEYINPUT53), .A3(new_n800), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G171), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n963), .A2(new_n968), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1004), .B1(new_n1016), .B2(G2090), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(new_n988), .A3(G8), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n956), .A2(new_n937), .A3(new_n957), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n704), .A2(G1976), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n589), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G305), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n517), .A2(G86), .B1(new_n518), .B2(G48), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n589), .C1(new_n1026), .C2(new_n1025), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT49), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1030), .A3(KEYINPUT49), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1028), .A2(new_n1030), .A3(KEYINPUT117), .A4(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1019), .A2(G8), .A3(new_n1021), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1020), .A2(new_n1036), .B1(new_n1037), .B2(KEYINPUT52), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1018), .A2(new_n1024), .A3(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1006), .A2(new_n1015), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n978), .A2(new_n980), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n961), .A2(new_n970), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(G8), .A3(G168), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1038), .A2(new_n1024), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1017), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n988), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1045), .A2(new_n1018), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1006), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(KEYINPUT63), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1020), .A2(new_n1036), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n1022), .A3(new_n704), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(G1981), .B2(G305), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1018), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1055), .A2(new_n1020), .B1(new_n1046), .B2(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1041), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n567), .A2(new_n569), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n567), .B2(new_n569), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n564), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT120), .B1(new_n1063), .B2(KEYINPUT57), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(new_n564), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1060), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n570), .A2(KEYINPUT57), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1064), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n805), .B1(new_n989), .B2(new_n990), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT56), .B(G2072), .Z(new_n1073));
  OR2_X1    g648(.A1(new_n1003), .A2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1019), .A2(G2067), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1016), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1075), .A2(new_n608), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1071), .A2(KEYINPUT121), .ZN(new_n1080));
  AOI22_X1  g655(.A1(KEYINPUT121), .A2(new_n1071), .B1(new_n1074), .B2(new_n1072), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1071), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1075), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1075), .B2(new_n1083), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(new_n760), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1019), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1001), .A2(new_n940), .A3(new_n937), .A4(new_n1002), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n822), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1085), .A2(new_n1087), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1078), .A2(KEYINPUT60), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n608), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n607), .B1(new_n1078), .B2(KEYINPUT60), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1082), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  AOI21_X1  g678(.A(G301), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1104));
  AND4_X1   g679(.A1(KEYINPUT53), .A2(new_n468), .A3(G40), .A4(new_n800), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n1106));
  OAI21_X1  g681(.A(G2105), .B1(new_n964), .B2(KEYINPUT124), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1002), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n935), .ZN(new_n1109));
  NOR4_X1   g684(.A1(new_n1009), .A2(new_n1010), .A3(new_n1109), .A4(G171), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1103), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT125), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1006), .A2(new_n1039), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1011), .A2(G301), .A3(new_n1013), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1009), .A2(new_n1010), .A3(new_n1109), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1114), .B(KEYINPUT54), .C1(G301), .C2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1113), .A2(new_n977), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1102), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n948), .B1(new_n1058), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n938), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n945), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT126), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n938), .A2(G1986), .A3(G290), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT48), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n938), .B1(new_n939), .B2(new_n740), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n938), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT46), .B1(new_n938), .B2(G1996), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT47), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n698), .A2(new_n701), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n943), .A2(new_n1131), .B1(G2067), .B2(new_n753), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1120), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1125), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n932), .B1(new_n1119), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n948), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1102), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1041), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1134), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT127), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g717(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1144));
  OAI211_X1 g718(.A(new_n869), .B(new_n1144), .C1(new_n928), .C2(new_n929), .ZN(G225));
  INV_X1    g719(.A(G225), .ZN(G308));
endmodule


