//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n196), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n195), .B1(new_n200), .B2(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n199), .A2(new_n208), .B1(KEYINPUT0), .B2(G128), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n199), .A2(new_n208), .A3(G128), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n206), .A2(new_n209), .B1(new_n210), .B2(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G224), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n213), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT83), .A2(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT83), .A2(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT84), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT84), .B1(new_n222), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT85), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT85), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n236), .A3(KEYINPUT4), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n244), .B1(new_n247), .B2(new_n243), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(G101), .C1(new_n228), .C2(new_n229), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT83), .A2(G107), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT83), .A2(G107), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n226), .B1(new_n255), .B2(G104), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n234), .A2(new_n235), .B1(G101), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(G113), .B1(new_n239), .B2(KEYINPUT5), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n247), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n244), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G122), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(KEYINPUT89), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n252), .B2(new_n263), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT6), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n252), .A2(new_n263), .ZN(new_n270));
  INV_X1    g084(.A(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n217), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n215), .A2(KEYINPUT7), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n203), .A2(new_n212), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT90), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n256), .A2(G101), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n255), .A2(new_n219), .B1(new_n226), .B2(new_n225), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT85), .B1(new_n281), .B2(new_n231), .ZN(new_n282));
  INV_X1    g096(.A(new_n235), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n262), .A3(new_n261), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n242), .A2(new_n260), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n262), .B1(new_n286), .B2(new_n258), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n257), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n264), .B(KEYINPUT8), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n213), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n279), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n276), .B1(new_n292), .B2(new_n266), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n190), .B1(new_n275), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n273), .B1(new_n272), .B2(new_n265), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n268), .A2(KEYINPUT6), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n216), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n279), .A2(new_n290), .A3(new_n291), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n298), .B2(new_n265), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n189), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n188), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT91), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n237), .A2(new_n211), .A3(new_n251), .ZN(new_n306));
  AOI21_X1  g120(.A(G128), .B1(new_n199), .B2(new_n208), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n207), .A2(KEYINPUT1), .A3(G146), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT86), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n311), .B(new_n308), .C1(new_n194), .C2(G128), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n195), .A3(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n280), .C1(new_n282), .C2(new_n283), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n199), .B1(new_n191), .B2(new_n192), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n194), .B1(new_n318), .B2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n199), .A2(new_n208), .A3(G128), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n197), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT69), .B(new_n195), .C1(new_n200), .C2(new_n194), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n306), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT11), .A3(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n330), .A3(new_n334), .A4(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n336), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n306), .A2(new_n338), .A3(new_n316), .A4(new_n324), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G140), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT82), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n214), .A2(G227), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT12), .ZN(new_n348));
  INV_X1    g162(.A(new_n201), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n284), .A2(new_n349), .ZN(new_n350));
  AOI211_X1 g164(.A(new_n348), .B(new_n338), .C1(new_n350), .C2(new_n314), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n314), .B1(new_n201), .B2(new_n257), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT12), .B1(new_n352), .B2(new_n336), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n339), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT87), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n339), .C1(new_n351), .C2(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n345), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n347), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G469), .B1(new_n360), .B2(G902), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n339), .B(new_n345), .C1(new_n351), .C2(new_n353), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n314), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n201), .B1(new_n236), .B2(new_n280), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n336), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n348), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n352), .A2(KEYINPUT12), .A3(new_n336), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT88), .A3(new_n339), .A4(new_n345), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n345), .B1(new_n337), .B2(new_n339), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G469), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n276), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n305), .B1(new_n361), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT13), .B1(new_n196), .B2(G143), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(new_n327), .ZN(new_n380));
  XNOR2_X1  g194(.A(G128), .B(G143), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G116), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n240), .A2(G122), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n255), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n220), .A2(new_n221), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT94), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n386), .B2(new_n389), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n382), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n303), .A2(new_n394), .A3(G953), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n381), .B(new_n327), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n385), .A2(KEYINPUT14), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n384), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n385), .A2(KEYINPUT14), .ZN(new_n399));
  OAI21_X1  g213(.A(G107), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT95), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n386), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n255), .A2(KEYINPUT95), .A3(new_n384), .A4(new_n385), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n396), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n393), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n395), .B1(new_n393), .B2(new_n404), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G902), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT96), .B1(new_n408), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  OR3_X1    g229(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n419), .A2(G952), .A3(new_n214), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT97), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT98), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G475), .ZN(new_n427));
  INV_X1    g241(.A(G140), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n202), .A2(G140), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT16), .ZN(new_n431));
  OR3_X1    g245(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n431), .A2(G146), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(G146), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(G237), .A2(G953), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(G143), .A3(G214), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G143), .B1(new_n436), .B2(G214), .ZN(new_n439));
  OAI21_X1  g253(.A(G131), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT17), .ZN(new_n441));
  INV_X1    g255(.A(G237), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n214), .A3(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n207), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n334), .A3(new_n437), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT17), .B(G131), .C1(new_n438), .C2(new_n439), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n437), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(KEYINPUT92), .A3(KEYINPUT17), .A4(G131), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n435), .A2(new_n446), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G113), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n218), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n429), .A2(new_n430), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G146), .ZN(new_n456));
  XNOR2_X1  g270(.A(G125), .B(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n198), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT18), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n334), .ZN(new_n461));
  OAI221_X1 g275(.A(new_n459), .B1(new_n450), .B2(new_n461), .C1(new_n440), .C2(new_n460), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n452), .A2(new_n454), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n452), .A2(new_n462), .ZN(new_n465));
  INV_X1    g279(.A(new_n454), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(KEYINPUT93), .B(new_n454), .C1(new_n452), .C2(new_n462), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n427), .B1(new_n469), .B2(new_n276), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n440), .A2(new_n445), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n457), .A2(KEYINPUT19), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n457), .A2(KEYINPUT19), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n198), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n431), .A2(new_n432), .A3(G146), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT79), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT79), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n431), .A2(new_n432), .A3(new_n479), .A4(G146), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n473), .A2(new_n476), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n466), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n463), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n472), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  AOI211_X1 g301(.A(KEYINPUT20), .B(new_n487), .C1(new_n483), .C2(new_n463), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n471), .A2(new_n490), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n418), .A2(new_n426), .A3(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n302), .A2(new_n378), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT80), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n495));
  OAI211_X1 g309(.A(KEYINPUT77), .B(KEYINPUT23), .C1(new_n196), .C2(G119), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n196), .B(G119), .C1(KEYINPUT77), .C2(KEYINPUT23), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT78), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(KEYINPUT78), .A3(G110), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G119), .B(G128), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT24), .B(G110), .Z(new_n505));
  AOI21_X1  g319(.A(new_n435), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n498), .A2(G110), .B1(new_n504), .B2(new_n505), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(new_n478), .A3(new_n480), .A4(new_n458), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G137), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n507), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n507), .B2(new_n509), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n495), .B(new_n276), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n394), .B1(G234), .B2(new_n276), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n512), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n507), .A2(new_n509), .A3(new_n513), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n495), .B1(new_n522), .B2(new_n276), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n494), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT25), .B1(new_n525), .B2(G902), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n516), .A4(new_n517), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n517), .A2(G902), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  XNOR2_X1  g345(.A(G134), .B(G137), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT65), .B1(new_n532), .B2(new_n334), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT65), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n327), .A2(G137), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n329), .A2(G134), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n534), .B(G131), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n335), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT68), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT68), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n533), .A2(new_n540), .A3(new_n537), .A4(new_n335), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n539), .A2(new_n322), .A3(new_n323), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n211), .A2(new_n336), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n531), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n201), .A2(new_n335), .A3(new_n533), .A4(new_n537), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(new_n531), .A3(new_n543), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n249), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n248), .A3(new_n543), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT70), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT26), .B(G101), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n436), .A2(G210), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n549), .B(new_n249), .C1(new_n544), .C2(new_n546), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n545), .A2(new_n543), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n548), .B1(new_n248), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT28), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT28), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT74), .B1(new_n548), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n548), .A2(KEYINPUT74), .A3(new_n563), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n559), .A2(KEYINPUT31), .B1(new_n567), .B2(new_n556), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n551), .A2(new_n557), .A3(new_n558), .A4(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(KEYINPUT73), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(KEYINPUT73), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G472), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n276), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT32), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT32), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n573), .A2(new_n577), .A3(new_n574), .A4(new_n276), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT76), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n248), .B1(new_n542), .B2(new_n543), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n548), .B1(new_n581), .B2(KEYINPUT75), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n583), .B(new_n248), .C1(new_n542), .C2(new_n543), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT28), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n548), .A2(KEYINPUT74), .A3(new_n563), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(new_n564), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n556), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n590), .A2(new_n276), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n551), .A2(new_n558), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n556), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(new_n557), .A3(new_n562), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n588), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n580), .B1(new_n596), .B2(G472), .ZN(new_n597));
  AOI211_X1 g411(.A(KEYINPUT76), .B(new_n574), .C1(new_n591), .C2(new_n595), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n530), .B1(new_n579), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n493), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  XNOR2_X1  g416(.A(new_n570), .B(KEYINPUT73), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n603), .B2(new_n568), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G472), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n356), .B1(new_n370), .B2(new_n339), .ZN(new_n606));
  INV_X1    g420(.A(new_n357), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n359), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(G469), .A3(new_n346), .ZN(new_n609));
  NAND2_X1  g423(.A1(G469), .A2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n373), .B1(new_n364), .B2(new_n371), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n612), .A2(G469), .A3(G902), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n304), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n530), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n393), .A2(new_n404), .ZN(new_n616));
  INV_X1    g430(.A(new_n395), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(G478), .B(G902), .C1(new_n618), .C2(new_n405), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT33), .B1(new_n395), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n406), .B2(new_n407), .ZN(new_n622));
  INV_X1    g436(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n618), .A2(new_n405), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n624), .A3(new_n276), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n619), .B1(new_n625), .B2(G478), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n491), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n301), .A2(new_n425), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n605), .A2(new_n615), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NOR2_X1   g445(.A1(new_n491), .A2(new_n417), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n301), .A2(new_n425), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n605), .A2(new_n615), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND3_X1  g450(.A1(new_n302), .A2(new_n378), .A3(new_n492), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n513), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n519), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n528), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n524), .A2(new_n527), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n605), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n574), .B1(new_n573), .B2(new_n276), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n575), .A3(new_n643), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n637), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  AOI21_X1  g465(.A(new_n577), .B1(new_n604), .B2(new_n574), .ZN(new_n652));
  INV_X1    g466(.A(new_n578), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n599), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n420), .B1(new_n422), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n491), .A2(new_n417), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n301), .A2(new_n657), .A3(new_n643), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n614), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  OAI21_X1  g475(.A(new_n556), .B1(new_n582), .B2(new_n584), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n559), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n574), .B1(new_n663), .B2(new_n276), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n652), .B2(new_n653), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n418), .A2(new_n491), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n643), .A3(new_n188), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n294), .A2(new_n300), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT38), .Z(new_n672));
  OR3_X1    g486(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT103), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n656), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n378), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  INV_X1    g494(.A(new_n656), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n626), .B(new_n681), .C1(new_n470), .C2(new_n489), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n275), .A2(new_n190), .A3(new_n293), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n189), .B1(new_n297), .B2(new_n299), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n683), .B(new_n187), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT104), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n301), .A2(new_n688), .A3(new_n683), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n378), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n654), .A3(new_n643), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OAI21_X1  g506(.A(G469), .B1(new_n612), .B2(G902), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n377), .A2(new_n304), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n377), .A2(new_n693), .A3(new_n696), .A4(new_n304), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n530), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n654), .A3(new_n699), .A4(new_n628), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n698), .A2(new_n654), .A3(new_n699), .A4(new_n633), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  AND4_X1   g518(.A1(new_n301), .A2(new_n695), .A3(new_n492), .A4(new_n697), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n524), .A2(new_n527), .A3(new_n642), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n579), .B2(new_n599), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NAND2_X1  g523(.A1(new_n574), .A2(new_n276), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n557), .B1(new_n585), .B2(new_n587), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(KEYINPUT31), .B2(new_n559), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n710), .B1(new_n603), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n645), .A2(new_n713), .A3(new_n530), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n187), .A2(new_n671), .A3(new_n491), .A4(new_n418), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n698), .A2(new_n425), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NOR4_X1   g531(.A1(new_n645), .A2(new_n713), .A3(new_n706), .A4(new_n682), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n301), .A3(new_n697), .A4(new_n695), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND3_X1  g534(.A1(new_n294), .A2(new_n300), .A3(new_n187), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n614), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n654), .A2(new_n699), .A3(new_n683), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n600), .A2(KEYINPUT42), .A3(new_n683), .A4(new_n722), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NAND4_X1  g542(.A1(new_n654), .A2(new_n699), .A3(new_n657), .A4(new_n722), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT106), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n600), .A2(new_n731), .A3(new_n657), .A4(new_n722), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  OAI21_X1  g548(.A(G469), .B1(new_n360), .B2(KEYINPUT45), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n360), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n610), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  OR3_X1    g555(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT108), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n613), .B1(new_n740), .B2(new_n741), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n304), .A3(new_n676), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT109), .Z(new_n747));
  NAND3_X1  g561(.A1(new_n471), .A2(new_n490), .A3(new_n626), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT43), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT110), .Z(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n605), .A3(new_n706), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(KEYINPUT44), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(KEYINPUT44), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n752), .A2(new_n753), .A3(new_n721), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  NAND2_X1  g570(.A1(new_n745), .A2(new_n304), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n745), .A2(KEYINPUT111), .A3(KEYINPUT47), .A4(new_n304), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n654), .A2(new_n699), .A3(new_n682), .A4(new_n721), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT112), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  NAND2_X1  g583(.A1(new_n377), .A2(new_n693), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT113), .Z(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT49), .Z(new_n772));
  NOR4_X1   g586(.A1(new_n530), .A2(new_n188), .A3(new_n305), .A4(new_n748), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n667), .A3(new_n672), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n721), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n698), .A2(new_n775), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n699), .A2(new_n776), .A3(new_n420), .A4(new_n667), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n491), .A2(new_n626), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n645), .A2(new_n713), .A3(new_n706), .ZN(new_n779));
  INV_X1    g593(.A(new_n420), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n749), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n777), .A2(new_n778), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n698), .A2(new_n188), .A3(new_n672), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n714), .A2(new_n781), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n786), .A2(KEYINPUT50), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT50), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n783), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n763), .B(new_n764), .C1(new_n304), .C2(new_n771), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n775), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT116), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n782), .A2(new_n600), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT48), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n777), .A2(new_n627), .ZN(new_n798));
  INV_X1    g612(.A(G952), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n695), .A2(new_n301), .A3(new_n697), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n799), .B(G953), .C1(new_n787), .C2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n794), .B2(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n524), .A2(new_n527), .A3(new_n642), .A4(new_n681), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n806), .B(new_n304), .C1(new_n611), .C2(new_n613), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n301), .A2(new_n491), .A3(new_n418), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n666), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n691), .A2(new_n660), .A3(new_n719), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n800), .A2(new_n718), .B1(new_n654), .B2(new_n659), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .A3(new_n691), .A4(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n418), .A2(new_n491), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n654), .A2(new_n817), .A3(new_n643), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n779), .A2(new_n627), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n614), .A2(new_n656), .A3(new_n721), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n732), .A2(new_n730), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n727), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n708), .A2(new_n700), .A3(new_n703), .A4(new_n716), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n627), .A2(new_n632), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n426), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n605), .A2(new_n615), .A3(new_n302), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n601), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n649), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n425), .A2(new_n695), .A3(new_n697), .A4(new_n715), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n707), .A2(new_n705), .B1(new_n832), .B2(new_n714), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n700), .A4(new_n703), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n805), .B1(new_n823), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n820), .A2(new_n821), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n733), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n644), .A2(new_n648), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n493), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n601), .A4(new_n829), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n725), .A2(new_n726), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n844), .A3(new_n824), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n700), .A2(new_n708), .A3(new_n703), .A4(new_n716), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n846), .B2(new_n727), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n816), .B(new_n842), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n836), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n823), .A2(new_n835), .A3(new_n805), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT118), .B1(new_n804), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT119), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n804), .A2(KEYINPUT118), .A3(new_n855), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n774), .B1(new_n859), .B2(new_n860), .ZN(G75));
  NOR2_X1   g675(.A1(new_n214), .A2(G952), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n849), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n276), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT56), .B1(new_n865), .B2(G210), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n295), .A2(new_n296), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n217), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n297), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT55), .Z(new_n870));
  OAI21_X1  g684(.A(new_n863), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n866), .B2(new_n870), .ZN(G51));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n836), .A2(new_n848), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT120), .B1(new_n849), .B2(KEYINPUT54), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n850), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n610), .B(KEYINPUT57), .Z(new_n878));
  AOI21_X1  g692(.A(new_n612), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n864), .A2(new_n276), .A3(new_n739), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n863), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT121), .B(new_n863), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(G54));
  AND3_X1   g699(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n863), .B1(new_n886), .B2(new_n484), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n484), .B2(new_n886), .ZN(G60));
  AND2_X1   g702(.A1(new_n622), .A2(new_n624), .ZN(new_n889));
  NAND2_X1  g703(.A1(G478), .A2(G902), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT59), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n855), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n877), .A2(new_n889), .A3(new_n891), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n863), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(new_n896), .A3(new_n863), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n892), .B1(new_n895), .B2(new_n897), .ZN(G63));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT60), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n864), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n863), .B1(new_n901), .B2(new_n522), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n641), .B2(new_n901), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g718(.A1(G224), .A2(G953), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n835), .A2(G953), .B1(new_n423), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n867), .B1(G898), .B2(new_n214), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT124), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n907), .B(new_n909), .ZN(G69));
  NAND2_X1  g724(.A1(new_n814), .A2(new_n691), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n727), .A3(new_n733), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n747), .B2(new_n754), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n747), .A2(new_n600), .A3(new_n715), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n214), .A4(new_n768), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n544), .A2(new_n546), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n474), .A2(new_n475), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT125), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n917), .B(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n916), .B(new_n920), .C1(new_n655), .C2(new_n214), .ZN(new_n921));
  INV_X1    g735(.A(new_n600), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n922), .A2(new_n677), .A3(new_n721), .A4(new_n827), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT126), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n679), .A2(new_n912), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n679), .A2(KEYINPUT62), .A3(new_n912), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n755), .A3(new_n768), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n214), .ZN(new_n931));
  INV_X1    g745(.A(new_n920), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n921), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n921), .A2(new_n937), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G72));
  INV_X1    g753(.A(new_n835), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n914), .A2(new_n915), .A3(new_n768), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT63), .Z(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT127), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n556), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n557), .B(new_n944), .C1(new_n930), .C2(new_n835), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n593), .A2(new_n559), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n852), .B2(new_n853), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n862), .B1(new_n950), .B2(new_n952), .ZN(G57));
endmodule


