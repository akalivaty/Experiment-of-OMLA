//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(G155gat), .B(G162gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n206), .B(new_n207), .C1(KEYINPUT2), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT2), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT76), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(G148gat), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  INV_X1    g021(.A(G155gat), .ZN(new_n223));
  INV_X1    g022(.A(G162gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n221), .A2(KEYINPUT78), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT78), .B1(new_n221), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n217), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n217), .B(new_n232), .C1(new_n228), .C2(new_n229), .ZN(new_n233));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G113gat), .B(G120gat), .Z(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n231), .A2(new_n233), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n241), .B(new_n217), .C1(new_n228), .C2(new_n229), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n221), .A2(new_n227), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT78), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n221), .A2(KEYINPUT78), .A3(new_n227), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n250), .A2(new_n251), .B1(new_n216), .B2(new_n209), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n243), .A2(new_n244), .A3(new_n247), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n230), .A2(new_n242), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n245), .ZN(new_n257));
  INV_X1    g056(.A(new_n244), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n253), .A2(new_n247), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(new_n255), .A3(new_n244), .A4(new_n243), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n205), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT39), .ZN(new_n264));
  INV_X1    g063(.A(new_n243), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n253), .A2(new_n247), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n264), .B(new_n258), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n244), .A3(new_n245), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n269), .B2(new_n268), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n244), .B1(new_n261), .B2(new_n243), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n205), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT40), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n205), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n272), .B2(new_n264), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n277), .B(KEYINPUT40), .C1(new_n272), .C2(new_n271), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G197gat), .ZN(new_n280));
  INV_X1    g079(.A(G204gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G211gat), .A2(G218gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(G211gat), .A2(G218gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT73), .B1(new_n289), .B2(new_n285), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(KEYINPUT72), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n282), .A2(new_n283), .B1(new_n286), .B2(new_n285), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n285), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G226gat), .ZN(new_n298));
  INV_X1    g097(.A(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n307), .A2(KEYINPUT67), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT67), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT66), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n318), .A2(new_n313), .A3(new_n315), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(G190gat), .B1(new_n313), .B2(KEYINPUT65), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT28), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n303), .B(new_n311), .C1(new_n323), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n307), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n303), .A2(KEYINPUT24), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT64), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n335), .B2(new_n337), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n333), .B1(new_n332), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n302), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n348), .A2(new_n298), .A3(new_n299), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n297), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n300), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n301), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n296), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G8gat), .B(G36gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT75), .ZN(new_n359));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n354), .A2(new_n357), .ZN(new_n365));
  INV_X1    g164(.A(new_n361), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n354), .A2(KEYINPUT30), .A3(new_n357), .A4(new_n361), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT31), .B(G50gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n297), .B1(new_n233), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n295), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n377), .B2(new_n292), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n288), .A2(new_n295), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT3), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n252), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G22gat), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n291), .B(new_n375), .C1(new_n294), .C2(new_n295), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n232), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n374), .B1(new_n385), .B2(new_n230), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n376), .B2(new_n387), .ZN(new_n388));
  AOI211_X1 g187(.A(KEYINPUT79), .B(new_n297), .C1(new_n233), .C2(new_n375), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n382), .B(new_n383), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n373), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G22gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n395), .A2(new_n396), .A3(new_n390), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n395), .B2(new_n390), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n390), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT81), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n396), .A3(new_n390), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n279), .A2(new_n369), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n260), .A2(new_n262), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n276), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n260), .A2(new_n262), .A3(new_n205), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n354), .A2(new_n416), .A3(new_n357), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n366), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n354), .B2(new_n357), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT38), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n362), .ZN(new_n421));
  INV_X1    g220(.A(new_n418), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n355), .A2(new_n297), .A3(new_n356), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n423), .A2(KEYINPUT37), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n296), .B1(new_n352), .B2(new_n353), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT38), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n421), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n412), .A2(new_n415), .A3(new_n420), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n399), .A2(new_n403), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n369), .B1(new_n410), .B2(new_n413), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n404), .A2(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G227gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n299), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n328), .A2(new_n347), .A3(new_n241), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n241), .B1(new_n328), .B2(new_n347), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  XOR2_X1   g239(.A(G15gat), .B(G43gat), .Z(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT70), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n439), .B(KEYINPUT32), .C1(new_n440), .C2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n447));
  INV_X1    g246(.A(new_n435), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n311), .A2(new_n303), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n320), .A2(new_n322), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n325), .A2(new_n326), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n317), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n345), .ZN(new_n454));
  INV_X1    g253(.A(new_n307), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n305), .A2(KEYINPUT23), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n329), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(new_n333), .B1(new_n334), .B2(new_n343), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n242), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n448), .B1(new_n460), .B2(new_n436), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT68), .B1(new_n461), .B2(KEYINPUT33), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT32), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n439), .A2(new_n467), .A3(new_n440), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n444), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n446), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n460), .A2(new_n448), .A3(new_n436), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT34), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n472), .B(new_n446), .C1(new_n466), .C2(new_n469), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT36), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n475), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n461), .A2(KEYINPUT33), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n445), .B1(new_n485), .B2(new_n467), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n486), .A2(new_n447), .A3(new_n462), .A4(new_n465), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n472), .B1(new_n487), .B2(new_n446), .ZN(new_n488));
  INV_X1    g287(.A(new_n475), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n429), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n369), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT83), .B1(new_n494), .B2(new_n408), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n411), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n415), .A2(new_n410), .A3(new_n409), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n492), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n479), .A2(new_n431), .A3(new_n429), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n433), .A2(new_n484), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n506));
  INV_X1    g305(.A(G57gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G64gat), .ZN(new_n508));
  INV_X1    g307(.A(G64gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G57gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512));
  AND2_X1   g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(G71gat), .A2(G78gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT89), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n520), .B(new_n512), .C1(new_n521), .C2(new_n506), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT90), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G127gat), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT86), .ZN(new_n536));
  INV_X1    g335(.A(G1gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(KEYINPUT86), .A3(G1gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT16), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n535), .A2(new_n540), .B1(new_n541), .B2(G8gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(G8gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n526), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT90), .B1(new_n519), .B2(new_n522), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT91), .B1(new_n525), .B2(new_n526), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n545), .B1(new_n551), .B2(new_n528), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n533), .A2(new_n534), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n533), .B2(new_n534), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n223), .ZN(new_n558));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G29gat), .A2(G36gat), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G43gat), .B(G50gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT15), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G43gat), .B(G50gat), .Z(new_n573));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n566), .A3(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT85), .B1(new_n578), .B2(G36gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n568), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n572), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT17), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n585), .B(new_n572), .C1(new_n577), .C2(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n545), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n544), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n543), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n583), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT18), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n589), .B(KEYINPUT13), .Z(new_n597));
  INV_X1    g396(.A(new_n592), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n591), .A2(new_n583), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n595), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n588), .A2(new_n589), .A3(new_n592), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G197gat), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT11), .B(G169gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n603), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT7), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n611), .A2(new_n613), .A3(G85gat), .A4(G92gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(KEYINPUT92), .A3(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT93), .B1(G99gat), .B2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT8), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT94), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT93), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(KEYINPUT8), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n629));
  INV_X1    g428(.A(new_n622), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n617), .B1(new_n623), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G99gat), .B(G106gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT95), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(new_n617), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n633), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n583), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n587), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n648));
  AND2_X1   g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n647), .A2(new_n648), .B1(KEYINPUT41), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n647), .A2(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n652), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n644), .A2(new_n646), .A3(new_n657), .A4(new_n650), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n653), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n653), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n527), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n637), .B(new_n664), .C1(new_n638), .C2(new_n639), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n523), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n623), .A2(new_n631), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n667), .B2(new_n637), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n662), .A2(new_n663), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT10), .B1(new_n549), .B2(new_n550), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n645), .A3(KEYINPUT98), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n548), .B1(new_n546), .B2(new_n547), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n525), .A2(KEYINPUT91), .A3(new_n526), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n663), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n643), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n671), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n669), .B1(new_n645), .B2(new_n527), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n683), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n565), .A2(new_n609), .A3(new_n661), .A4(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n505), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n413), .A2(new_n410), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(new_n369), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n693), .A2(new_n369), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n699), .A2(new_n700), .B1(new_n701), .B2(G8gat), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(KEYINPUT99), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(KEYINPUT99), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n693), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n707), .A2(G15gat), .A3(new_n481), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n480), .A2(new_n709), .A3(new_n483), .ZN(new_n710));
  INV_X1    g509(.A(new_n483), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n482), .B1(new_n476), .B2(new_n478), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT100), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G15gat), .B1(new_n707), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n708), .A2(new_n716), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n693), .A2(new_n430), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(new_n661), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n501), .A2(new_n503), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n369), .A2(new_n275), .A3(new_n278), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n427), .A2(new_n420), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n429), .B(new_n723), .C1(new_n724), .C2(new_n498), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n432), .A2(new_n430), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n484), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n721), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n564), .A2(new_n609), .A3(new_n691), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(G29gat), .A3(new_n694), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT45), .Z(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT101), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n735), .B(KEYINPUT44), .C1(new_n504), .C2(new_n721), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n725), .A2(new_n726), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n713), .B2(new_n710), .ZN(new_n738));
  INV_X1    g537(.A(new_n722), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n733), .B(new_n661), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n734), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n695), .A3(new_n729), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G29gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n743), .ZN(G1328gat));
  NOR3_X1   g543(.A1(new_n730), .A2(G36gat), .A3(new_n493), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n741), .A2(new_n369), .A3(new_n729), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G36gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1329gat));
  NAND3_X1  g549(.A1(new_n741), .A2(new_n714), .A3(new_n729), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  OR3_X1    g551(.A1(new_n730), .A2(G43gat), .A3(new_n481), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT47), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n754), .B(new_n756), .ZN(G1330gat));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  INV_X1    g557(.A(new_n730), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n429), .A2(G50gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT104), .Z(new_n762));
  NAND3_X1  g561(.A1(new_n741), .A2(new_n430), .A3(new_n729), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(G50gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n759), .A2(KEYINPUT105), .A3(new_n760), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT105), .B1(new_n759), .B2(new_n760), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT48), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(G50gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n763), .B2(KEYINPUT106), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n741), .A2(new_n771), .A3(new_n430), .A4(new_n729), .ZN(new_n772));
  AOI211_X1 g571(.A(KEYINPUT107), .B(new_n768), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n763), .A2(KEYINPUT106), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(G50gat), .A3(new_n772), .ZN(new_n776));
  INV_X1    g575(.A(new_n768), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n765), .B1(new_n773), .B2(new_n778), .ZN(G1331gat));
  OAI21_X1  g578(.A(new_n722), .B1(new_n714), .B2(new_n737), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n661), .B1(new_n562), .B2(new_n563), .ZN(new_n781));
  AND4_X1   g580(.A1(new_n609), .A2(new_n780), .A3(new_n781), .A4(new_n691), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n695), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g583(.A(new_n493), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT108), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1333gat));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n714), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n481), .A2(G71gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(G71gat), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g592(.A1(new_n782), .A2(new_n430), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G78gat), .ZN(G1335gat));
  INV_X1    g594(.A(new_n609), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n564), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n661), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n661), .A3(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n799), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n691), .ZN(new_n806));
  INV_X1    g605(.A(G85gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n695), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n797), .ZN(new_n809));
  INV_X1    g608(.A(new_n691), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n741), .A2(new_n695), .A3(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n806), .A2(new_n808), .B1(new_n807), .B2(new_n812), .ZN(G1336gat));
  NOR2_X1   g612(.A1(new_n493), .A2(G92gat), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n806), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n741), .A2(new_n369), .A3(new_n811), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G92gat), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n798), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n815), .A2(new_n810), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n817), .A2(G92gat), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n816), .A2(new_n820), .B1(new_n823), .B2(new_n819), .ZN(G1337gat));
  XOR2_X1   g623(.A(KEYINPUT111), .B(G99gat), .Z(new_n825));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n481), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT112), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n805), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n741), .A2(new_n714), .A3(new_n811), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n825), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(G1338gat));
  NOR3_X1   g633(.A1(new_n810), .A2(new_n429), .A3(G106gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n805), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n741), .A2(new_n430), .A3(new_n811), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n835), .B(KEYINPUT113), .Z(new_n841));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT114), .B1(new_n843), .B2(KEYINPUT53), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845));
  AOI211_X1 g644(.A(new_n845), .B(new_n837), .C1(new_n839), .C2(new_n842), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n844), .B2(new_n846), .ZN(G1339gat));
  OAI21_X1  g646(.A(KEYINPUT98), .B1(new_n672), .B2(new_n645), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n642), .A2(new_n636), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n677), .A2(new_n849), .A3(new_n674), .A4(new_n635), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n848), .A2(new_n850), .B1(new_n682), .B2(new_n663), .ZN(new_n851));
  INV_X1    g650(.A(new_n680), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n681), .A2(new_n853), .A3(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n850), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n671), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n687), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n858), .A3(KEYINPUT55), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n690), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT54), .B1(new_n851), .B2(new_n852), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n855), .A2(new_n852), .A3(new_n671), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n679), .A2(new_n857), .A3(new_n680), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n688), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n596), .A2(new_n608), .A3(new_n600), .A4(new_n602), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n598), .A2(new_n599), .A3(new_n597), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n589), .B1(new_n588), .B2(new_n592), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n607), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n659), .A2(new_n660), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n860), .A2(new_n861), .A3(new_n868), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n868), .A2(new_n690), .A3(new_n859), .A4(new_n874), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n868), .A2(new_n796), .A3(new_n690), .A4(new_n859), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n691), .A2(new_n869), .A3(new_n872), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n661), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n565), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n781), .A2(new_n609), .A3(new_n810), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT115), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n781), .A2(new_n885), .A3(new_n609), .A4(new_n810), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n430), .B(new_n481), .C1(new_n882), .C2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n695), .A3(new_n493), .ZN(new_n889));
  INV_X1    g688(.A(G113gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n889), .A2(new_n890), .A3(new_n609), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n694), .B1(new_n882), .B2(new_n887), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n479), .A2(new_n429), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n369), .ZN(new_n895));
  AOI21_X1  g694(.A(G113gat), .B1(new_n895), .B2(new_n796), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n891), .A2(new_n896), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n889), .A2(new_n898), .A3(new_n810), .ZN(new_n899));
  AOI21_X1  g698(.A(G120gat), .B1(new_n895), .B2(new_n691), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1341gat));
  OAI21_X1  g700(.A(G127gat), .B1(new_n889), .B2(new_n565), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(new_n532), .A3(new_n564), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1342gat));
  NAND2_X1  g703(.A1(new_n493), .A2(new_n661), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT117), .Z(new_n906));
  OR3_X1    g705(.A1(new_n894), .A2(G134gat), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g707(.A(G134gat), .B1(new_n889), .B2(new_n721), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G1343gat));
  NOR3_X1   g710(.A1(new_n714), .A2(new_n694), .A3(new_n369), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n882), .A2(new_n887), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n430), .ZN(new_n914));
  INV_X1    g713(.A(new_n887), .ZN(new_n915));
  INV_X1    g714(.A(new_n878), .ZN(new_n916));
  INV_X1    g715(.A(new_n880), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n796), .A2(new_n859), .A3(new_n690), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n865), .B2(new_n867), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n854), .A2(new_n858), .A3(KEYINPUT119), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n862), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(KEYINPUT120), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n920), .A2(new_n924), .A3(new_n862), .A4(new_n921), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n917), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n916), .B1(new_n926), .B2(new_n661), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n915), .B1(new_n927), .B2(new_n565), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n430), .A2(KEYINPUT57), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n914), .A2(KEYINPUT118), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n430), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n931), .A2(KEYINPUT118), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n796), .B(new_n912), .C1(new_n930), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n218), .A2(new_n219), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT121), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n714), .A2(new_n429), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n892), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n369), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n212), .A3(new_n796), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n942), .A3(KEYINPUT58), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n936), .B(new_n941), .C1(KEYINPUT121), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1344gat));
  OAI21_X1  g745(.A(new_n912), .B1(new_n930), .B2(new_n933), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n810), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n210), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n912), .B(KEYINPUT122), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n876), .B1(new_n926), .B2(new_n661), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n565), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n883), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT57), .B1(new_n953), .B2(new_n430), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n931), .A2(new_n932), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n691), .B(new_n950), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n210), .B1(new_n956), .B2(KEYINPUT59), .ZN(new_n957));
  AOI21_X1  g756(.A(G148gat), .B1(new_n940), .B2(new_n691), .ZN(new_n958));
  OAI22_X1  g757(.A1(new_n949), .A2(KEYINPUT59), .B1(new_n957), .B2(new_n958), .ZN(G1345gat));
  OAI21_X1  g758(.A(G155gat), .B1(new_n947), .B2(new_n565), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n940), .A2(new_n223), .A3(new_n564), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1346gat));
  OAI21_X1  g761(.A(G162gat), .B1(new_n947), .B2(new_n721), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n906), .A2(G162gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n939), .B2(new_n964), .ZN(G1347gat));
  AOI21_X1  g764(.A(new_n695), .B1(new_n882), .B2(new_n887), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n893), .A2(new_n369), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G169gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n970), .A3(new_n796), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n695), .A2(new_n493), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n888), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n888), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n796), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n972), .B1(new_n980), .B2(G169gat), .ZN(new_n981));
  AOI211_X1 g780(.A(KEYINPUT124), .B(new_n970), .C1(new_n979), .C2(new_n796), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n971), .B1(new_n981), .B2(new_n982), .ZN(G1348gat));
  OAI21_X1  g782(.A(G176gat), .B1(new_n978), .B2(new_n810), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n968), .A2(G176gat), .A3(new_n810), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1349gat));
  OAI21_X1  g785(.A(G183gat), .B1(new_n978), .B2(new_n565), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n968), .A2(new_n316), .A3(new_n565), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT60), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n987), .A2(new_n992), .A3(new_n989), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1350gat));
  INV_X1    g793(.A(G190gat), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n995), .B1(new_n979), .B2(new_n661), .ZN(new_n996));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n969), .A2(new_n995), .A3(new_n661), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(KEYINPUT125), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n998), .B(new_n999), .C1(new_n996), .C2(new_n1001), .ZN(G1351gat));
  AND3_X1   g801(.A1(new_n966), .A2(new_n369), .A3(new_n938), .ZN(new_n1003));
  AOI21_X1  g802(.A(G197gat), .B1(new_n1003), .B2(new_n796), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n954), .A2(new_n955), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n715), .A2(new_n973), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n609), .A2(new_n280), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G1352gat));
  NAND3_X1  g808(.A1(new_n1003), .A2(new_n281), .A3(new_n691), .ZN(new_n1010));
  XOR2_X1   g809(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1011));
  XNOR2_X1  g810(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NOR3_X1   g811(.A1(new_n1005), .A2(new_n810), .A3(new_n1006), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1012), .B1(new_n1013), .B2(new_n281), .ZN(G1353gat));
  INV_X1    g813(.A(G211gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1003), .A2(new_n1015), .A3(new_n564), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1006), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n564), .B(new_n1017), .C1(new_n954), .C2(new_n955), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(G1354gat));
  AOI21_X1  g820(.A(G218gat), .B1(new_n1003), .B2(new_n661), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n661), .A2(G218gat), .ZN(new_n1023));
  XNOR2_X1  g822(.A(new_n1023), .B(KEYINPUT127), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1022), .B1(new_n1007), .B2(new_n1024), .ZN(G1355gat));
endmodule


