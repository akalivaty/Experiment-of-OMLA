

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799;

  INV_X1 U377 ( .A(n583), .ZN(n355) );
  INV_X1 U378 ( .A(n729), .ZN(n575) );
  XNOR2_X1 U379 ( .A(n372), .B(n492), .ZN(n594) );
  AND2_X1 U380 ( .A1(n552), .A2(n722), .ZN(n728) );
  XNOR2_X1 U381 ( .A(n483), .B(KEYINPUT95), .ZN(n787) );
  XNOR2_X1 U382 ( .A(n440), .B(G146), .ZN(n499) );
  INV_X1 U383 ( .A(n643), .ZN(n755) );
  NAND2_X1 U384 ( .A1(n356), .A2(n643), .ZN(n651) );
  XNOR2_X2 U385 ( .A(n584), .B(n355), .ZN(n643) );
  NOR2_X1 U386 ( .A1(n641), .A2(n384), .ZN(n356) );
  NOR2_X1 U387 ( .A1(n556), .A2(n564), .ZN(n569) );
  XNOR2_X2 U388 ( .A(n549), .B(KEYINPUT22), .ZN(n556) );
  XNOR2_X1 U389 ( .A(G101), .B(G107), .ZN(n464) );
  NAND2_X1 U390 ( .A1(n573), .A2(n566), .ZN(n740) );
  BUF_X1 U391 ( .A(n552), .Z(n723) );
  INV_X1 U392 ( .A(G953), .ZN(n789) );
  AND2_X2 U393 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X2 U394 ( .A(n776), .B(n410), .ZN(n689) );
  XNOR2_X1 U395 ( .A(n568), .B(KEYINPUT35), .ZN(n425) );
  NAND2_X2 U396 ( .A1(n398), .A2(n395), .ZN(n761) );
  XNOR2_X1 U397 ( .A(n787), .B(n470), .ZN(n682) );
  INV_X1 U398 ( .A(KEYINPUT16), .ZN(n381) );
  INV_X1 U399 ( .A(KEYINPUT45), .ZN(n583) );
  INV_X1 U400 ( .A(G125), .ZN(n440) );
  AND2_X1 U401 ( .A1(n424), .A2(n582), .ZN(n383) );
  AND2_X1 U402 ( .A1(n394), .A2(n389), .ZN(n393) );
  XNOR2_X1 U403 ( .A(n510), .B(KEYINPUT39), .ZN(n585) );
  XNOR2_X1 U404 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U405 ( .A(n487), .B(n486), .ZN(n497) );
  XOR2_X1 U406 ( .A(G113), .B(G104), .Z(n523) );
  XNOR2_X1 U407 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n500) );
  XNOR2_X1 U408 ( .A(G137), .B(G134), .ZN(n460) );
  INV_X1 U409 ( .A(G131), .ZN(n459) );
  XNOR2_X1 U410 ( .A(n775), .B(n462), .ZN(n357) );
  INV_X2 U411 ( .A(KEYINPUT73), .ZN(n413) );
  XNOR2_X1 U412 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n462) );
  XNOR2_X1 U413 ( .A(n380), .B(n523), .ZN(n422) );
  XNOR2_X1 U414 ( .A(n514), .B(n381), .ZN(n380) );
  XNOR2_X1 U415 ( .A(n589), .B(n588), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n589), .B(n588), .ZN(n688) );
  XNOR2_X1 U417 ( .A(n555), .B(KEYINPUT106), .ZN(n798) );
  NAND2_X1 U418 ( .A1(n585), .A2(n711), .ZN(n589) );
  BUF_X1 U419 ( .A(n798), .Z(n359) );
  XNOR2_X1 U420 ( .A(n775), .B(n462), .ZN(n504) );
  INV_X2 U421 ( .A(n562), .ZN(n548) );
  XNOR2_X1 U422 ( .A(n594), .B(n371), .ZN(n609) );
  INV_X1 U423 ( .A(KEYINPUT6), .ZN(n371) );
  NOR2_X1 U424 ( .A1(n622), .A2(n607), .ZN(n407) );
  NAND2_X1 U425 ( .A1(n624), .A2(n623), .ZN(n388) );
  AND2_X1 U426 ( .A1(n606), .A2(n406), .ZN(n623) );
  XNOR2_X1 U427 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n445) );
  XNOR2_X1 U428 ( .A(G104), .B(KEYINPUT75), .ZN(n463) );
  XNOR2_X1 U429 ( .A(G146), .B(G140), .ZN(n466) );
  AND2_X1 U430 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U431 ( .A1(n575), .A2(n368), .ZN(n396) );
  INV_X1 U432 ( .A(n565), .ZN(n397) );
  NAND2_X1 U433 ( .A1(n669), .A2(n534), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n455), .B(n454), .ZN(n552) );
  NAND2_X1 U435 ( .A1(n665), .A2(n534), .ZN(n455) );
  XOR2_X1 U436 ( .A(G146), .B(G113), .Z(n489) );
  XOR2_X1 U437 ( .A(KEYINPUT3), .B(G119), .Z(n486) );
  INV_X1 U438 ( .A(KEYINPUT70), .ZN(n484) );
  XNOR2_X1 U439 ( .A(G128), .B(G119), .ZN(n443) );
  XNOR2_X1 U440 ( .A(G137), .B(G110), .ZN(n448) );
  XNOR2_X1 U441 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n447) );
  INV_X1 U442 ( .A(KEYINPUT10), .ZN(n441) );
  AND2_X1 U443 ( .A1(n657), .A2(n360), .ZN(n659) );
  XNOR2_X1 U444 ( .A(n411), .B(n369), .ZN(n762) );
  NOR2_X1 U445 ( .A1(n740), .A2(n625), .ZN(n412) );
  NAND2_X1 U446 ( .A1(n390), .A2(n548), .ZN(n382) );
  XNOR2_X1 U447 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n599) );
  AND2_X1 U448 ( .A1(n618), .A2(n367), .ZN(n406) );
  NAND2_X1 U449 ( .A1(n425), .A2(n373), .ZN(n427) );
  INV_X1 U450 ( .A(KEYINPUT44), .ZN(n373) );
  AND2_X1 U451 ( .A1(n434), .A2(n545), .ZN(n431) );
  INV_X1 U452 ( .A(G902), .ZN(n534) );
  XNOR2_X1 U453 ( .A(G116), .B(G101), .ZN(n485) );
  XNOR2_X1 U454 ( .A(G143), .B(G131), .ZN(n524) );
  INV_X1 U455 ( .A(KEYINPUT65), .ZN(n652) );
  XOR2_X1 U456 ( .A(KEYINPUT76), .B(KEYINPUT89), .Z(n501) );
  OR2_X1 U457 ( .A1(G237), .A2(G902), .ZN(n506) );
  AND2_X1 U458 ( .A1(n479), .A2(n481), .ZN(n419) );
  NAND2_X1 U459 ( .A1(n625), .A2(n362), .ZN(n437) );
  NAND2_X1 U460 ( .A1(n430), .A2(n365), .ZN(n435) );
  INV_X1 U461 ( .A(n609), .ZN(n564) );
  AND2_X1 U462 ( .A1(n546), .A2(n722), .ZN(n547) );
  XNOR2_X1 U463 ( .A(G134), .B(G116), .ZN(n515) );
  NAND2_X1 U464 ( .A1(n379), .A2(n361), .ZN(n510) );
  NOR2_X1 U465 ( .A1(n612), .A2(n611), .ZN(n627) );
  NOR2_X1 U466 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U467 ( .A(n491), .B(n490), .ZN(n669) );
  XNOR2_X1 U468 ( .A(n483), .B(n482), .ZN(n491) );
  XNOR2_X1 U469 ( .A(n405), .B(n402), .ZN(n665) );
  AND2_X1 U470 ( .A1(n666), .A2(G953), .ZN(n774) );
  XNOR2_X1 U471 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U472 ( .A(n689), .B(n690), .ZN(n691) );
  INV_X1 U473 ( .A(n660), .ZN(n760) );
  NOR2_X1 U474 ( .A1(n408), .A2(n601), .ZN(n709) );
  INV_X1 U475 ( .A(G122), .ZN(n374) );
  AND2_X1 U476 ( .A1(n656), .A2(KEYINPUT2), .ZN(n360) );
  XOR2_X1 U477 ( .A(n508), .B(n509), .Z(n361) );
  XNOR2_X1 U478 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n362) );
  OR2_X1 U479 ( .A1(n656), .A2(n637), .ZN(n363) );
  AND2_X1 U480 ( .A1(n435), .A2(n433), .ZN(n364) );
  NAND2_X1 U481 ( .A1(n436), .A2(n435), .ZN(n601) );
  NOR2_X1 U482 ( .A1(n625), .A2(n362), .ZN(n365) );
  NAND2_X1 U483 ( .A1(n640), .A2(n639), .ZN(n366) );
  AND2_X1 U484 ( .A1(n605), .A2(n407), .ZN(n367) );
  XNOR2_X1 U485 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n368) );
  XOR2_X1 U486 ( .A(KEYINPUT112), .B(KEYINPUT41), .Z(n369) );
  INV_X1 U487 ( .A(KEYINPUT34), .ZN(n401) );
  OR2_X1 U488 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n370) );
  XNOR2_X1 U489 ( .A(KEYINPUT15), .B(G902), .ZN(n647) );
  XNOR2_X2 U490 ( .A(n414), .B(n461), .ZN(n483) );
  XNOR2_X2 U491 ( .A(n376), .B(KEYINPUT4), .ZN(n414) );
  XNOR2_X2 U492 ( .A(G143), .B(G128), .ZN(n376) );
  XNOR2_X1 U493 ( .A(n425), .B(n374), .ZN(G24) );
  XNOR2_X1 U494 ( .A(n376), .B(n375), .ZN(n516) );
  INV_X1 U495 ( .A(KEYINPUT103), .ZN(n375) );
  NAND2_X1 U496 ( .A1(n657), .A2(n656), .ZN(n377) );
  XNOR2_X1 U497 ( .A(n377), .B(KEYINPUT82), .ZN(n788) );
  NAND2_X1 U498 ( .A1(n728), .A2(n378), .ZN(n472) );
  XNOR2_X2 U499 ( .A(n378), .B(KEYINPUT1), .ZN(n729) );
  NAND2_X1 U500 ( .A1(n596), .A2(n378), .ZN(n408) );
  XNOR2_X2 U501 ( .A(n471), .B(G469), .ZN(n378) );
  NAND2_X1 U502 ( .A1(n379), .A2(n621), .ZN(n707) );
  NOR2_X2 U503 ( .A1(n415), .A2(n420), .ZN(n379) );
  NAND2_X1 U504 ( .A1(n385), .A2(n386), .ZN(n562) );
  NOR2_X2 U505 ( .A1(n556), .A2(n729), .ZN(n551) );
  NAND2_X1 U506 ( .A1(n393), .A2(n382), .ZN(n567) );
  NAND2_X1 U507 ( .A1(n383), .A2(n426), .ZN(n584) );
  NAND2_X1 U508 ( .A1(n387), .A2(n363), .ZN(n384) );
  INV_X1 U509 ( .A(n388), .ZN(n655) );
  NAND2_X1 U510 ( .A1(n659), .A2(n643), .ZN(n660) );
  NAND2_X1 U511 ( .A1(n432), .A2(n431), .ZN(n385) );
  NAND2_X1 U512 ( .A1(n429), .A2(n428), .ZN(n386) );
  NAND2_X1 U513 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U514 ( .A1(n388), .A2(n366), .ZN(n387) );
  NAND2_X1 U515 ( .A1(n565), .A2(n368), .ZN(n400) );
  NAND2_X1 U516 ( .A1(n575), .A2(n368), .ZN(n399) );
  NAND2_X1 U517 ( .A1(n761), .A2(n401), .ZN(n389) );
  INV_X1 U518 ( .A(n395), .ZN(n391) );
  NAND2_X1 U519 ( .A1(n398), .A2(KEYINPUT34), .ZN(n392) );
  NAND2_X1 U520 ( .A1(n563), .A2(n401), .ZN(n394) );
  NAND2_X1 U521 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U522 ( .A(n531), .ZN(n786) );
  XNOR2_X1 U523 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X1 U524 ( .A(n449), .B(n448), .ZN(n403) );
  NAND2_X1 U525 ( .A1(n511), .A2(G221), .ZN(n404) );
  XNOR2_X1 U526 ( .A(n531), .B(n444), .ZN(n405) );
  NOR2_X1 U527 ( .A1(n762), .A2(n408), .ZN(n598) );
  XNOR2_X2 U528 ( .A(n409), .B(n507), .ZN(n538) );
  NAND2_X1 U529 ( .A1(n689), .A2(n647), .ZN(n409) );
  XNOR2_X1 U530 ( .A(n421), .B(n505), .ZN(n410) );
  XNOR2_X2 U531 ( .A(n422), .B(n497), .ZN(n776) );
  NOR2_X1 U532 ( .A1(n620), .A2(n508), .ZN(n621) );
  NAND2_X1 U533 ( .A1(n629), .A2(n508), .ZN(n721) );
  NAND2_X1 U534 ( .A1(n361), .A2(n412), .ZN(n411) );
  NAND2_X1 U535 ( .A1(n361), .A2(n738), .ZN(n741) );
  XNOR2_X2 U536 ( .A(n413), .B(G110), .ZN(n775) );
  XNOR2_X1 U537 ( .A(n414), .B(n504), .ZN(n421) );
  NAND2_X1 U538 ( .A1(n418), .A2(n416), .ZN(n415) );
  AND2_X1 U539 ( .A1(n496), .A2(n417), .ZN(n416) );
  OR2_X1 U540 ( .A1(n479), .A2(n481), .ZN(n417) );
  NAND2_X1 U541 ( .A1(n480), .A2(n419), .ZN(n418) );
  NOR2_X1 U542 ( .A1(n480), .A2(n481), .ZN(n420) );
  NAND2_X1 U543 ( .A1(n427), .A2(n425), .ZN(n424) );
  NAND2_X1 U544 ( .A1(n423), .A2(n427), .ZN(n426) );
  XNOR2_X1 U545 ( .A(n561), .B(n370), .ZN(n423) );
  NAND2_X1 U546 ( .A1(n433), .A2(n545), .ZN(n428) );
  NAND2_X1 U547 ( .A1(n364), .A2(n436), .ZN(n429) );
  INV_X1 U548 ( .A(n538), .ZN(n430) );
  INV_X1 U549 ( .A(n601), .ZN(n432) );
  NAND2_X1 U550 ( .A1(n544), .A2(KEYINPUT0), .ZN(n433) );
  NOR2_X1 U551 ( .A1(n508), .A2(n625), .ZN(n613) );
  INV_X1 U552 ( .A(n544), .ZN(n434) );
  NAND2_X1 U553 ( .A1(n538), .A2(n362), .ZN(n438) );
  XNOR2_X2 U554 ( .A(n663), .B(n662), .ZN(n769) );
  XOR2_X1 U555 ( .A(n489), .B(n488), .Z(n439) );
  NAND2_X1 U556 ( .A1(n688), .A2(n797), .ZN(n600) );
  INV_X1 U557 ( .A(KEYINPUT108), .ZN(n473) );
  INV_X1 U558 ( .A(n591), .ZN(n479) );
  XNOR2_X1 U559 ( .A(n497), .B(n439), .ZN(n490) );
  NAND2_X1 U560 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U561 ( .A(n441), .B(G140), .ZN(n442) );
  XNOR2_X1 U562 ( .A(n499), .B(n442), .ZN(n531) );
  XNOR2_X1 U563 ( .A(n443), .B(KEYINPUT24), .ZN(n444) );
  NAND2_X1 U564 ( .A1(n789), .A2(G234), .ZN(n446) );
  XNOR2_X1 U565 ( .A(n446), .B(n445), .ZN(n511) );
  XNOR2_X1 U566 ( .A(n447), .B(KEYINPUT23), .ZN(n449) );
  NAND2_X1 U567 ( .A1(n647), .A2(G234), .ZN(n451) );
  INV_X1 U568 ( .A(KEYINPUT20), .ZN(n450) );
  XNOR2_X1 U569 ( .A(n451), .B(n450), .ZN(n457) );
  INV_X1 U570 ( .A(n457), .ZN(n452) );
  AND2_X1 U571 ( .A1(n452), .A2(G217), .ZN(n453) );
  XNOR2_X1 U572 ( .A(n453), .B(KEYINPUT25), .ZN(n454) );
  INV_X1 U573 ( .A(G221), .ZN(n456) );
  OR2_X1 U574 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U575 ( .A(n458), .B(KEYINPUT21), .ZN(n590) );
  INV_X1 U576 ( .A(n590), .ZN(n722) );
  XNOR2_X1 U577 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U578 ( .A(n464), .B(n463), .ZN(n468) );
  NAND2_X1 U579 ( .A1(n789), .A2(G227), .ZN(n465) );
  XNOR2_X1 U580 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U581 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U582 ( .A(n357), .B(n469), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n682), .A2(n534), .ZN(n471) );
  XNOR2_X2 U584 ( .A(n472), .B(KEYINPUT98), .ZN(n577) );
  XNOR2_X1 U585 ( .A(n577), .B(n473), .ZN(n480) );
  XOR2_X1 U586 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n475) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n474) );
  XNOR2_X1 U588 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U589 ( .A1(G952), .A2(n476), .ZN(n751) );
  NOR2_X1 U590 ( .A1(n751), .A2(G953), .ZN(n543) );
  NAND2_X1 U591 ( .A1(G902), .A2(n476), .ZN(n540) );
  OR2_X1 U592 ( .A1(n789), .A2(n540), .ZN(n477) );
  NOR2_X1 U593 ( .A1(n477), .A2(G900), .ZN(n478) );
  NOR2_X1 U594 ( .A1(n543), .A2(n478), .ZN(n591) );
  INV_X1 U595 ( .A(KEYINPUT74), .ZN(n481) );
  NOR2_X1 U596 ( .A1(G953), .A2(G237), .ZN(n529) );
  NAND2_X1 U597 ( .A1(n529), .A2(G210), .ZN(n482) );
  XNOR2_X1 U598 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U599 ( .A(KEYINPUT5), .B(KEYINPUT100), .ZN(n488) );
  INV_X1 U600 ( .A(G472), .ZN(n492) );
  NAND2_X1 U601 ( .A1(n506), .A2(G214), .ZN(n493) );
  XOR2_X1 U602 ( .A(KEYINPUT90), .B(n493), .Z(n625) );
  OR2_X1 U603 ( .A1(n594), .A2(n625), .ZN(n495) );
  XNOR2_X1 U604 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n494) );
  XNOR2_X1 U605 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X2 U606 ( .A(G107), .B(G122), .Z(n514) );
  NAND2_X1 U607 ( .A1(G224), .A2(n789), .ZN(n498) );
  XNOR2_X1 U608 ( .A(n499), .B(n498), .ZN(n503) );
  XNOR2_X1 U609 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U610 ( .A(n503), .B(n502), .ZN(n505) );
  NAND2_X1 U611 ( .A1(n506), .A2(G210), .ZN(n507) );
  BUF_X1 U612 ( .A(n538), .Z(n508) );
  INV_X1 U613 ( .A(KEYINPUT38), .ZN(n509) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n513) );
  NAND2_X1 U615 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U616 ( .A(n513), .B(n512), .ZN(n519) );
  XNOR2_X1 U617 ( .A(n515), .B(n514), .ZN(n517) );
  XNOR2_X1 U618 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U619 ( .A(n519), .B(n518), .ZN(n771) );
  NOR2_X1 U620 ( .A1(G902), .A2(n771), .ZN(n520) );
  XOR2_X1 U621 ( .A(n520), .B(KEYINPUT104), .Z(n522) );
  INV_X1 U622 ( .A(G478), .ZN(n521) );
  XNOR2_X1 U623 ( .A(n522), .B(n521), .ZN(n573) );
  XNOR2_X1 U624 ( .A(n524), .B(n523), .ZN(n528) );
  XOR2_X1 U625 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n526) );
  XNOR2_X1 U626 ( .A(G122), .B(KEYINPUT12), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U628 ( .A(n528), .B(n527), .Z(n533) );
  NAND2_X1 U629 ( .A1(G214), .A2(n529), .ZN(n530) );
  XNOR2_X1 U630 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n533), .B(n532), .ZN(n675) );
  NAND2_X1 U632 ( .A1(n675), .A2(n534), .ZN(n537) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n535), .B(G475), .ZN(n536) );
  XNOR2_X1 U635 ( .A(n537), .B(n536), .ZN(n566) );
  INV_X1 U636 ( .A(n566), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n714) );
  NAND2_X1 U638 ( .A1(n585), .A2(n714), .ZN(n630) );
  XNOR2_X1 U639 ( .A(n630), .B(G134), .ZN(G36) );
  XOR2_X1 U640 ( .A(G898), .B(KEYINPUT92), .Z(n781) );
  NAND2_X1 U641 ( .A1(n781), .A2(G953), .ZN(n539) );
  XOR2_X1 U642 ( .A(KEYINPUT93), .B(n539), .Z(n777) );
  NOR2_X1 U643 ( .A1(n540), .A2(n777), .ZN(n541) );
  XNOR2_X1 U644 ( .A(n541), .B(KEYINPUT94), .ZN(n542) );
  NOR2_X1 U645 ( .A1(n543), .A2(n542), .ZN(n544) );
  INV_X1 U646 ( .A(KEYINPUT0), .ZN(n545) );
  INV_X1 U647 ( .A(n740), .ZN(n546) );
  NAND2_X1 U648 ( .A1(n548), .A2(n547), .ZN(n549) );
  INV_X1 U649 ( .A(KEYINPUT105), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n551), .B(n550), .ZN(n554) );
  INV_X1 U651 ( .A(n594), .ZN(n726) );
  NOR2_X1 U652 ( .A1(n726), .A2(n723), .ZN(n553) );
  XNOR2_X1 U653 ( .A(n729), .B(KEYINPUT88), .ZN(n616) );
  INV_X1 U654 ( .A(n616), .ZN(n557) );
  NOR2_X1 U655 ( .A1(n557), .A2(n723), .ZN(n558) );
  AND2_X1 U656 ( .A1(n569), .A2(n558), .ZN(n560) );
  XNOR2_X1 U657 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n559) );
  XNOR2_X1 U658 ( .A(n560), .B(n559), .ZN(n799) );
  NAND2_X1 U659 ( .A1(n798), .A2(n799), .ZN(n561) );
  BUF_X1 U660 ( .A(n562), .Z(n563) );
  NAND2_X1 U661 ( .A1(n564), .A2(n728), .ZN(n565) );
  NOR2_X1 U662 ( .A1(n573), .A2(n566), .ZN(n619) );
  NAND2_X1 U663 ( .A1(n567), .A2(n619), .ZN(n568) );
  INV_X1 U664 ( .A(n569), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n575), .A2(n723), .ZN(n570) );
  NOR2_X1 U666 ( .A1(n571), .A2(n570), .ZN(n697) );
  AND2_X1 U667 ( .A1(n573), .A2(n572), .ZN(n711) );
  NOR2_X1 U668 ( .A1(n711), .A2(n714), .ZN(n742) );
  NAND2_X1 U669 ( .A1(n726), .A2(n728), .ZN(n574) );
  NOR2_X1 U670 ( .A1(n575), .A2(n574), .ZN(n735) );
  NAND2_X1 U671 ( .A1(n735), .A2(n548), .ZN(n576) );
  XNOR2_X1 U672 ( .A(KEYINPUT31), .B(n576), .ZN(n715) );
  NOR2_X1 U673 ( .A1(n563), .A2(n577), .ZN(n578) );
  XNOR2_X1 U674 ( .A(n578), .B(KEYINPUT99), .ZN(n579) );
  NOR2_X1 U675 ( .A1(n726), .A2(n579), .ZN(n699) );
  NOR2_X1 U676 ( .A1(n715), .A2(n699), .ZN(n580) );
  NOR2_X1 U677 ( .A1(n742), .A2(n580), .ZN(n581) );
  NOR2_X1 U678 ( .A1(n697), .A2(n581), .ZN(n582) );
  XNOR2_X1 U679 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n587) );
  INV_X1 U680 ( .A(KEYINPUT110), .ZN(n586) );
  XNOR2_X1 U681 ( .A(n587), .B(n586), .ZN(n588) );
  INV_X1 U682 ( .A(n625), .ZN(n738) );
  OR2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U684 ( .A1(n723), .A2(n592), .ZN(n593) );
  XNOR2_X1 U685 ( .A(n593), .B(KEYINPUT69), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n594), .A2(n608), .ZN(n595) );
  XNOR2_X1 U687 ( .A(KEYINPUT28), .B(n595), .ZN(n596) );
  INV_X1 U688 ( .A(KEYINPUT42), .ZN(n597) );
  XNOR2_X1 U689 ( .A(n598), .B(n597), .ZN(n797) );
  XNOR2_X1 U690 ( .A(n600), .B(n599), .ZN(n624) );
  INV_X1 U691 ( .A(KEYINPUT47), .ZN(n602) );
  NOR2_X1 U692 ( .A1(n709), .A2(n602), .ZN(n603) );
  XOR2_X1 U693 ( .A(n603), .B(KEYINPUT78), .Z(n606) );
  NOR2_X1 U694 ( .A1(KEYINPUT47), .A2(n742), .ZN(n604) );
  NAND2_X1 U695 ( .A1(n709), .A2(n604), .ZN(n605) );
  AND2_X1 U696 ( .A1(KEYINPUT47), .A2(n742), .ZN(n607) );
  XOR2_X1 U697 ( .A(KEYINPUT86), .B(KEYINPUT36), .Z(n615) );
  INV_X1 U698 ( .A(n711), .ZN(n612) );
  NOR2_X1 U699 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U700 ( .A(n610), .B(KEYINPUT107), .ZN(n611) );
  NAND2_X1 U701 ( .A1(n627), .A2(n613), .ZN(n614) );
  XNOR2_X1 U702 ( .A(n615), .B(n614), .ZN(n617) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n718) );
  XNOR2_X1 U704 ( .A(n718), .B(KEYINPUT84), .ZN(n618) );
  INV_X1 U705 ( .A(n619), .ZN(n620) );
  INV_X1 U706 ( .A(n707), .ZN(n622) );
  NOR2_X1 U707 ( .A1(n729), .A2(n625), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  AND2_X1 U710 ( .A1(n721), .A2(n630), .ZN(n656) );
  XNOR2_X1 U711 ( .A(KEYINPUT68), .B(KEYINPUT48), .ZN(n654) );
  INV_X1 U712 ( .A(n654), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n632), .A2(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n656), .A2(n631), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n632), .A2(KEYINPUT82), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n655), .A2(n635), .ZN(n636) );
  INV_X1 U718 ( .A(n647), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n636), .A2(n644), .ZN(n641) );
  INV_X1 U720 ( .A(KEYINPUT82), .ZN(n637) );
  NOR2_X1 U721 ( .A1(n654), .A2(KEYINPUT82), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n656), .A2(n638), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n654), .A2(KEYINPUT82), .ZN(n639) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n658) );
  OR2_X1 U725 ( .A1(n658), .A2(KEYINPUT81), .ZN(n645) );
  OR2_X1 U726 ( .A1(n647), .A2(n645), .ZN(n649) );
  AND2_X1 U727 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n648) );
  AND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n655), .B(n654), .ZN(n657) );
  INV_X1 U733 ( .A(KEYINPUT64), .ZN(n662) );
  AND2_X1 U734 ( .A1(n770), .A2(G217), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n664), .B(n665), .ZN(n667) );
  INV_X1 U736 ( .A(G952), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n667), .A2(n774), .ZN(G66) );
  NAND2_X1 U738 ( .A1(n769), .A2(G472), .ZN(n671) );
  XOR2_X1 U739 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n668) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n672) );
  INV_X1 U741 ( .A(n774), .ZN(n693) );
  NAND2_X1 U742 ( .A1(n672), .A2(n693), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U744 ( .A1(n769), .A2(G475), .ZN(n677) );
  XOR2_X1 U745 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n674) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n678), .A2(n693), .ZN(n680) );
  INV_X1 U748 ( .A(KEYINPUT60), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(G60) );
  NAND2_X1 U750 ( .A1(n769), .A2(G469), .ZN(n684) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  XNOR2_X1 U752 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n685), .A2(n693), .ZN(n687) );
  INV_X1 U755 ( .A(KEYINPUT126), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(n686), .ZN(G54) );
  XNOR2_X1 U757 ( .A(n358), .B(G131), .ZN(G33) );
  NAND2_X1 U758 ( .A1(n769), .A2(G210), .ZN(n692) );
  XOR2_X1 U759 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n690) );
  XNOR2_X1 U760 ( .A(n692), .B(n691), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U762 ( .A(KEYINPUT125), .B(KEYINPUT56), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n696), .B(n695), .ZN(G51) );
  XOR2_X1 U764 ( .A(G101), .B(n697), .Z(G3) );
  NAND2_X1 U765 ( .A1(n699), .A2(n711), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n698), .B(G104), .ZN(G6) );
  XNOR2_X1 U767 ( .A(G107), .B(KEYINPUT27), .ZN(n703) );
  XOR2_X1 U768 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n701) );
  NAND2_X1 U769 ( .A1(n699), .A2(n714), .ZN(n700) );
  XNOR2_X1 U770 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U771 ( .A(n703), .B(n702), .ZN(G9) );
  XOR2_X1 U772 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n705) );
  NAND2_X1 U773 ( .A1(n714), .A2(n709), .ZN(n704) );
  XNOR2_X1 U774 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U775 ( .A(G128), .B(n706), .Z(G30) );
  XNOR2_X1 U776 ( .A(G143), .B(KEYINPUT116), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n708), .B(n707), .ZN(G45) );
  NAND2_X1 U778 ( .A1(n709), .A2(n711), .ZN(n710) );
  XNOR2_X1 U779 ( .A(n710), .B(G146), .ZN(G48) );
  XOR2_X1 U780 ( .A(G113), .B(KEYINPUT117), .Z(n713) );
  NAND2_X1 U781 ( .A1(n715), .A2(n711), .ZN(n712) );
  XNOR2_X1 U782 ( .A(n713), .B(n712), .ZN(G15) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U784 ( .A(n716), .B(KEYINPUT118), .ZN(n717) );
  XNOR2_X1 U785 ( .A(G116), .B(n717), .ZN(G18) );
  XNOR2_X1 U786 ( .A(KEYINPUT37), .B(KEYINPUT119), .ZN(n719) );
  XNOR2_X1 U787 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U788 ( .A(G125), .B(n720), .ZN(G27) );
  XNOR2_X1 U789 ( .A(G140), .B(n721), .ZN(G42) );
  XOR2_X1 U790 ( .A(KEYINPUT53), .B(KEYINPUT124), .Z(n768) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U792 ( .A(KEYINPUT49), .B(n724), .Z(n725) );
  NOR2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U794 ( .A(KEYINPUT120), .B(n727), .Z(n733) );
  NOR2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U796 ( .A(KEYINPUT121), .B(n730), .Z(n731) );
  XNOR2_X1 U797 ( .A(KEYINPUT50), .B(n731), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U799 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U800 ( .A(KEYINPUT51), .B(n736), .Z(n737) );
  NOR2_X1 U801 ( .A1(n762), .A2(n737), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n738), .A2(n361), .ZN(n739) );
  NOR2_X1 U803 ( .A1(n740), .A2(n739), .ZN(n744) );
  NOR2_X1 U804 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U805 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U806 ( .A1(n761), .A2(n745), .ZN(n746) );
  NOR2_X1 U807 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U808 ( .A(n748), .B(KEYINPUT122), .ZN(n749) );
  XNOR2_X1 U809 ( .A(KEYINPUT52), .B(n749), .ZN(n750) );
  NOR2_X1 U810 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U811 ( .A(KEYINPUT123), .B(n752), .Z(n753) );
  NOR2_X1 U812 ( .A1(G953), .A2(n753), .ZN(n766) );
  NAND2_X1 U813 ( .A1(n788), .A2(n658), .ZN(n754) );
  XNOR2_X1 U814 ( .A(n754), .B(KEYINPUT80), .ZN(n758) );
  BUF_X1 U815 ( .A(n755), .Z(n756) );
  NAND2_X1 U816 ( .A1(n658), .A2(n756), .ZN(n757) );
  NAND2_X1 U817 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U818 ( .A1(n760), .A2(n759), .ZN(n764) );
  NOR2_X1 U819 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U820 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U821 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U822 ( .A(n768), .B(n767), .ZN(G75) );
  BUF_X1 U823 ( .A(n769), .Z(n770) );
  NAND2_X1 U824 ( .A1(n770), .A2(G478), .ZN(n772) );
  XNOR2_X1 U825 ( .A(n772), .B(n771), .ZN(n773) );
  NOR2_X1 U826 ( .A1(n774), .A2(n773), .ZN(G63) );
  XNOR2_X1 U827 ( .A(n776), .B(n775), .ZN(n778) );
  NAND2_X1 U828 ( .A1(n778), .A2(n777), .ZN(n785) );
  NAND2_X1 U829 ( .A1(G953), .A2(G224), .ZN(n779) );
  XOR2_X1 U830 ( .A(KEYINPUT61), .B(n779), .Z(n780) );
  NOR2_X1 U831 ( .A1(n781), .A2(n780), .ZN(n783) );
  NOR2_X1 U832 ( .A1(G953), .A2(n756), .ZN(n782) );
  NOR2_X1 U833 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U834 ( .A(n785), .B(n784), .ZN(G69) );
  XNOR2_X1 U835 ( .A(n787), .B(n786), .ZN(n791) );
  XNOR2_X1 U836 ( .A(n788), .B(n791), .ZN(n790) );
  NAND2_X1 U837 ( .A1(n790), .A2(n789), .ZN(n796) );
  XOR2_X1 U838 ( .A(G227), .B(n791), .Z(n792) );
  XNOR2_X1 U839 ( .A(n792), .B(KEYINPUT127), .ZN(n793) );
  NAND2_X1 U840 ( .A1(n793), .A2(G900), .ZN(n794) );
  NAND2_X1 U841 ( .A1(n794), .A2(G953), .ZN(n795) );
  NAND2_X1 U842 ( .A1(n796), .A2(n795), .ZN(G72) );
  XNOR2_X1 U843 ( .A(G137), .B(n797), .ZN(G39) );
  XNOR2_X1 U844 ( .A(n359), .B(G110), .ZN(G12) );
  XNOR2_X1 U845 ( .A(n799), .B(G119), .ZN(G21) );
endmodule

