//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G77), .A2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G238), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n219), .A3(G68), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n215), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n210), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G250), .ZN(new_n231));
  NOR2_X1   g0031(.A1(G257), .A2(G264), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n204), .A2(new_n205), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n212), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  INV_X1    g0036(.A(G20), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI22_X1  g0038(.A1(new_n233), .A2(KEYINPUT0), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g0039(.A(new_n228), .B(new_n239), .C1(KEYINPUT0), .C2(new_n233), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G250), .B(G257), .Z(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT66), .ZN(new_n251));
  XOR2_X1   g0051(.A(G50), .B(G58), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n237), .A2(G33), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n259), .B1(new_n260), .B2(new_n261), .C1(new_n206), .C2(new_n237), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n236), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(new_n268), .B2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n264), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n212), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n267), .A2(new_n270), .A3(new_n271), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT9), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n271), .A2(new_n274), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(new_n270), .A4(new_n267), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G77), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT67), .B(G1698), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n285), .B2(new_n282), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n287), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI211_X1 g0094(.A(G1), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(G226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n276), .A2(new_n279), .B1(G200), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n291), .A2(G190), .A3(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n303));
  OR2_X1    g0103(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n291), .A2(new_n306), .A3(new_n298), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT70), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n310), .A3(new_n275), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n300), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n301), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n269), .A2(G68), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT12), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n268), .A2(G13), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n203), .A2(G20), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G13), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G1), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n321), .A2(KEYINPUT12), .A3(G20), .A4(new_n203), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  INV_X1    g0125(.A(new_n258), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n318), .B1(new_n261), .B2(new_n207), .C1(new_n326), .C2(new_n212), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n264), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n327), .B2(new_n264), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n331), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT11), .A3(new_n329), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n324), .A2(new_n332), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n338));
  OAI21_X1  g0138(.A(G226), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G232), .A2(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n282), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n289), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n295), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n297), .A2(G238), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n344), .A2(new_n349), .A3(new_n345), .A4(new_n346), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n309), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT78), .B(KEYINPUT14), .Z(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n350), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n306), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n336), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n336), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(G200), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n348), .A2(G190), .A3(new_n350), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  INV_X1    g0164(.A(new_n260), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n273), .ZN(new_n366));
  INV_X1    g0166(.A(new_n264), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G1), .B2(new_n237), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n368), .B2(new_n365), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g0173(.A(G33), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n237), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT79), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n237), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT80), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n280), .A2(new_n281), .A3(new_n378), .A4(G20), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n377), .A2(KEYINPUT79), .A3(new_n378), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n381), .A2(new_n383), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n372), .B1(new_n388), .B2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n367), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n282), .B2(new_n237), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n391), .B2(new_n384), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT16), .B1(new_n392), .B2(new_n371), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n369), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n297), .A2(G232), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n284), .A2(G223), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G226), .A2(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n375), .A2(new_n376), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(G33), .B2(G87), .ZN(new_n401));
  OAI211_X1 g0201(.A(G1), .B(G13), .C1(new_n374), .C2(new_n293), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n345), .B(new_n396), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n306), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(G169), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n364), .B1(new_n395), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n388), .A2(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n371), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n264), .A3(new_n394), .ZN(new_n409));
  INV_X1    g0209(.A(new_n369), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n403), .A2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n306), .B2(new_n403), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(KEYINPUT18), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n406), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n403), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n403), .A2(G200), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n409), .A2(new_n417), .A3(new_n410), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n395), .A2(KEYINPUT17), .A3(new_n417), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G232), .B1(new_n337), .B2(new_n338), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n217), .A2(new_n219), .A3(G1698), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n400), .ZN(new_n427));
  INV_X1    g0227(.A(G107), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n282), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n289), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT71), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n295), .B1(new_n297), .B2(G244), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n430), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n306), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT73), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT73), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n306), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n433), .A2(new_n434), .A3(G169), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n272), .A2(G77), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n368), .A2(new_n207), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n260), .A2(new_n326), .B1(new_n237), .B2(new_n207), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT72), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g0245(.A(KEYINPUT15), .B(G87), .Z(new_n446));
  INV_X1    g0246(.A(new_n261), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI221_X1 g0248(.A(KEYINPUT72), .B1(new_n237), .B2(new_n207), .C1(new_n260), .C2(new_n326), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI211_X1 g0250(.A(new_n441), .B(new_n442), .C1(new_n450), .C2(new_n264), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT74), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n440), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n441), .B1(new_n450), .B2(new_n264), .ZN(new_n454));
  INV_X1    g0254(.A(new_n442), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n430), .A2(new_n432), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT71), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n309), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT74), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n439), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n433), .A2(new_n434), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G200), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n451), .C1(new_n416), .C2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AND4_X1   g0267(.A1(new_n314), .A2(new_n363), .A3(new_n424), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT89), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n237), .B1(new_n342), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G87), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n224), .A3(new_n428), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n472), .A2(KEYINPUT87), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT87), .B1(new_n472), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n400), .A2(new_n237), .A3(G68), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n237), .A2(G33), .A3(G97), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n479), .A2(KEYINPUT88), .A3(new_n471), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT88), .B1(new_n479), .B2(new_n471), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n470), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n471), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(KEYINPUT88), .A3(new_n471), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(new_n375), .B2(new_n376), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n486), .A2(new_n487), .B1(G68), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n472), .A2(new_n474), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n472), .A2(KEYINPUT87), .A3(new_n474), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n494), .A3(KEYINPUT89), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n483), .A2(new_n495), .A3(new_n264), .ZN(new_n496));
  INV_X1    g0296(.A(new_n446), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n273), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G238), .B1(new_n337), .B2(new_n338), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G244), .A2(G1698), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n282), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT85), .B(G116), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n374), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n289), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n268), .A2(G45), .A3(G274), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT84), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n268), .A2(G45), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n402), .A2(G250), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n416), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n268), .A2(G33), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n272), .A2(new_n513), .A3(new_n236), .A4(new_n263), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(G200), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n499), .A2(new_n512), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n446), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n496), .A2(new_n498), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n510), .A2(new_n309), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n505), .A2(new_n306), .A3(new_n507), .A4(new_n509), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G250), .B1(new_n337), .B2(new_n338), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G257), .A2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n282), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n374), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n289), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g0331(.A1(KEYINPUT5), .A2(G41), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT5), .A2(G41), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n508), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n289), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G264), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(G274), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n531), .A2(new_n416), .A3(new_n536), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n317), .A2(new_n237), .A3(G107), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n543), .B(KEYINPUT25), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n428), .B2(new_n514), .ZN(new_n545));
  AND2_X1   g0345(.A1(KEYINPUT85), .A2(G116), .ZN(new_n546));
  NOR2_X1   g0346(.A1(KEYINPUT85), .A2(G116), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT23), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n237), .B2(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n428), .A2(KEYINPUT23), .A3(G20), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n548), .A2(new_n447), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n237), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n400), .A2(KEYINPUT22), .A3(new_n237), .A4(G87), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n552), .A2(new_n555), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n545), .B1(new_n561), .B2(new_n264), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n542), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n538), .A2(new_n309), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n531), .A2(new_n306), .A3(new_n536), .A4(new_n537), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n367), .B1(new_n558), .B2(new_n560), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n545), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n564), .B1(new_n563), .B2(new_n568), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n518), .B(new_n525), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(KEYINPUT5), .A2(G41), .ZN(new_n572));
  NOR2_X1   g0372(.A1(KEYINPUT5), .A2(G41), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n402), .B1(new_n574), .B2(new_n508), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n537), .B1(new_n575), .B2(new_n225), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n400), .A2(new_n284), .A3(G244), .ZN(new_n578));
  NOR2_X1   g0378(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(G244), .B1(KEYINPUT82), .B2(KEYINPUT4), .ZN(new_n581));
  OR2_X1    g0381(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(G250), .A2(G1698), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n400), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G283), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n580), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT83), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(new_n289), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n588), .B2(new_n289), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n577), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n514), .A2(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n272), .A2(new_n224), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT81), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n428), .B1(new_n379), .B2(new_n382), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n224), .A2(new_n428), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G97), .A2(G107), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n428), .A2(KEYINPUT6), .A3(G97), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n237), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n326), .A2(new_n207), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n600), .B1(new_n609), .B2(new_n367), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n416), .B(new_n576), .C1(new_n588), .C2(new_n289), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n588), .A2(new_n289), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n577), .ZN(new_n614));
  OAI21_X1  g0414(.A(G107), .B1(new_n391), .B2(new_n384), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n605), .A2(new_n606), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G20), .ZN(new_n617));
  INV_X1    g0417(.A(new_n608), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n264), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n614), .A2(new_n309), .B1(new_n620), .B2(new_n600), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n306), .B(new_n577), .C1(new_n590), .C2(new_n591), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n593), .A2(new_n612), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(G257), .B1(new_n337), .B2(new_n338), .ZN(new_n624));
  NAND2_X1  g0424(.A1(G264), .A2(G1698), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n400), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G303), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n282), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n626), .A2(new_n289), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G270), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n537), .B1(new_n575), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(G169), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n503), .A2(G20), .B1(new_n236), .B2(new_n263), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT20), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n587), .B(new_n237), .C1(G33), .C2(new_n224), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n633), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n321), .B(G20), .C1(new_n547), .C2(new_n546), .ZN(new_n638));
  INV_X1    g0438(.A(G116), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n514), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(G20), .B1(new_n546), .B2(new_n547), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n264), .A3(new_n636), .ZN(new_n643));
  NAND2_X1  g0443(.A1(KEYINPUT90), .A2(KEYINPUT20), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(new_n635), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n637), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT91), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT91), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n637), .A2(new_n641), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n632), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g0452(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n650), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT21), .B(G169), .C1(new_n629), .C2(new_n631), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n535), .A2(G270), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n626), .A2(new_n289), .A3(new_n628), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(G179), .A4(new_n537), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n652), .A2(new_n653), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n631), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n657), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G200), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(G190), .A3(new_n657), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n650), .A3(new_n648), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n623), .A2(new_n660), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n469), .A2(new_n571), .A3(new_n666), .ZN(G372));
  OAI21_X1  g0467(.A(new_n452), .B1(new_n440), .B2(new_n451), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n456), .A2(new_n460), .A3(KEYINPUT74), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n361), .A2(new_n670), .A3(new_n439), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n357), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT96), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n421), .A2(new_n422), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n357), .A3(KEYINPUT96), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n406), .A2(new_n414), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n305), .A2(new_n312), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT97), .B1(new_n682), .B2(new_n311), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n680), .B1(new_n677), .B2(new_n678), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT97), .ZN(new_n685));
  INV_X1    g0485(.A(new_n311), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT94), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n520), .A2(KEYINPUT94), .A3(new_n521), .A4(new_n522), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n496), .A2(new_n517), .A3(new_n516), .A4(new_n498), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n511), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n654), .A2(new_n659), .ZN(new_n697));
  INV_X1    g0497(.A(new_n653), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n697), .B(new_n568), .C1(new_n651), .C2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n696), .A2(new_n563), .A3(new_n623), .A4(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n621), .A2(new_n622), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT26), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n703));
  AND4_X1   g0503(.A1(new_n518), .A2(new_n701), .A3(new_n525), .A4(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n692), .B(new_n700), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n683), .A2(new_n687), .B1(new_n469), .B2(new_n706), .ZN(G369));
  OAI211_X1 g0507(.A(new_n697), .B(new_n665), .C1(new_n651), .C2(new_n698), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n320), .A2(G20), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n268), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n654), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT98), .ZN(new_n717));
  MUX2_X1   g0517(.A(new_n660), .B(new_n708), .S(new_n717), .Z(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n715), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n568), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n563), .A2(new_n568), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT93), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n715), .B1(new_n567), .B2(new_n545), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n569), .A2(new_n570), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n568), .B1(new_n732), .B2(new_n660), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n722), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(G399));
  NOR2_X1   g0535(.A1(new_n230), .A2(G41), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n474), .A2(G116), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n235), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n737), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  AND4_X1   g0543(.A1(new_n520), .A2(new_n521), .A3(new_n524), .A4(new_n523), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n621), .A2(new_n622), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n744), .A2(new_n695), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n703), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n701), .A2(new_n518), .A3(new_n688), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT26), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n692), .B(new_n700), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n743), .B1(new_n751), .B2(new_n722), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n705), .A2(new_n743), .A3(new_n722), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n571), .A2(new_n666), .A3(new_n715), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n510), .A2(new_n658), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n576), .B1(new_n588), .B2(new_n289), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n757), .A2(new_n531), .A3(new_n536), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n510), .A2(new_n306), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n592), .A2(new_n538), .A3(new_n662), .A4(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT30), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n759), .A2(KEYINPUT99), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n761), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(new_n715), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT31), .B1(new_n756), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n715), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT31), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n719), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n755), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n742), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n718), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n709), .A2(G45), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n737), .A2(G1), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n236), .B1(G20), .B2(new_n309), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n282), .B1(new_n787), .B2(new_n529), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n237), .A2(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n539), .A2(G179), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n237), .A2(new_n416), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n306), .A2(new_n539), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G283), .A2(new_n792), .B1(new_n795), .B2(G326), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n790), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n627), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n789), .A2(new_n784), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT102), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n788), .B(new_n798), .C1(G329), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n306), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G322), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n794), .A2(new_n789), .A3(KEYINPUT101), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT101), .B1(new_n794), .B2(new_n789), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT33), .B(G317), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT103), .Z(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n802), .A2(new_n789), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n801), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n795), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n816), .A2(new_n212), .B1(new_n814), .B2(new_n207), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n791), .A2(new_n428), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n797), .A2(new_n473), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n809), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n803), .B(KEYINPUT100), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n821), .A2(G68), .B1(new_n822), .B2(G58), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n787), .A2(new_n224), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n282), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n799), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT32), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n820), .A2(new_n823), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n783), .B1(new_n815), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n253), .A2(G45), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n230), .A2(new_n400), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(G45), .C2(new_n740), .ZN(new_n833));
  INV_X1    g0633(.A(G355), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n400), .A2(new_n229), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(G116), .B2(new_n229), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n777), .A2(new_n782), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n778), .A2(new_n781), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT104), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n721), .A2(new_n780), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n719), .B2(new_n718), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n840), .A2(new_n842), .ZN(G396));
  NAND2_X1  g0643(.A1(new_n456), .A2(new_n715), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n670), .B2(new_n439), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n466), .B2(new_n844), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n746), .A2(new_n703), .B1(new_n748), .B2(new_n749), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n588), .A2(new_n589), .A3(new_n289), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n576), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n612), .B1(new_n850), .B2(new_n539), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n699), .A2(new_n851), .A3(new_n563), .A4(new_n745), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n518), .A2(new_n688), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n692), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n722), .B(new_n846), .C1(new_n847), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT106), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT106), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n705), .A2(new_n857), .A3(new_n722), .A4(new_n846), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n706), .A2(new_n715), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(new_n846), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(new_n772), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n780), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n792), .A2(G68), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n212), .B2(new_n797), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT105), .Z(new_n866));
  AOI211_X1 g0666(.A(new_n282), .B(new_n866), .C1(G132), .C2(new_n800), .ZN(new_n867));
  INV_X1    g0667(.A(new_n814), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n821), .A2(G150), .B1(G159), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n822), .A2(G143), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n816), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT34), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n867), .B(new_n873), .C1(new_n202), .C2(new_n787), .ZN(new_n874));
  INV_X1    g0674(.A(G283), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n809), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n791), .A2(new_n473), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G303), .B2(new_n795), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n428), .B2(new_n797), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n824), .B(new_n879), .C1(new_n548), .C2(new_n868), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n800), .A2(G311), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n400), .B1(new_n804), .B2(G294), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n874), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n782), .A2(new_n775), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n884), .A2(new_n782), .B1(new_n207), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(new_n781), .C1(new_n776), .C2(new_n846), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n863), .A2(new_n887), .ZN(G384));
  INV_X1    g0688(.A(new_n754), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n468), .B1(new_n752), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n683), .B2(new_n687), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT108), .Z(new_n892));
  NAND3_X1  g0692(.A1(new_n362), .A2(new_n336), .A3(new_n715), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n336), .A2(new_n715), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n357), .A2(new_n361), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n462), .A2(new_n715), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n859), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n408), .A2(new_n264), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n389), .A2(KEYINPUT16), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n410), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n713), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n413), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n901), .B1(new_n906), .B2(new_n419), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n367), .B(new_n393), .C1(new_n389), .C2(KEYINPUT16), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n908), .A2(new_n369), .B1(new_n413), .B2(new_n905), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n909), .A2(new_n901), .A3(new_n419), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n905), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT38), .B(new_n911), .C1(new_n424), .C2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n675), .B2(new_n678), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n907), .A2(new_n910), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n900), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n678), .A2(new_n905), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n357), .A2(new_n715), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n913), .A2(new_n917), .A3(KEYINPUT39), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n915), .A2(new_n916), .A3(new_n914), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n395), .A2(new_n713), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n415), .B2(new_n423), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n909), .A2(new_n419), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n909), .A2(new_n901), .A3(new_n419), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n932), .B2(KEYINPUT39), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n919), .B(new_n921), .C1(new_n922), .C2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n892), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n768), .A2(new_n771), .ZN(new_n936));
  OR2_X1    g0736(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n936), .A2(new_n846), .A3(new_n896), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n848), .A2(new_n849), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n539), .B1(new_n939), .B2(new_n577), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n610), .A2(new_n611), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n745), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n708), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n744), .A2(new_n695), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(new_n727), .A3(new_n944), .A4(new_n722), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n770), .B1(new_n945), .B2(new_n769), .ZN(new_n946));
  INV_X1    g0746(.A(new_n771), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n846), .B(new_n896), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n938), .A2(new_n918), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT40), .B1(new_n932), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n468), .A2(new_n936), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(G330), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n935), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n268), .B2(new_n709), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n639), .B1(new_n616), .B2(KEYINPUT35), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n959), .B(new_n238), .C1(KEYINPUT35), .C2(new_n616), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  OAI21_X1  g0761(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n740), .A2(new_n962), .B1(G50), .B2(new_n203), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(G1), .A3(new_n320), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(new_n961), .A3(new_n964), .ZN(G367));
  INV_X1    g0765(.A(G317), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n816), .A2(new_n813), .B1(new_n799), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n797), .A2(new_n968), .A3(new_n639), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n821), .A2(G294), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n822), .A2(G303), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n968), .B1(new_n797), .B2(new_n503), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n791), .A2(new_n224), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n868), .A2(G283), .B1(new_n786), .B2(G107), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT110), .ZN(new_n977));
  OR4_X1    g0777(.A1(new_n400), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n787), .A2(new_n203), .ZN(new_n979));
  INV_X1    g0779(.A(new_n799), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G50), .A2(new_n868), .B1(new_n980), .B2(G137), .ZN(new_n981));
  INV_X1    g0781(.A(G143), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n981), .B1(new_n982), .B2(new_n816), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n979), .B(new_n983), .C1(G150), .C2(new_n804), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n202), .B2(new_n797), .C1(new_n826), .C2(new_n809), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n400), .B1(new_n791), .B2(new_n207), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT111), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n978), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n780), .B1(new_n989), .B2(new_n782), .ZN(new_n990));
  INV_X1    g0790(.A(new_n832), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n837), .B1(new_n229), .B2(new_n497), .C1(new_n248), .C2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n777), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n499), .A2(new_n516), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n715), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n696), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n692), .B2(new_n995), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n990), .B(new_n992), .C1(new_n993), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n779), .A2(G1), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n610), .A2(new_n715), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n623), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n701), .A2(new_n715), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n734), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT45), .Z(new_n1005));
  NAND3_X1  g0805(.A1(new_n733), .A2(new_n942), .A3(new_n722), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT44), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n731), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n730), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n660), .A2(new_n715), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n729), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n732), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n720), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n773), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n773), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n736), .B(KEYINPUT41), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n999), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n730), .A2(new_n1003), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n732), .B(new_n1013), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT42), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n568), .B1(new_n593), .B2(new_n612), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n722), .B1(new_n1025), .B2(new_n701), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1022), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT109), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1027), .A2(new_n1022), .A3(new_n1028), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1032), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n998), .B1(new_n1021), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(KEYINPUT112), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT112), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n998), .C1(new_n1021), .C2(new_n1038), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1042), .ZN(G387));
  OR2_X1    g0843(.A1(new_n773), .A2(new_n1017), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n736), .A3(new_n1018), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1017), .A2(new_n999), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n822), .A2(G317), .B1(G322), .B2(new_n795), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n627), .B2(new_n814), .C1(new_n813), .C2(new_n809), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT48), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n875), .B2(new_n787), .C1(new_n529), .C2(new_n797), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n980), .A2(G326), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n400), .B1(new_n792), .B2(new_n548), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n803), .A2(new_n212), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n816), .A2(new_n826), .B1(new_n814), .B2(new_n203), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n821), .B2(new_n365), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n797), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n282), .B(new_n975), .C1(G77), .C2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT113), .B(G150), .Z(new_n1062));
  AOI22_X1  g0862(.A1(new_n980), .A2(new_n1062), .B1(new_n786), .B2(new_n446), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n832), .B1(new_n245), .B2(new_n294), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n738), .B2(new_n835), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n203), .A2(new_n207), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n365), .A2(new_n212), .ZN(new_n1069));
  AOI211_X1 g0869(.A(G116), .B(new_n474), .C1(new_n1069), .C2(KEYINPUT50), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n294), .C1(KEYINPUT50), .C2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1067), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(G107), .B2(new_n229), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1065), .A2(new_n782), .B1(new_n837), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n729), .A2(new_n777), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n781), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1045), .A2(new_n1046), .A3(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(KEYINPUT114), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1009), .A2(new_n1078), .A3(new_n1011), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1005), .A2(new_n731), .A3(KEYINPUT114), .A4(new_n1008), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1018), .A3(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n736), .C1(new_n1018), .C2(new_n1012), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n837), .B1(new_n224), .B2(new_n229), .C1(new_n256), .C2(new_n991), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n804), .A2(G159), .B1(new_n795), .B2(G150), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n821), .A2(G50), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n814), .A2(new_n260), .B1(new_n799), .B2(new_n982), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n787), .A2(new_n207), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G68), .C2(new_n1060), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n400), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n816), .A2(new_n966), .B1(new_n803), .B2(new_n813), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT52), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1092), .A2(new_n1091), .B1(new_n821), .B2(G303), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n400), .B1(new_n786), .B2(new_n548), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n797), .A2(new_n875), .B1(new_n814), .B2(new_n529), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n818), .B(new_n1096), .C1(G322), .C2(new_n980), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1090), .A2(new_n877), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n780), .B1(new_n1099), .B2(new_n782), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1083), .B(new_n1100), .C1(new_n1003), .C2(new_n993), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1082), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT115), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1079), .A2(new_n1104), .A3(new_n1080), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n999), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1103), .A2(new_n1109), .ZN(G390));
  AOI21_X1  g0910(.A(new_n898), .B1(new_n856), .B2(new_n858), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n846), .C1(new_n946), .C2(new_n947), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n897), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n897), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1113), .A2(new_n897), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n751), .A2(new_n722), .A3(new_n846), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(new_n899), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1120), .A3(new_n1114), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n468), .A2(new_n936), .A3(G330), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n890), .B(new_n1123), .C1(new_n683), .C2(new_n687), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n922), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n933), .B1(new_n900), .B2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n922), .B1(new_n924), .B2(new_n931), .C1(new_n1120), .C2(new_n897), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1118), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1126), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1116), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1124), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1137), .A3(new_n736), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n933), .A2(new_n775), .ZN(new_n1139));
  INV_X1    g0939(.A(G132), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n803), .A2(new_n1140), .B1(new_n791), .B2(new_n212), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n809), .A2(new_n871), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G125), .C2(new_n800), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1144), .A2(KEYINPUT53), .B1(new_n826), .B2(new_n787), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n282), .B(new_n1145), .C1(KEYINPUT53), .C2(new_n1144), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n795), .A2(G128), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n868), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n864), .B1(new_n224), .B2(new_n814), .C1(new_n639), .C2(new_n803), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n819), .B(new_n1151), .C1(G283), .C2(new_n795), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n821), .A2(G107), .B1(G294), .B2(new_n800), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n207), .C2(new_n787), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1150), .B1(new_n1154), .B2(new_n400), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1155), .A2(new_n782), .B1(new_n260), .B2(new_n885), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1139), .A2(new_n781), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT116), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n999), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT116), .A4(new_n1107), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1138), .B(new_n1157), .C1(new_n1160), .C2(new_n1161), .ZN(G378));
  NAND2_X1  g0962(.A1(new_n953), .A2(G330), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n313), .A2(KEYINPUT55), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT55), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n305), .A2(new_n1165), .A3(new_n311), .A4(new_n312), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n275), .A2(new_n905), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT56), .Z(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT118), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n934), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1173), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n953), .A2(G330), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n953), .B2(G330), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n719), .B(new_n1173), .C1(new_n951), .C2(new_n952), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n934), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1137), .A2(new_n1125), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1183), .A3(KEYINPUT57), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n736), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1175), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1179), .A2(new_n1180), .A3(new_n934), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n999), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1171), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n775), .A3(new_n1169), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n885), .A2(new_n212), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n809), .A2(new_n1140), .B1(new_n871), .B2(new_n814), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT117), .Z(new_n1196));
  NAND2_X1  g0996(.A1(new_n804), .A2(G128), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n786), .A2(G150), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1060), .A2(new_n1148), .B1(new_n795), .B2(G125), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT59), .Z(new_n1201));
  AOI21_X1  g1001(.A(G41), .B1(new_n980), .B2(G124), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G33), .B1(new_n792), .B2(G159), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n212), .B1(new_n280), .B2(G41), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n809), .A2(new_n224), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n816), .A2(new_n639), .B1(new_n803), .B2(new_n428), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G58), .B2(new_n792), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n979), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n868), .A2(new_n446), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G41), .B(new_n400), .C1(new_n1060), .C2(G77), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1206), .B(new_n1212), .C1(G283), .C2(new_n800), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT58), .Z(new_n1214));
  NAND3_X1  g1014(.A1(new_n1204), .A2(new_n1205), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n780), .B1(new_n1215), .B2(new_n782), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1193), .A2(new_n1194), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1191), .A2(KEYINPUT119), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT119), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1107), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1217), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1188), .A2(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n885), .A2(new_n203), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n896), .A2(new_n776), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n804), .A2(G283), .B1(new_n795), .B2(G294), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n224), .B2(new_n797), .C1(new_n428), .C2(new_n814), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G77), .B2(new_n792), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n400), .B1(new_n786), .B2(new_n446), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n821), .A2(new_n548), .B1(G303), .B2(new_n800), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT120), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G159), .A2(new_n1060), .B1(new_n868), .B2(G150), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n212), .B2(new_n787), .C1(new_n1140), .C2(new_n816), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n282), .B(new_n1235), .C1(G58), .C2(new_n792), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n821), .A2(new_n1148), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n822), .A2(G137), .B1(new_n800), .B2(G128), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n783), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1226), .A2(new_n780), .A3(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1122), .A2(new_n999), .B1(new_n1225), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1124), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1020), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1244), .B2(new_n1136), .ZN(G381));
  INV_X1    g1045(.A(G378), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1188), .A2(new_n1223), .A3(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1247), .A2(G384), .A3(G381), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1040), .A2(new_n1249), .A3(new_n1042), .A4(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT121), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT121), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1248), .A2(new_n1254), .A3(new_n1251), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1253), .A2(new_n1255), .ZN(G407));
  OR2_X1    g1056(.A1(new_n1247), .A2(G343), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G213), .B(new_n1257), .C1(new_n1253), .C2(new_n1255), .ZN(G409));
  INV_X1    g1058(.A(new_n1039), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1250), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G390), .A2(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1249), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n998), .B1(new_n1021), .B2(new_n1038), .C1(new_n1102), .C2(new_n1108), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1249), .A2(new_n1039), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1261), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(new_n1250), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1260), .A2(KEYINPUT125), .A3(new_n1261), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1262), .A2(new_n1263), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1243), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1124), .A2(new_n1117), .A3(new_n1121), .A4(KEYINPUT60), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1126), .A3(new_n736), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1242), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(G384), .A3(new_n1242), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n714), .A2(G213), .A3(G2897), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT122), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1279), .A2(KEYINPUT122), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1281), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1276), .A2(G384), .A3(new_n1242), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1276), .B2(new_n1242), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT123), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT123), .A3(new_n1287), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1246), .B1(new_n1188), .B2(new_n1223), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n714), .A2(G213), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1182), .A2(new_n1183), .A3(new_n1020), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1191), .A3(new_n1217), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1299), .B2(G378), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1286), .B(new_n1295), .C1(new_n1296), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1296), .A2(new_n1293), .A3(new_n1300), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1301), .B(new_n1302), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1296), .A2(new_n1300), .A3(new_n1293), .A4(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1272), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1295), .A2(new_n1286), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT124), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1295), .A2(new_n1286), .A3(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1303), .B1(new_n1314), .B2(KEYINPUT63), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1272), .B2(KEYINPUT61), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1264), .A2(new_n1265), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1319));
  OAI211_X1 g1119(.A(KEYINPUT126), .B(new_n1302), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1303), .A2(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1308), .B1(new_n1315), .B2(new_n1323), .ZN(G405));
  NOR2_X1   g1124(.A1(G375), .A2(G378), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1279), .B(new_n1280), .C1(new_n1325), .C2(new_n1296), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G375), .A2(G378), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(new_n1247), .A3(new_n1293), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1272), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1329), .B(new_n1330), .ZN(G402));
endmodule


