//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(G22gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(G204gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G197gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G197gat), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n207), .C1(KEYINPUT22), .C2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G141gat), .B(G148gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n220), .B1(new_n224), .B2(KEYINPUT2), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n217), .B(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n216), .B1(KEYINPUT29), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n211), .B(new_n212), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT74), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n228), .B(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G228gat), .A3(G233gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT31), .B(G50gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n215), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT78), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n213), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT29), .B1(new_n214), .B2(KEYINPUT78), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT3), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n243), .B(new_n233), .C1(new_n248), .C2(new_n229), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n240), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n242), .B1(new_n240), .B2(new_n249), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n204), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n241), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n240), .A2(new_n242), .A3(new_n249), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n203), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n229), .A2(new_n237), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n228), .A2(KEYINPUT74), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n230), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G134gat), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT65), .B(G134gat), .Z(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  INV_X1    g064(.A(G113gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G120gat), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(G113gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n265), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n261), .A2(G134gat), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n272), .A2(new_n265), .A3(new_n262), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT66), .B1(new_n266), .B2(G120gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n268), .A3(G113gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n274), .B(new_n276), .C1(G113gat), .C2(new_n268), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n231), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n260), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n279), .B2(new_n228), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n264), .A2(new_n270), .B1(new_n273), .B2(new_n277), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n229), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G225gat), .A2(G233gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(KEYINPUT75), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n286), .A2(KEYINPUT39), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G1gat), .B(G29gat), .Z(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n295), .B(KEYINPUT79), .Z(new_n296));
  NOR2_X1   g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n279), .A2(new_n228), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n258), .A2(new_n259), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n279), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n289), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT39), .B(new_n301), .C1(new_n286), .C2(new_n289), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT40), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(G183gat), .B(G190gat), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n315));
  OR2_X1    g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT25), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(new_n313), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n308), .A2(new_n321), .A3(new_n322), .A4(new_n309), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n304), .A2(KEYINPUT26), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(new_n311), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n309), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n332), .A2(new_n304), .A3(KEYINPUT26), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n318), .B(new_n323), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(new_n235), .B1(G226gat), .B2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(G226gat), .A3(G233gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n234), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n216), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343));
  INV_X1    g142(.A(G64gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G92gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n338), .A2(new_n342), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT72), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n338), .A2(new_n342), .A3(new_n352), .A4(new_n348), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n234), .B1(new_n336), .B2(new_n337), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n341), .A2(new_n335), .A3(new_n216), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n348), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT71), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n303), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n282), .A2(new_n285), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n289), .C1(new_n260), .C2(new_n280), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n298), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(new_n238), .B2(new_n283), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n365), .B1(new_n369), .B2(new_n288), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT5), .B1(new_n300), .B2(new_n289), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n364), .A3(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n373), .A3(new_n296), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n371), .A2(new_n373), .A3(new_n376), .A4(new_n296), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n297), .A2(KEYINPUT40), .A3(new_n302), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n257), .B1(new_n362), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n295), .B1(new_n371), .B2(new_n373), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(KEYINPUT6), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n373), .A3(new_n295), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT6), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n350), .A2(new_n353), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT37), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT83), .B(new_n347), .C1(new_n357), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n338), .B2(new_n342), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n348), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n357), .A2(new_n392), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n378), .A2(KEYINPUT81), .A3(new_n383), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n386), .A2(new_n390), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n397), .ZN(new_n403));
  NOR4_X1   g202(.A1(new_n403), .A2(new_n348), .A3(new_n395), .A4(new_n399), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n381), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n339), .A2(new_n283), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n334), .A2(new_n279), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT34), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n406), .A2(new_n412), .A3(new_n409), .A4(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n406), .B2(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT32), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT67), .B(G71gat), .ZN(new_n419));
  INV_X1    g218(.A(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n415), .B2(KEYINPUT33), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n411), .B(new_n413), .C1(new_n416), .C2(new_n415), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n418), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n418), .B2(new_n426), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT69), .B1(new_n430), .B2(KEYINPUT36), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT36), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n432), .B(new_n433), .C1(new_n428), .C2(new_n429), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(KEYINPUT68), .A3(KEYINPUT36), .ZN(new_n436));
  INV_X1    g235(.A(new_n429), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT36), .A3(new_n427), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n359), .A2(new_n361), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n383), .A2(new_n387), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n389), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n257), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n405), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n252), .A2(new_n256), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT35), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n386), .A2(new_n390), .A3(new_n401), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT35), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .A4(new_n444), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT16), .ZN(new_n459));
  AOI21_X1  g258(.A(G1gat), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n460), .B(new_n462), .Z(new_n463));
  NAND2_X1  g262(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n460), .B(new_n462), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT89), .B(G8gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n472));
  INV_X1    g271(.A(G57gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G64gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n344), .A2(G57gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT92), .B(new_n471), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n479));
  XNOR2_X1  g278(.A(G57gat), .B(G64gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n472), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT91), .B1(new_n480), .B2(new_n472), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n471), .B1(new_n483), .B2(KEYINPUT92), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT21), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n208), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n208), .B1(new_n470), .B2(new_n486), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n488), .A2(new_n489), .B1(KEYINPUT21), .B2(new_n485), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n485), .A2(KEYINPUT21), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G127gat), .B(G155gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(KEYINPUT20), .Z(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT19), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT93), .B(G183gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n497), .B2(new_n499), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G134gat), .B(G162gat), .Z(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT94), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT41), .ZN(new_n513));
  INV_X1    g312(.A(G50gat), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n514), .A2(G43gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(G43gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT15), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(G43gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n514), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT15), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT85), .B(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n523), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n517), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n517), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(new_n524), .A3(new_n522), .A4(new_n525), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT87), .A3(KEYINPUT17), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n529), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G99gat), .B(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(G99gat), .B2(G106gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n346), .A2(KEYINPUT95), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G92gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G85gat), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n538), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(G85gat), .B1(new_n541), .B2(new_n543), .ZN(new_n554));
  NOR4_X1   g353(.A1(new_n554), .A2(new_n551), .A3(new_n537), .A4(new_n540), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n536), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT97), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n527), .B(new_n529), .C1(new_n553), .C2(new_n555), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n512), .A2(KEYINPUT41), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT96), .B1(new_n563), .B2(new_n564), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n513), .B1(new_n558), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n567), .A2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(new_n513), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n572), .A3(new_n557), .A4(new_n562), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n509), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n560), .A2(new_n561), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n570), .A2(new_n573), .A3(new_n509), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n570), .A2(new_n573), .A3(new_n509), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n579), .A2(new_n574), .B1(new_n561), .B2(new_n560), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n507), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n469), .B1(new_n531), .B2(new_n535), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n533), .B1(new_n465), .B2(new_n468), .ZN(new_n587));
  NOR4_X1   g386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n585), .B(KEYINPUT13), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n470), .A2(new_n533), .ZN(new_n590));
  INV_X1    g389(.A(new_n587), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT90), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n583), .A2(new_n587), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n585), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n584), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n591), .ZN(new_n597));
  INV_X1    g396(.A(new_n589), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n536), .A2(new_n470), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(KEYINPUT18), .A3(new_n585), .A4(new_n591), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n593), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT11), .B(G169gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G197gat), .ZN(new_n606));
  XOR2_X1   g405(.A(G113gat), .B(G141gat), .Z(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT84), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n596), .A2(new_n609), .A3(new_n599), .A4(new_n601), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT10), .B1(new_n553), .B2(new_n555), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT92), .B1(new_n476), .B2(new_n477), .ZN(new_n617));
  INV_X1    g416(.A(new_n471), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n481), .A3(new_n478), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n615), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  INV_X1    g421(.A(G106gat), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT8), .B1(new_n420), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT95), .B(G92gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(G85gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n537), .B1(new_n626), .B2(new_n551), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n546), .A2(new_n538), .A3(new_n552), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n485), .A2(new_n629), .A3(KEYINPUT101), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n554), .A2(new_n551), .A3(new_n540), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n538), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT99), .B(new_n537), .C1(new_n626), .C2(new_n551), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n485), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n482), .A2(new_n484), .B1(new_n553), .B2(new_n555), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G230gat), .ZN(new_n641));
  INV_X1    g440(.A(G233gat), .ZN(new_n642));
  OAI22_X1  g441(.A1(new_n631), .A2(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n644), .A3(new_n639), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  INV_X1    g446(.A(G176gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT103), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT104), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n643), .A2(new_n645), .A3(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT102), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n643), .A2(new_n656), .A3(new_n645), .A4(new_n650), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n614), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n457), .A2(new_n582), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n445), .A2(new_n389), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n661), .A2(KEYINPUT42), .A3(new_n443), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n443), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT105), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(G8gat), .ZN(new_n671));
  OAI221_X1 g470(.A(new_n667), .B1(KEYINPUT42), .B2(new_n666), .C1(new_n669), .C2(new_n671), .ZN(G1325gat));
  AOI21_X1  g471(.A(G15gat), .B1(new_n661), .B2(new_n430), .ZN(new_n673));
  INV_X1    g472(.A(new_n442), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n661), .A2(G15gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n257), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  AND2_X1   g478(.A1(new_n578), .A2(new_n580), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n448), .B2(new_n456), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n660), .A2(new_n507), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n662), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G29gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n685), .ZN(new_n689));
  INV_X1    g488(.A(new_n662), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(G29gat), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT45), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(G1328gat));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n443), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n521), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n689), .A2(new_n521), .A3(new_n444), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1329gat));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n674), .A3(new_n685), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n683), .A2(new_n701), .A3(new_n674), .A4(new_n685), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n518), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n689), .ZN(new_n704));
  INV_X1    g503(.A(new_n518), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n430), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(KEYINPUT47), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n706), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n699), .B2(new_n518), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(KEYINPUT47), .B2(new_n709), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n686), .A2(G50gat), .A3(new_n257), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n514), .B1(new_n689), .B2(new_n449), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g513(.A1(new_n582), .A2(new_n457), .A3(new_n614), .A4(new_n659), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n662), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G57gat), .ZN(G1332gat));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n715), .B(new_n443), .C1(new_n718), .C2(new_n344), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n344), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1333gat));
  NAND3_X1  g520(.A1(new_n715), .A2(G71gat), .A3(new_n674), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n715), .A2(new_n430), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(G71gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n726), .B(new_n722), .C1(new_n723), .C2(G71gat), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(KEYINPUT50), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT50), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1334gat));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n257), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g531(.A1(new_n457), .A2(new_n581), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n682), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n506), .A2(new_n613), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n734), .A2(new_n659), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n690), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n457), .A2(new_n581), .A3(new_n736), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n681), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n659), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n662), .A2(new_n545), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n744), .B2(new_n745), .ZN(G1336gat));
  INV_X1    g545(.A(new_n659), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(new_n444), .A3(G92gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n741), .B2(new_n742), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n625), .B1(new_n737), .B2(new_n444), .ZN(new_n753));
  INV_X1    g552(.A(new_n742), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n681), .B2(new_n736), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n748), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT110), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n752), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n748), .B(KEYINPUT108), .Z(new_n760));
  AOI21_X1  g559(.A(KEYINPUT109), .B1(new_n741), .B2(new_n742), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(new_n753), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT111), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n757), .A3(new_n753), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n754), .B2(new_n755), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n683), .A2(new_n659), .A3(new_n443), .A4(new_n736), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(new_n760), .B1(new_n772), .B2(new_n625), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n767), .B(new_n768), .C1(new_n773), .C2(new_n759), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n766), .A2(new_n774), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n737), .B2(new_n442), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n659), .A2(new_n420), .A3(new_n430), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT112), .Z(new_n778));
  NAND2_X1  g577(.A1(new_n743), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1338gat));
  OR2_X1    g579(.A1(new_n623), .A2(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n623), .A2(KEYINPUT113), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n781), .B(new_n782), .C1(new_n737), .C2(new_n449), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n449), .A2(G106gat), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n783), .B(new_n784), .C1(new_n744), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n659), .A3(new_n785), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n783), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n789), .B2(new_n784), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n453), .A2(new_n662), .A3(new_n444), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n594), .A2(new_n585), .B1(new_n597), .B2(new_n598), .ZN(new_n792));
  INV_X1    g591(.A(new_n608), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n612), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n636), .A2(new_n637), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n639), .B1(new_n796), .B2(new_n620), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n632), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n621), .A2(new_n630), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n644), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT114), .A4(new_n644), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n643), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n644), .B1(new_n798), .B2(new_n799), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n650), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n658), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n581), .A2(new_n795), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n613), .A2(new_n813), .B1(new_n659), .B2(new_n795), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n581), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n507), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n582), .A2(new_n614), .A3(new_n747), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n791), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n613), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n659), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n506), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g624(.A1(new_n819), .A2(new_n581), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n263), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT56), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(G134gat), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n817), .A2(new_n818), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n257), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n674), .A2(new_n690), .A3(new_n443), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(G141gat), .A3(new_n614), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT58), .B1(new_n837), .B2(KEYINPUT119), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n257), .A2(KEYINPUT57), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n812), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n810), .A2(KEYINPUT116), .A3(new_n658), .A4(new_n811), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n613), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n659), .A2(new_n795), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n680), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n506), .B1(new_n846), .B2(new_n814), .ZN(new_n847));
  NOR4_X1   g646(.A1(new_n507), .A2(new_n581), .A3(new_n613), .A4(new_n659), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n839), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT117), .ZN(new_n850));
  XOR2_X1   g649(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n851));
  NAND2_X1  g650(.A1(new_n832), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n839), .C1(new_n847), .C2(new_n848), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n613), .A3(new_n833), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n838), .B(new_n857), .C1(KEYINPUT119), .C2(new_n837), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n856), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT118), .B1(new_n856), .B2(G141gat), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n837), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(G1344gat));
  INV_X1    g662(.A(G148gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n835), .A2(new_n864), .A3(new_n659), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT120), .B1(new_n680), .B2(new_n812), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n581), .A2(new_n868), .A3(new_n813), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n867), .A2(new_n795), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n846), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n507), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n818), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n257), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n832), .A2(new_n851), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n659), .A3(new_n833), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n866), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n855), .A2(new_n833), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n864), .C1(new_n879), .C2(new_n659), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n865), .B1(new_n878), .B2(new_n880), .ZN(G1345gat));
  AOI21_X1  g680(.A(G155gat), .B1(new_n835), .B2(new_n506), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n879), .A2(G155gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n506), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n835), .B2(new_n581), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n879), .A2(new_n581), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n444), .A2(new_n662), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n430), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n257), .B1(new_n889), .B2(KEYINPUT121), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n831), .B(new_n890), .C1(KEYINPUT121), .C2(new_n889), .ZN(new_n891));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n614), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n662), .B1(new_n817), .B2(new_n818), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n450), .A2(new_n444), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(G169gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n892), .B1(new_n896), .B2(new_n614), .ZN(G1348gat));
  INV_X1    g696(.A(new_n895), .ZN(new_n898));
  AOI21_X1  g697(.A(G176gat), .B1(new_n898), .B2(new_n659), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n891), .A2(new_n648), .A3(new_n747), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1349gat));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n506), .A3(new_n324), .ZN(new_n902));
  OAI21_X1  g701(.A(G183gat), .B1(new_n891), .B2(new_n507), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT60), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n904), .B(new_n906), .Z(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n891), .B2(new_n680), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT61), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n325), .A3(new_n581), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1351gat));
  AND2_X1   g710(.A1(new_n442), .A2(new_n888), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n876), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n913), .B2(new_n614), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n876), .A2(new_n915), .A3(new_n613), .A4(new_n912), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(G197gat), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n442), .A2(new_n443), .A3(new_n257), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n893), .A3(new_n921), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n922), .A2(G197gat), .A3(new_n614), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n917), .A2(new_n923), .ZN(G1352gat));
  INV_X1    g723(.A(new_n922), .ZN(new_n925));
  INV_X1    g724(.A(G204gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n659), .ZN(new_n927));
  AND2_X1   g726(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n928));
  NOR2_X1   g727(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n876), .A2(new_n659), .A3(new_n912), .ZN(new_n931));
  OAI221_X1 g730(.A(new_n930), .B1(new_n928), .B2(new_n927), .C1(new_n931), .C2(new_n926), .ZN(G1353gat));
  OAI211_X1 g731(.A(new_n506), .B(new_n912), .C1(new_n874), .C2(new_n875), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G211gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(KEYINPUT126), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n925), .A2(new_n208), .A3(new_n506), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n940), .A3(new_n935), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n913), .B2(new_n680), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n209), .A3(new_n581), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


