//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n214), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  AND2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT67), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(new_n215), .A3(KEYINPUT8), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n207), .A2(G33), .ZN(new_n255));
  OR2_X1    g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n249), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n249), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n206), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G50), .B2(new_n261), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n276), .A2(G223), .B1(G77), .B2(new_n274), .ZN(new_n277));
  INV_X1    g0077(.A(G222), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n213), .A2(KEYINPUT66), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT66), .B1(new_n213), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n213), .B2(new_n282), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n290), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n292), .B1(G226), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n286), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n268), .A2(new_n269), .B1(new_n297), .B2(G190), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n286), .A2(new_n296), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n267), .A2(KEYINPUT9), .B1(new_n299), .B2(G200), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(new_n303), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n268), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT68), .ZN(new_n311));
  INV_X1    g0111(.A(new_n285), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n279), .A2(G232), .A3(new_n275), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n274), .A2(G107), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n279), .A2(G1698), .ZN(new_n315));
  INV_X1    g0115(.A(G238), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n318), .B2(new_n317), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n295), .A2(G244), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n291), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(G169), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n207), .A2(new_n270), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n250), .A2(new_n326), .B1(new_n207), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n255), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n260), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n249), .A2(new_n261), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n264), .A2(G77), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n331), .B1(G77), .B2(new_n261), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n324), .A2(new_n325), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n325), .B1(new_n324), .B2(new_n335), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n320), .A2(new_n306), .A3(new_n323), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n320), .A2(new_n323), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n335), .C1(new_n342), .C2(new_n340), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n305), .A2(new_n311), .A3(new_n339), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  INV_X1    g0146(.A(G226), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n346), .C1(new_n280), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n285), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n292), .B1(G238), .B2(new_n295), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n349), .A2(new_n350), .A3(new_n352), .A4(KEYINPUT13), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(G200), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n349), .A2(new_n350), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n349), .B2(new_n350), .ZN(new_n361));
  OAI21_X1  g0161(.A(G190), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n262), .A2(new_n216), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT12), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n326), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n255), .A2(new_n327), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n260), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n364), .B(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n357), .A2(new_n362), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n357), .A2(new_n362), .A3(KEYINPUT73), .A4(new_n372), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n355), .A2(G169), .A3(new_n356), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n384));
  OAI21_X1  g0184(.A(G179), .B1(new_n360), .B2(new_n361), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n371), .B2(new_n370), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n251), .A2(new_n253), .A3(new_n264), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n251), .A2(KEYINPUT77), .A3(new_n253), .A4(new_n264), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n263), .ZN(new_n394));
  INV_X1    g0194(.A(new_n254), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n392), .A2(new_n394), .B1(new_n261), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n279), .B2(G20), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n272), .A2(G33), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT7), .B(new_n207), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(KEYINPUT76), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT76), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n397), .C1(new_n279), .C2(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(G68), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n207), .B1(new_n217), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G159), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n326), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n398), .A2(new_n401), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n407), .B2(new_n409), .ZN(new_n416));
  INV_X1    g0216(.A(new_n406), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n417), .B2(new_n201), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n257), .A2(G159), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(KEYINPUT75), .A3(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n414), .A2(G68), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n249), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n396), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(G1698), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n271), .A2(new_n273), .A3(G223), .A4(new_n275), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n285), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n293), .A2(G232), .A3(new_n289), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n291), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n430), .A3(new_n342), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n291), .A2(new_n429), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n285), .B2(new_n427), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n431), .B1(new_n433), .B2(G200), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n423), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n394), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n391), .B1(new_n262), .B2(new_n254), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT7), .B1(new_n274), .B2(new_n207), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n397), .B(G20), .C1(new_n271), .C2(new_n273), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n416), .A2(new_n420), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n260), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT16), .B1(new_n405), .B2(new_n410), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n437), .B(new_n434), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT79), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n413), .A2(new_n422), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n437), .A4(new_n434), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n435), .B1(new_n450), .B2(KEYINPUT17), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n428), .A2(new_n430), .A3(new_n306), .ZN(new_n452));
  AOI21_X1  g0252(.A(G169), .B1(new_n428), .B2(new_n430), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT78), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n428), .A2(new_n430), .A3(new_n306), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT78), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n455), .B(new_n456), .C1(new_n433), .C2(G169), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT18), .B1(new_n423), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n437), .B1(new_n443), .B2(new_n444), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n454), .A4(new_n457), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n451), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NOR4_X1   g0263(.A1(new_n344), .A2(new_n381), .A3(new_n388), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n261), .A2(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT25), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G33), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n249), .A2(new_n467), .A3(new_n261), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n261), .A2(new_n468), .A3(new_n248), .A4(new_n247), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G107), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n279), .A2(KEYINPUT86), .A3(new_n207), .A4(G87), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT22), .ZN(new_n476));
  OR2_X1    g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n476), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G116), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n207), .B2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(KEYINPUT23), .A3(G20), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT24), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n477), .A2(new_n487), .A3(new_n478), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n474), .B1(new_n489), .B2(new_n260), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n275), .A2(G257), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G250), .B2(G1698), .ZN(new_n492));
  INV_X1    g0292(.A(G294), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n492), .A2(new_n274), .B1(new_n270), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n285), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT82), .B1(new_n496), .B2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  INV_X1    g0298(.A(G41), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n206), .A2(G45), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n504), .A3(new_n288), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n294), .B1(new_n501), .B2(new_n504), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n506), .A2(new_n507), .A3(G264), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n506), .B2(G264), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n495), .B(new_n505), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n510), .A2(KEYINPUT88), .A3(new_n306), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT88), .B1(new_n510), .B2(new_n306), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(G264), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n495), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G169), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n490), .B1(new_n516), .B2(KEYINPUT89), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT89), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n511), .A2(new_n518), .A3(new_n512), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G200), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n510), .A2(KEYINPUT90), .A3(new_n521), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n514), .A2(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT90), .B1(new_n510), .B2(new_n521), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n490), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n528), .B(KEYINPUT81), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(new_n275), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n285), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n506), .A2(G257), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n505), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n308), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n535), .A2(new_n306), .A3(new_n505), .A4(new_n536), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n402), .A2(G107), .A3(new_n404), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n473), .A2(KEYINPUT6), .A3(G97), .ZN(new_n541));
  XOR2_X1   g0341(.A(G97), .B(G107), .Z(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(KEYINPUT6), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n249), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n469), .A2(new_n471), .A3(G97), .ZN(new_n546));
  INV_X1    g0346(.A(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n262), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n538), .B(new_n539), .C1(new_n545), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n537), .A2(G200), .ZN(new_n551));
  INV_X1    g0351(.A(new_n545), .ZN(new_n552));
  INV_X1    g0352(.A(new_n549), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n535), .A2(G190), .A3(new_n505), .A4(new_n536), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n207), .B1(new_n346), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n547), .A3(new_n473), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n271), .A2(new_n273), .A3(new_n207), .A4(G68), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n557), .B1(new_n255), .B2(new_n547), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n260), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n329), .A2(new_n262), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n472), .C2(new_n329), .ZN(new_n567));
  INV_X1    g0367(.A(G45), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G1), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n293), .A2(G274), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n293), .A2(G250), .A3(new_n503), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n271), .A2(new_n273), .A3(G238), .A4(new_n275), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n479), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n285), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n306), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n567), .B(new_n577), .C1(G169), .C2(new_n576), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT83), .B1(new_n472), .B2(new_n559), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT83), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n469), .A2(new_n471), .A3(new_n580), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n565), .A2(new_n566), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n576), .A2(G190), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n521), .B2(new_n576), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n578), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n556), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n506), .A2(G270), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n591), .A2(new_n505), .ZN(new_n592));
  INV_X1    g0392(.A(G264), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n315), .A2(new_n593), .B1(new_n594), .B2(new_n279), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n279), .A2(new_n596), .A3(G257), .A4(new_n275), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n279), .A2(G257), .A3(new_n275), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT84), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n592), .B(G179), .C1(new_n600), .C2(new_n312), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n470), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n262), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n249), .B1(G20), .B2(new_n602), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(new_n270), .B2(G97), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n529), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n608), .A3(KEYINPUT20), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT85), .B1(new_n601), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n613), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n591), .A2(new_n505), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n599), .A2(new_n597), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n276), .A2(G264), .B1(G303), .B2(new_n274), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n285), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n615), .A2(new_n616), .A3(new_n621), .A4(G179), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n613), .A2(new_n308), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n592), .B1(new_n600), .B2(new_n312), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(G190), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n629), .B(new_n613), .C1(new_n521), .C2(new_n621), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(KEYINPUT21), .A3(new_n625), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n623), .A2(new_n628), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n590), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n464), .A2(new_n527), .A3(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n311), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n339), .B1(new_n375), .B2(new_n377), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n451), .B1(new_n636), .B2(new_n388), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n459), .A2(KEYINPUT94), .A3(new_n462), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT94), .B1(new_n459), .B2(new_n462), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n635), .B1(new_n640), .B2(new_n305), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT91), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n575), .A2(new_n285), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n642), .B(G200), .C1(new_n643), .C2(new_n572), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT91), .B1(new_n576), .B2(new_n521), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n586), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n578), .B1(new_n646), .B2(new_n585), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT92), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n578), .B(new_n649), .C1(new_n646), .C2(new_n585), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n550), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT93), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(new_n550), .ZN(new_n653));
  INV_X1    g0453(.A(new_n650), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n583), .B1(new_n579), .B2(new_n581), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(new_n586), .A3(new_n644), .A4(new_n645), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n656), .B2(new_n578), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT93), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n550), .A2(new_n588), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT26), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n652), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n578), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n556), .A2(new_n526), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n654), .A2(new_n657), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n490), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n516), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n623), .A3(new_n628), .A4(new_n631), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n665), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n464), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n641), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n490), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT95), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n527), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n517), .A2(new_n519), .A3(new_n681), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n623), .A2(new_n628), .A3(new_n631), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n613), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n632), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n682), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n527), .A2(new_n684), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n516), .A2(new_n669), .A3(new_n682), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT96), .ZN(G399));
  INV_X1    g0502(.A(new_n210), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n560), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n218), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n673), .A2(new_n682), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT98), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT98), .B(new_n660), .C1(new_n550), .C2(new_n588), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n714), .B(new_n715), .C1(new_n658), .C2(new_n660), .ZN(new_n716));
  INV_X1    g0516(.A(new_n668), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n688), .B1(new_n517), .B2(new_n519), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n716), .B(new_n578), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n712), .B1(new_n719), .B2(new_n682), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n621), .A2(G179), .A3(new_n576), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n510), .A3(new_n537), .ZN(new_n723));
  INV_X1    g0523(.A(new_n601), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n508), .A2(new_n509), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n285), .B2(new_n494), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n535), .A2(new_n536), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n724), .A2(new_n726), .A3(new_n727), .A4(new_n576), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT97), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n728), .B2(new_n729), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n728), .A2(new_n729), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n731), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n682), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n633), .A2(new_n520), .A3(new_n526), .A4(new_n682), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(KEYINPUT31), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n734), .A2(new_n730), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n739), .A2(new_n740), .A3(new_n682), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n721), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n709), .B1(new_n745), .B2(G1), .ZN(G364));
  INV_X1    g0546(.A(G13), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n206), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n704), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n693), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n691), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n248), .B1(G20), .B2(new_n308), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n207), .A2(new_n306), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n342), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n207), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n342), .A3(G200), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n202), .B1(new_n761), .B2(new_n473), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n757), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n342), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n207), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n216), .B1(new_n547), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n756), .A2(G190), .A3(new_n521), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n279), .B1(new_n769), .B2(new_n327), .C1(new_n215), .C2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n762), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(new_n768), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G159), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(KEYINPUT32), .B1(new_n777), .B2(G87), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n772), .B(new_n778), .C1(KEYINPUT32), .C2(new_n775), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n274), .B1(new_n769), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n781), .B(new_n783), .C1(G329), .C2(new_n774), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n758), .A2(G326), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n763), .A2(new_n786), .B1(new_n777), .B2(G303), .ZN(new_n787));
  INV_X1    g0587(.A(new_n766), .ZN(new_n788));
  INV_X1    g0588(.A(new_n761), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n788), .A2(G294), .B1(new_n789), .B2(G283), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n755), .B1(new_n779), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n703), .A2(new_n274), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G355), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G116), .B2(new_n210), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n703), .A2(new_n279), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n218), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n568), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n242), .A2(new_n568), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n754), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n751), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n792), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n804), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n691), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n753), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n335), .A2(new_n682), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n339), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(new_n339), .B2(new_n343), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n710), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n681), .B1(new_n664), .B2(new_n672), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n814), .A2(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n751), .B1(new_n743), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n743), .B2(new_n821), .ZN(new_n823));
  INV_X1    g0623(.A(new_n751), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n754), .A2(new_n802), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n327), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n769), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n763), .A2(G283), .B1(new_n827), .B2(G116), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT100), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n766), .A2(new_n547), .B1(new_n770), .B2(new_n493), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n828), .A2(new_n829), .B1(KEYINPUT101), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT101), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n828), .A2(new_n829), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n274), .B1(new_n773), .B2(new_n782), .C1(new_n559), .C2(new_n761), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n759), .A2(new_n594), .B1(new_n776), .B2(new_n473), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n279), .B1(new_n773), .B2(new_n837), .C1(new_n202), .C2(new_n776), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n766), .A2(new_n215), .B1(new_n761), .B2(new_n216), .ZN(new_n839));
  INV_X1    g0639(.A(new_n770), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(G143), .B1(new_n827), .B2(G159), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G137), .A2(new_n758), .B1(new_n763), .B2(G150), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT34), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n838), .B(new_n839), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n836), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n826), .B1(new_n755), .B2(new_n850), .C1(new_n819), .C2(new_n803), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n823), .A2(new_n851), .ZN(G384));
  NAND2_X1  g0652(.A1(new_n406), .A2(G77), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n218), .A2(new_n853), .B1(G50), .B2(new_n216), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(G1), .A3(new_n747), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT103), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n602), .B(new_n214), .C1(new_n543), .C2(KEYINPUT35), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(KEYINPUT35), .B2(new_n543), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT36), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n638), .A2(new_n639), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n679), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n339), .A2(new_n681), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT104), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n818), .B2(new_n819), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n372), .A2(new_n682), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n375), .B2(new_n377), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n387), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n380), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n386), .B1(new_n872), .B2(new_n378), .ZN(new_n873));
  INV_X1    g0673(.A(new_n869), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n440), .A2(new_n441), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT105), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n421), .A2(KEYINPUT105), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n443), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT106), .B1(new_n882), .B2(new_n396), .ZN(new_n883));
  INV_X1    g0683(.A(new_n679), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n412), .B1(new_n421), .B2(KEYINPUT105), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n878), .A2(new_n879), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n422), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT106), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n437), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n877), .B1(new_n463), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n446), .A2(new_n449), .ZN(new_n893));
  INV_X1    g0693(.A(new_n458), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n883), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n460), .A2(new_n454), .A3(new_n457), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n460), .A2(new_n884), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n893), .A3(KEYINPUT108), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT108), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n450), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT107), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n892), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT109), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT109), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n892), .B(new_n911), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n463), .A2(new_n891), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n907), .B2(new_n908), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n910), .A2(new_n912), .B1(new_n877), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n863), .B1(new_n876), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT110), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n451), .B1(new_n638), .B2(new_n639), .ZN(new_n919));
  INV_X1    g0719(.A(new_n900), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n898), .A2(new_n445), .A3(new_n900), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT108), .B1(new_n901), .B2(new_n893), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n904), .A2(new_n450), .A3(new_n903), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT111), .B1(new_n927), .B2(new_n877), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT111), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n929), .B(KEYINPUT38), .C1(new_n921), .C2(new_n926), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n918), .B(new_n909), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n915), .B2(new_n918), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n387), .A2(new_n681), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT110), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n863), .C1(new_n876), .C2(new_n915), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n917), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n464), .B1(new_n711), .B2(new_n720), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n641), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n736), .A2(KEYINPUT31), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n875), .B(new_n819), .C1(new_n738), .C2(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n906), .A2(new_n923), .B1(new_n919), .B2(new_n920), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n929), .B1(new_n943), .B2(KEYINPUT38), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n927), .A2(KEYINPUT111), .A3(new_n877), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n946), .B2(new_n909), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n869), .B1(new_n381), .B2(new_n386), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n816), .B1(new_n949), .B2(new_n871), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n948), .C1(new_n738), .C2(new_n941), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n947), .A2(new_n948), .B1(new_n915), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n464), .B1(new_n738), .B2(new_n941), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(G330), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n206), .B2(new_n748), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n940), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n861), .B1(new_n959), .B2(new_n960), .ZN(G367));
  INV_X1    g0761(.A(KEYINPUT113), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n653), .A2(new_n681), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT112), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n681), .B1(new_n545), .B2(new_n549), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n556), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n698), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n550), .B1(new_n968), .B2(new_n520), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n969), .A2(KEYINPUT42), .B1(new_n682), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n585), .A2(new_n681), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n578), .ZN(new_n975));
  INV_X1    g0775(.A(new_n667), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n970), .A2(new_n972), .A3(new_n978), .A4(new_n977), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n694), .A2(new_n968), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n962), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n986), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n982), .A2(KEYINPUT113), .A3(new_n985), .A4(new_n983), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n704), .B(KEYINPUT41), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n700), .A2(new_n968), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n698), .A2(new_n699), .A3(new_n967), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n695), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n698), .B1(new_n687), .B2(new_n697), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(new_n692), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n994), .A2(new_n997), .A3(new_n694), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n999), .A2(new_n745), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n991), .B1(new_n1004), .B2(new_n745), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n990), .B1(new_n750), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n234), .A2(new_n797), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n805), .B1(new_n210), .B2(new_n329), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n751), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n764), .A2(new_n408), .B1(new_n776), .B2(new_n215), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G68), .B2(new_n788), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n274), .B1(new_n827), .B2(G50), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(KEYINPUT114), .B(G137), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n840), .A2(G150), .B1(new_n774), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n761), .A2(new_n327), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G143), .B2(new_n758), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n776), .A2(new_n602), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT46), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G107), .A2(new_n788), .B1(new_n758), .B2(G311), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n279), .B1(new_n840), .B2(G303), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G283), .A2(new_n827), .B1(new_n774), .B2(G317), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n763), .A2(G294), .B1(new_n789), .B2(G97), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1018), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1009), .B1(new_n1027), .B2(new_n754), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n980), .B2(new_n809), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1006), .A2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n1002), .A2(new_n750), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n706), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n793), .A2(new_n1032), .B1(new_n473), .B2(new_n703), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n238), .A2(new_n568), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n250), .A2(G50), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT50), .Z(new_n1036));
  OAI211_X1 g0836(.A(new_n706), .B(new_n568), .C1(new_n216), .C2(new_n327), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n796), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n824), .B1(new_n1039), .B2(new_n805), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G68), .A2(new_n827), .B1(new_n774), .B2(G150), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n274), .B1(new_n840), .B2(G50), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n254), .C2(new_n764), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n759), .A2(new_n408), .B1(new_n776), .B2(new_n327), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n761), .A2(new_n547), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n766), .A2(new_n329), .ZN(new_n1046));
  NOR4_X1   g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n840), .A2(G317), .B1(new_n827), .B2(G303), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n759), .B2(new_n780), .C1(new_n782), .C2(new_n764), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n788), .A2(G283), .B1(new_n777), .B2(G294), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT116), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n279), .B1(new_n774), .B2(G326), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n602), .B2(new_n761), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1056), .B2(KEYINPUT116), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1047), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1040), .B1(new_n755), .B2(new_n1061), .C1(new_n687), .C2(new_n809), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1031), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1002), .A2(new_n745), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1001), .B1(new_n744), .B2(new_n721), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n704), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n999), .A2(new_n1003), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n1064), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n1004), .A3(new_n704), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n999), .A2(new_n750), .A3(new_n1003), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G317), .A2(new_n758), .B1(new_n840), .B2(G311), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n274), .B1(new_n773), .B2(new_n780), .C1(new_n493), .C2(new_n769), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n764), .A2(new_n594), .B1(new_n761), .B2(new_n473), .ZN(new_n1075));
  INV_X1    g0875(.A(G283), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n766), .A2(new_n602), .B1(new_n776), .B2(new_n1076), .ZN(new_n1077));
  OR4_X1    g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(G150), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n759), .A2(new_n1079), .B1(new_n408), .B2(new_n770), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  INV_X1    g0881(.A(G143), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n279), .B1(new_n773), .B2(new_n1082), .C1(new_n250), .C2(new_n769), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n766), .A2(new_n327), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G87), .B2(new_n789), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n763), .A2(G50), .B1(new_n777), .B2(G68), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1081), .A2(new_n1084), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n755), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n797), .A2(new_n245), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n806), .B1(G97), .B2(new_n703), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n824), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n967), .B2(new_n809), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1071), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1070), .A2(new_n1094), .ZN(G390));
  INV_X1    g0895(.A(new_n933), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n875), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n867), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n931), .B(new_n1098), .C1(new_n915), .C2(new_n918), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n909), .B1(new_n928), .B2(new_n930), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n719), .A2(new_n682), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n864), .B1(new_n1101), .B2(new_n819), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1100), .B(new_n1096), .C1(new_n1102), .C2(new_n1097), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(G330), .B1(new_n738), .B2(new_n941), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n875), .A2(new_n819), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(G330), .B(new_n819), .C1(new_n738), .C2(new_n741), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(new_n1097), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1099), .A2(new_n1103), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1112), .A2(new_n749), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n932), .A2(new_n803), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n825), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n751), .B1(new_n395), .B2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n758), .A2(G283), .B1(new_n827), .B2(G97), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n473), .B2(new_n764), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT119), .Z(new_n1119));
  OAI221_X1 g0919(.A(new_n274), .B1(new_n773), .B2(new_n493), .C1(new_n770), .C2(new_n602), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n216), .A2(new_n761), .B1(new_n776), .B2(new_n559), .ZN(new_n1121));
  OR3_X1    g0921(.A1(new_n1120), .A2(new_n1085), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT118), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n776), .A2(new_n1079), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT53), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n770), .A2(new_n837), .B1(new_n773), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n279), .B1(new_n769), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n758), .A2(G128), .B1(new_n789), .B2(G50), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G159), .A2(new_n788), .B1(new_n763), .B2(new_n1014), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1126), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1123), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1116), .B1(new_n1136), .B2(new_n754), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1113), .B1(new_n1114), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1109), .A2(new_n1097), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n868), .B1(new_n1140), .B2(new_n1107), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1097), .B1(new_n1105), .B2(new_n816), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1110), .A2(new_n1102), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n464), .B(G330), .C1(new_n738), .C2(new_n941), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n938), .A2(new_n641), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n705), .B1(new_n1112), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1108), .A2(new_n1111), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1139), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1111), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1107), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1148), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AND4_X1   g0956(.A1(new_n1139), .A2(new_n1156), .A3(new_n704), .A4(new_n1151), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1138), .B1(new_n1152), .B2(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(new_n942), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n948), .B1(new_n1100), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n915), .A2(new_n951), .ZN(new_n1161));
  OAI21_X1  g0961(.A(G330), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n305), .A2(new_n310), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n268), .A2(new_n884), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1165), .B(new_n1166), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n914), .A2(new_n877), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n912), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT107), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n906), .A3(new_n897), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n911), .B1(new_n1174), .B2(new_n892), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1169), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n867), .A2(new_n1097), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1176), .A2(new_n1177), .B1(new_n862), .B2(new_n679), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n935), .A2(new_n1178), .B1(new_n932), .B2(new_n933), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1167), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n952), .A2(G330), .A3(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1168), .A2(new_n917), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G330), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n944), .A2(new_n945), .B1(new_n1174), .B2(new_n892), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT40), .B1(new_n1184), .B2(new_n942), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n942), .A2(KEYINPUT40), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1183), .B(new_n1167), .C1(new_n1185), .C2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1180), .B1(new_n952), .B2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n937), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1182), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n750), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1180), .A2(new_n803), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n751), .B1(G50), .B2(new_n1115), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n274), .B2(new_n499), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n759), .A2(new_n602), .B1(new_n761), .B2(new_n215), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G97), .B2(new_n763), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G41), .B(new_n279), .C1(new_n774), .C2(G283), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n769), .A2(new_n329), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G107), .B2(new_n840), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n788), .A2(G68), .B1(new_n777), .B2(G77), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT58), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1206));
  INV_X1    g1006(.A(G128), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n770), .A2(new_n1207), .B1(new_n776), .B2(new_n1129), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT120), .Z(new_n1209));
  AOI22_X1  g1009(.A1(new_n758), .A2(G125), .B1(new_n827), .B2(G137), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G150), .A2(new_n788), .B1(new_n763), .B2(G132), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1206), .B1(new_n408), .B2(new_n761), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1205), .B1(new_n1204), .B2(new_n1203), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1194), .B1(new_n1216), .B2(new_n754), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1193), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1192), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1151), .A2(new_n1147), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n937), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1168), .A2(new_n1181), .B1(new_n1179), .B2(new_n917), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n705), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1182), .A2(new_n1190), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1228), .A2(KEYINPUT121), .A3(new_n917), .A4(new_n1179), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1224), .B1(new_n1151), .B2(new_n1147), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1219), .B1(new_n1225), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(G375));
  NAND3_X1  g1033(.A1(new_n1141), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n991), .B(KEYINPUT122), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1148), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1097), .A2(new_n802), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G116), .A2(new_n763), .B1(new_n758), .B2(G294), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n547), .B2(new_n776), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n279), .B1(new_n774), .B2(G303), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n473), .B2(new_n769), .C1(new_n1076), .C2(new_n770), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1240), .A2(new_n1242), .A3(new_n1016), .A4(new_n1046), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n788), .A2(G50), .B1(new_n777), .B2(G159), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n837), .B2(new_n759), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n764), .A2(new_n1129), .B1(new_n761), .B2(new_n215), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n279), .B1(new_n773), .B2(new_n1207), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n770), .A2(new_n1013), .B1(new_n769), .B2(new_n1079), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n754), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n751), .C1(G68), .C2(new_n1115), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1238), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1144), .B2(new_n750), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1236), .A2(new_n1253), .ZN(G381));
  XOR2_X1   g1054(.A(new_n1232), .B(KEYINPUT123), .Z(new_n1255));
  NAND2_X1  g1055(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1138), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OR3_X1    g1060(.A1(new_n1260), .A2(G390), .A3(G384), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1261), .A2(G387), .A3(G381), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1255), .A2(new_n1258), .A3(new_n1262), .ZN(G407));
  NAND2_X1  g1063(.A1(new_n680), .A2(G213), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT124), .Z(new_n1265));
  NAND3_X1  g1065(.A1(new_n1255), .A2(new_n1258), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(G407), .A2(new_n1266), .A3(G213), .ZN(G409));
  NAND2_X1  g1067(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n704), .A3(new_n1231), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1219), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(G378), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1227), .A2(new_n750), .A3(new_n1229), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1191), .A2(new_n1220), .A3(new_n1235), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1218), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1258), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1150), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1234), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n704), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(new_n1234), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1253), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G384), .B(KEYINPUT125), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1253), .B(new_n1286), .C1(new_n1280), .C2(new_n1282), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1276), .A2(new_n1264), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n811), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1260), .A2(G390), .A3(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1070), .B(new_n1094), .C1(new_n1259), .C2(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G387), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1295), .A2(new_n1296), .A3(new_n1006), .A4(new_n1029), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1265), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1289), .A2(KEYINPUT63), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1301), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1264), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1265), .A2(G2897), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1287), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1307), .A2(G2897), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1289), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1306), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1310), .A2(new_n1287), .A3(new_n1312), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1289), .B2(new_n1309), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1232), .A2(G378), .B1(new_n1258), .B2(new_n1274), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1316), .B(KEYINPUT126), .C1(new_n1317), .C2(new_n1307), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1292), .A2(new_n1305), .A3(new_n1314), .A4(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1299), .B1(new_n1302), .B2(new_n1313), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1290), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1302), .A2(KEYINPUT62), .A3(new_n1289), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1320), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1319), .B1(new_n1324), .B2(new_n1325), .ZN(G405));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1269), .A2(G378), .A3(new_n1270), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1257), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1327), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1271), .B(KEYINPUT127), .C1(new_n1232), .C2(new_n1257), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1289), .A3(new_n1331), .ZN(new_n1332));
  OAI221_X1 g1132(.A(new_n1327), .B1(new_n1288), .B2(new_n1285), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1332), .A2(new_n1325), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1325), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(G402));
endmodule


