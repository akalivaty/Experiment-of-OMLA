

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733;

  INV_X1 U365 ( .A(n654), .ZN(n343) );
  INV_X1 U366 ( .A(n654), .ZN(n347) );
  BUF_X1 U367 ( .A(G119), .Z(n350) );
  XNOR2_X1 U368 ( .A(n377), .B(n472), .ZN(n610) );
  INV_X1 U369 ( .A(n342), .ZN(n599) );
  NAND2_X1 U370 ( .A1(n344), .A2(n343), .ZN(n342) );
  XNOR2_X1 U371 ( .A(n595), .B(n345), .ZN(n344) );
  INV_X1 U372 ( .A(n594), .ZN(n345) );
  INV_X1 U373 ( .A(n346), .ZN(n649) );
  NAND2_X1 U374 ( .A1(n348), .A2(n347), .ZN(n346) );
  XNOR2_X1 U375 ( .A(n647), .B(n349), .ZN(n348) );
  INV_X1 U376 ( .A(n646), .ZN(n349) );
  NAND2_X1 U377 ( .A1(n351), .A2(G210), .ZN(n653) );
  AND2_X2 U378 ( .A1(n360), .A2(n361), .ZN(n351) );
  XNOR2_X2 U379 ( .A(n610), .B(n384), .ZN(n650) );
  INV_X1 U380 ( .A(n567), .ZN(n545) );
  INV_X2 U381 ( .A(G953), .ZN(n727) );
  XNOR2_X2 U382 ( .A(n500), .B(n499), .ZN(n606) );
  AND2_X2 U383 ( .A1(n517), .A2(n516), .ZN(n525) );
  NAND2_X2 U384 ( .A1(n525), .A2(n524), .ZN(n527) );
  NAND2_X2 U385 ( .A1(n501), .A2(n435), .ZN(n437) );
  OR2_X1 U386 ( .A1(n493), .A2(n564), .ZN(n494) );
  XNOR2_X1 U387 ( .A(n558), .B(n392), .ZN(n570) );
  NAND2_X1 U388 ( .A1(n659), .A2(n484), .ZN(n486) );
  NOR2_X1 U389 ( .A1(n631), .A2(G902), .ZN(n465) );
  NOR2_X1 U390 ( .A1(n571), .A2(n690), .ZN(n551) );
  NOR2_X1 U391 ( .A1(n557), .A2(n543), .ZN(n544) );
  NOR2_X1 U392 ( .A1(n570), .A2(n396), .ZN(n362) );
  XNOR2_X1 U393 ( .A(n486), .B(n485), .ZN(n502) );
  XNOR2_X1 U394 ( .A(n476), .B(n475), .ZN(n567) );
  XNOR2_X1 U395 ( .A(KEYINPUT3), .B(G119), .ZN(n371) );
  OR2_X1 U396 ( .A1(n510), .A2(n672), .ZN(n515) );
  NAND2_X1 U397 ( .A1(n356), .A2(n363), .ZN(n609) );
  AND2_X1 U398 ( .A1(n365), .A2(n542), .ZN(n364) );
  XNOR2_X1 U399 ( .A(n362), .B(n397), .ZN(n498) );
  XNOR2_X2 U400 ( .A(n545), .B(KEYINPUT1), .ZN(n664) );
  XNOR2_X2 U401 ( .A(n596), .B(KEYINPUT86), .ZN(n654) );
  XNOR2_X1 U402 ( .A(n422), .B(KEYINPUT4), .ZN(n439) );
  XNOR2_X1 U403 ( .A(n378), .B(G128), .ZN(n422) );
  XNOR2_X1 U404 ( .A(n372), .B(n371), .ZN(n446) );
  XNOR2_X1 U405 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n373) );
  XNOR2_X1 U406 ( .A(G116), .B(G113), .ZN(n372) );
  XNOR2_X1 U407 ( .A(G146), .B(G125), .ZN(n405) );
  XNOR2_X1 U408 ( .A(G143), .B(KEYINPUT77), .ZN(n378) );
  NAND2_X1 U409 ( .A1(n361), .A2(n360), .ZN(n352) );
  NOR2_X2 U410 ( .A1(n591), .A2(n429), .ZN(n361) );
  INV_X1 U411 ( .A(n582), .ZN(n353) );
  INV_X1 U412 ( .A(n490), .ZN(n354) );
  AND2_X2 U413 ( .A1(n628), .A2(n521), .ZN(n482) );
  NAND2_X1 U414 ( .A1(n389), .A2(n674), .ZN(n390) );
  INV_X1 U415 ( .A(KEYINPUT38), .ZN(n370) );
  XNOR2_X1 U416 ( .A(n439), .B(n438), .ZN(n469) );
  XNOR2_X1 U417 ( .A(n409), .B(n634), .ZN(n410) );
  XNOR2_X1 U418 ( .A(n421), .B(n420), .ZN(n450) );
  XNOR2_X1 U419 ( .A(n419), .B(KEYINPUT79), .ZN(n421) );
  XNOR2_X1 U420 ( .A(n428), .B(n623), .ZN(n508) );
  AND2_X1 U421 ( .A1(n506), .A2(n508), .ZN(n676) );
  XNOR2_X1 U422 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U423 ( .A(n469), .B(n468), .ZN(n722) );
  XNOR2_X1 U424 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n379) );
  XNOR2_X1 U425 ( .A(n536), .B(KEYINPUT39), .ZN(n586) );
  AND2_X1 U426 ( .A1(n535), .A2(n502), .ZN(n536) );
  INV_X1 U427 ( .A(KEYINPUT65), .ZN(n366) );
  NAND2_X1 U428 ( .A1(n481), .A2(n366), .ZN(n365) );
  OR2_X1 U429 ( .A1(n514), .A2(n368), .ZN(n367) );
  NAND2_X1 U430 ( .A1(n369), .A2(KEYINPUT65), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U432 ( .A(n406), .B(n720), .ZN(n407) );
  XOR2_X1 U433 ( .A(n386), .B(KEYINPUT78), .Z(n355) );
  AND2_X1 U434 ( .A1(n367), .A2(n364), .ZN(n356) );
  AND2_X1 U435 ( .A1(n723), .A2(KEYINPUT81), .ZN(n357) );
  XOR2_X1 U436 ( .A(n479), .B(KEYINPUT32), .Z(n358) );
  AND2_X1 U437 ( .A1(n360), .A2(n359), .ZN(n657) );
  INV_X1 U438 ( .A(n591), .ZN(n359) );
  XNOR2_X2 U439 ( .A(n590), .B(KEYINPUT2), .ZN(n360) );
  AND2_X1 U440 ( .A1(n357), .A2(n612), .ZN(n591) );
  XNOR2_X2 U441 ( .A(n527), .B(n526), .ZN(n612) );
  INV_X1 U442 ( .A(n498), .ZN(n501) );
  NAND2_X1 U443 ( .A1(n514), .A2(n366), .ZN(n363) );
  INV_X1 U444 ( .A(n481), .ZN(n369) );
  XNOR2_X2 U445 ( .A(n437), .B(n436), .ZN(n514) );
  INV_X1 U446 ( .A(n389), .ZN(n563) );
  XNOR2_X1 U447 ( .A(n389), .B(n370), .ZN(n675) );
  XNOR2_X2 U448 ( .A(n387), .B(n355), .ZN(n389) );
  BUF_X1 U449 ( .A(n628), .Z(n629) );
  INV_X1 U450 ( .A(KEYINPUT98), .ZN(n414) );
  INV_X1 U451 ( .A(n467), .ZN(n468) );
  XNOR2_X1 U452 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U453 ( .A(n408), .B(n407), .ZN(n636) );
  XNOR2_X1 U454 ( .A(n411), .B(n410), .ZN(n509) );
  INV_X1 U455 ( .A(KEYINPUT63), .ZN(n598) );
  XNOR2_X1 U456 ( .A(n373), .B(G122), .ZN(n374) );
  XNOR2_X1 U457 ( .A(n446), .B(n374), .ZN(n377) );
  XNOR2_X1 U458 ( .A(G104), .B(G101), .ZN(n376) );
  XNOR2_X1 U459 ( .A(G110), .B(G107), .ZN(n375) );
  XNOR2_X1 U460 ( .A(n376), .B(n375), .ZN(n472) );
  XNOR2_X1 U461 ( .A(n405), .B(n379), .ZN(n382) );
  NAND2_X1 U462 ( .A1(n727), .A2(G224), .ZN(n380) );
  XNOR2_X1 U463 ( .A(n380), .B(KEYINPUT87), .ZN(n381) );
  XNOR2_X1 U464 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U465 ( .A(n439), .B(n383), .ZN(n384) );
  XNOR2_X1 U466 ( .A(KEYINPUT15), .B(G902), .ZN(n429) );
  INV_X1 U467 ( .A(n429), .ZN(n592) );
  OR2_X2 U468 ( .A1(n650), .A2(n592), .ZN(n387) );
  INV_X1 U469 ( .A(G902), .ZN(n427) );
  INV_X1 U470 ( .A(G237), .ZN(n385) );
  NAND2_X1 U471 ( .A1(n427), .A2(n385), .ZN(n388) );
  NAND2_X1 U472 ( .A1(n388), .A2(G210), .ZN(n386) );
  NAND2_X1 U473 ( .A1(n388), .A2(G214), .ZN(n674) );
  XNOR2_X2 U474 ( .A(n390), .B(KEYINPUT85), .ZN(n558) );
  XNOR2_X1 U475 ( .A(KEYINPUT73), .B(KEYINPUT19), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n391), .B(KEYINPUT67), .ZN(n392) );
  NAND2_X1 U477 ( .A1(G237), .A2(G234), .ZN(n393) );
  XNOR2_X1 U478 ( .A(n393), .B(KEYINPUT14), .ZN(n687) );
  NOR2_X1 U479 ( .A1(G898), .A2(n727), .ZN(n611) );
  NAND2_X1 U480 ( .A1(n611), .A2(G902), .ZN(n394) );
  NAND2_X1 U481 ( .A1(G952), .A2(n727), .ZN(n529) );
  NAND2_X1 U482 ( .A1(n394), .A2(n529), .ZN(n395) );
  NAND2_X1 U483 ( .A1(n687), .A2(n395), .ZN(n396) );
  INV_X1 U484 ( .A(KEYINPUT0), .ZN(n397) );
  NOR2_X1 U485 ( .A1(G953), .A2(G237), .ZN(n442) );
  NAND2_X1 U486 ( .A1(n442), .A2(G214), .ZN(n399) );
  XOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n398) );
  XNOR2_X1 U488 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U489 ( .A(n400), .B(KEYINPUT11), .Z(n408) );
  XOR2_X1 U490 ( .A(G113), .B(G104), .Z(n402) );
  XNOR2_X1 U491 ( .A(G122), .B(G131), .ZN(n401) );
  XNOR2_X1 U492 ( .A(n402), .B(n401), .ZN(n404) );
  XNOR2_X1 U493 ( .A(G143), .B(G140), .ZN(n403) );
  XNOR2_X1 U494 ( .A(n404), .B(n403), .ZN(n406) );
  XNOR2_X1 U495 ( .A(n405), .B(KEYINPUT10), .ZN(n720) );
  NOR2_X1 U496 ( .A1(G902), .A2(n636), .ZN(n411) );
  XNOR2_X1 U497 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n409) );
  INV_X1 U498 ( .A(G475), .ZN(n634) );
  INV_X1 U499 ( .A(n509), .ZN(n506) );
  XOR2_X1 U500 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n413) );
  XNOR2_X1 U501 ( .A(G116), .B(G122), .ZN(n412) );
  XNOR2_X1 U502 ( .A(n413), .B(n412), .ZN(n417) );
  XNOR2_X1 U503 ( .A(G134), .B(G107), .ZN(n415) );
  XOR2_X1 U504 ( .A(n418), .B(KEYINPUT9), .Z(n426) );
  NAND2_X1 U505 ( .A1(G234), .A2(n727), .ZN(n419) );
  XOR2_X1 U506 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n420) );
  NAND2_X1 U507 ( .A1(n450), .A2(G217), .ZN(n424) );
  XNOR2_X1 U508 ( .A(n422), .B(KEYINPUT7), .ZN(n423) );
  XNOR2_X1 U509 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n426), .B(n425), .ZN(n624) );
  NAND2_X1 U511 ( .A1(n624), .A2(n427), .ZN(n428) );
  INV_X1 U512 ( .A(G478), .ZN(n623) );
  XOR2_X1 U513 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n431) );
  NAND2_X1 U514 ( .A1(G234), .A2(n429), .ZN(n430) );
  XNOR2_X1 U515 ( .A(n431), .B(n430), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n460), .A2(G221), .ZN(n432) );
  XOR2_X1 U517 ( .A(KEYINPUT21), .B(n432), .Z(n434) );
  INV_X1 U518 ( .A(KEYINPUT91), .ZN(n433) );
  XNOR2_X1 U519 ( .A(n434), .B(n433), .ZN(n658) );
  XNOR2_X1 U520 ( .A(n658), .B(KEYINPUT92), .ZN(n484) );
  AND2_X1 U521 ( .A1(n676), .A2(n484), .ZN(n435) );
  XNOR2_X1 U522 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n436) );
  XNOR2_X1 U523 ( .A(G134), .B(G131), .ZN(n438) );
  XOR2_X1 U524 ( .A(KEYINPUT5), .B(G137), .Z(n441) );
  XNOR2_X1 U525 ( .A(G146), .B(G101), .ZN(n440) );
  XNOR2_X1 U526 ( .A(n441), .B(n440), .ZN(n444) );
  NAND2_X1 U527 ( .A1(G210), .A2(n442), .ZN(n443) );
  XNOR2_X1 U528 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U529 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U530 ( .A(n469), .B(n447), .ZN(n593) );
  OR2_X1 U531 ( .A1(n593), .A2(G902), .ZN(n448) );
  XNOR2_X2 U532 ( .A(n448), .B(G472), .ZN(n662) );
  INV_X1 U533 ( .A(KEYINPUT6), .ZN(n449) );
  XNOR2_X1 U534 ( .A(n662), .B(n449), .ZN(n555) );
  XNOR2_X1 U535 ( .A(n555), .B(KEYINPUT76), .ZN(n466) );
  NAND2_X1 U536 ( .A1(n450), .A2(G221), .ZN(n454) );
  XOR2_X1 U537 ( .A(KEYINPUT74), .B(KEYINPUT23), .Z(n452) );
  XNOR2_X1 U538 ( .A(G110), .B(KEYINPUT24), .ZN(n451) );
  XOR2_X1 U539 ( .A(n452), .B(n451), .Z(n453) );
  XNOR2_X1 U540 ( .A(n454), .B(n453), .ZN(n459) );
  XNOR2_X1 U541 ( .A(G128), .B(n720), .ZN(n457) );
  INV_X1 U542 ( .A(G140), .ZN(n455) );
  XNOR2_X1 U543 ( .A(n455), .B(G137), .ZN(n467) );
  XOR2_X1 U544 ( .A(n467), .B(n350), .Z(n456) );
  XNOR2_X1 U545 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U546 ( .A(n459), .B(n458), .ZN(n631) );
  NAND2_X1 U547 ( .A1(n460), .A2(G217), .ZN(n461) );
  XNOR2_X1 U548 ( .A(n461), .B(KEYINPUT90), .ZN(n463) );
  XNOR2_X1 U549 ( .A(KEYINPUT25), .B(KEYINPUT88), .ZN(n462) );
  XNOR2_X2 U550 ( .A(n465), .B(n464), .ZN(n659) );
  NOR2_X1 U551 ( .A1(n466), .A2(n659), .ZN(n477) );
  NAND2_X1 U552 ( .A1(n727), .A2(G227), .ZN(n470) );
  XNOR2_X1 U553 ( .A(n470), .B(G146), .ZN(n471) );
  XNOR2_X1 U554 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U555 ( .A(n722), .B(n473), .ZN(n645) );
  OR2_X1 U556 ( .A1(n645), .A2(G902), .ZN(n476) );
  INV_X1 U557 ( .A(KEYINPUT70), .ZN(n474) );
  XNOR2_X1 U558 ( .A(n474), .B(G469), .ZN(n475) );
  NAND2_X1 U559 ( .A1(n477), .A2(n353), .ZN(n478) );
  NOR2_X2 U560 ( .A1(n514), .A2(n478), .ZN(n480) );
  INV_X1 U561 ( .A(KEYINPUT75), .ZN(n479) );
  XNOR2_X2 U562 ( .A(n480), .B(n358), .ZN(n628) );
  INV_X1 U563 ( .A(KEYINPUT44), .ZN(n521) );
  OR2_X1 U564 ( .A1(n664), .A2(n662), .ZN(n481) );
  INV_X1 U565 ( .A(n659), .ZN(n542) );
  NAND2_X1 U566 ( .A1(n482), .A2(n609), .ZN(n483) );
  NAND2_X1 U567 ( .A1(n483), .A2(KEYINPUT84), .ZN(n496) );
  INV_X1 U568 ( .A(KEYINPUT68), .ZN(n485) );
  AND2_X1 U569 ( .A1(n502), .A2(n555), .ZN(n487) );
  NAND2_X1 U570 ( .A1(n487), .A2(n664), .ZN(n489) );
  XNOR2_X1 U571 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n488) );
  XNOR2_X2 U572 ( .A(n489), .B(n488), .ZN(n691) );
  BUF_X1 U573 ( .A(n498), .Z(n490) );
  NOR2_X1 U574 ( .A1(n691), .A2(n490), .ZN(n492) );
  INV_X1 U575 ( .A(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U576 ( .A(n492), .B(n491), .ZN(n493) );
  INV_X1 U577 ( .A(n508), .ZN(n507) );
  NAND2_X1 U578 ( .A1(n509), .A2(n507), .ZN(n564) );
  XNOR2_X2 U579 ( .A(n494), .B(KEYINPUT35), .ZN(n630) );
  INV_X1 U580 ( .A(n630), .ZN(n495) );
  NAND2_X1 U581 ( .A1(n496), .A2(n495), .ZN(n517) );
  AND2_X1 U582 ( .A1(n502), .A2(n662), .ZN(n497) );
  NAND2_X1 U583 ( .A1(n497), .A2(n664), .ZN(n668) );
  OR2_X1 U584 ( .A1(n668), .A2(n498), .ZN(n500) );
  INV_X1 U585 ( .A(KEYINPUT31), .ZN(n499) );
  INV_X1 U586 ( .A(n662), .ZN(n543) );
  AND2_X1 U587 ( .A1(n545), .A2(n543), .ZN(n503) );
  AND2_X1 U588 ( .A1(n502), .A2(n503), .ZN(n504) );
  NAND2_X1 U589 ( .A1(n354), .A2(n504), .ZN(n699) );
  NAND2_X1 U590 ( .A1(n606), .A2(n699), .ZN(n505) );
  XNOR2_X1 U591 ( .A(n505), .B(KEYINPUT93), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n507), .A2(n506), .ZN(n712) );
  NAND2_X1 U593 ( .A1(n509), .A2(n508), .ZN(n554) );
  AND2_X1 U594 ( .A1(n712), .A2(n554), .ZN(n672) );
  INV_X1 U595 ( .A(n555), .ZN(n511) );
  NAND2_X1 U596 ( .A1(n659), .A2(n511), .ZN(n512) );
  OR2_X1 U597 ( .A1(n512), .A2(n353), .ZN(n513) );
  OR2_X1 U598 ( .A1(n514), .A2(n513), .ZN(n605) );
  AND2_X1 U599 ( .A1(n515), .A2(n605), .ZN(n516) );
  NAND2_X1 U600 ( .A1(n630), .A2(KEYINPUT84), .ZN(n520) );
  AND2_X1 U601 ( .A1(n628), .A2(KEYINPUT44), .ZN(n518) );
  AND2_X1 U602 ( .A1(n609), .A2(n518), .ZN(n519) );
  NAND2_X1 U603 ( .A1(n520), .A2(n519), .ZN(n523) );
  NAND2_X1 U604 ( .A1(n521), .A2(KEYINPUT84), .ZN(n522) );
  NAND2_X1 U605 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U606 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n526) );
  NOR2_X1 U607 ( .A1(G900), .A2(n727), .ZN(n528) );
  NAND2_X1 U608 ( .A1(n528), .A2(G902), .ZN(n530) );
  NAND2_X1 U609 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U610 ( .A1(n531), .A2(n687), .ZN(n539) );
  INV_X1 U611 ( .A(n539), .ZN(n562) );
  AND2_X1 U612 ( .A1(n562), .A2(n675), .ZN(n533) );
  NAND2_X1 U613 ( .A1(n662), .A2(n674), .ZN(n532) );
  XOR2_X1 U614 ( .A(KEYINPUT30), .B(n532), .Z(n561) );
  NAND2_X1 U615 ( .A1(n533), .A2(n561), .ZN(n534) );
  NOR2_X1 U616 ( .A1(n534), .A2(n567), .ZN(n535) );
  NOR2_X1 U617 ( .A1(n586), .A2(n554), .ZN(n538) );
  XNOR2_X1 U618 ( .A(KEYINPUT101), .B(KEYINPUT40), .ZN(n537) );
  XNOR2_X1 U619 ( .A(n538), .B(n537), .ZN(n732) );
  INV_X1 U620 ( .A(n658), .ZN(n540) );
  NOR2_X1 U621 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U622 ( .A1(n542), .A2(n541), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n544), .B(KEYINPUT28), .ZN(n546) );
  NAND2_X1 U624 ( .A1(n546), .A2(n545), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n675), .A2(n674), .ZN(n547) );
  XNOR2_X1 U626 ( .A(n547), .B(KEYINPUT102), .ZN(n673) );
  INV_X1 U627 ( .A(n673), .ZN(n548) );
  NAND2_X1 U628 ( .A1(n548), .A2(n676), .ZN(n550) );
  XNOR2_X1 U629 ( .A(KEYINPUT103), .B(KEYINPUT41), .ZN(n549) );
  XNOR2_X1 U630 ( .A(n550), .B(n549), .ZN(n690) );
  XOR2_X1 U631 ( .A(KEYINPUT42), .B(n551), .Z(n622) );
  NAND2_X1 U632 ( .A1(n732), .A2(n622), .ZN(n553) );
  XOR2_X1 U633 ( .A(KEYINPUT83), .B(KEYINPUT46), .Z(n552) );
  XNOR2_X1 U634 ( .A(n553), .B(n552), .ZN(n577) );
  XNOR2_X1 U635 ( .A(n554), .B(KEYINPUT99), .ZN(n607) );
  NAND2_X1 U636 ( .A1(n555), .A2(n607), .ZN(n556) );
  NOR2_X1 U637 ( .A1(n557), .A2(n556), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n580), .A2(n558), .ZN(n559) );
  XNOR2_X1 U639 ( .A(n559), .B(KEYINPUT36), .ZN(n560) );
  INV_X1 U640 ( .A(n664), .ZN(n582) );
  NOR2_X1 U641 ( .A1(n560), .A2(n582), .ZN(n716) );
  AND2_X1 U642 ( .A1(n562), .A2(n561), .ZN(n566) );
  NOR2_X1 U643 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U644 ( .A1(n566), .A2(n565), .ZN(n568) );
  NOR2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U646 ( .A1(n569), .A2(n502), .ZN(n708) );
  NOR2_X1 U647 ( .A1(n716), .A2(n708), .ZN(n575) );
  NOR2_X1 U648 ( .A1(n571), .A2(n570), .ZN(n703) );
  INV_X1 U649 ( .A(n672), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n703), .A2(n572), .ZN(n573) );
  XOR2_X1 U651 ( .A(KEYINPUT47), .B(n573), .Z(n574) );
  NAND2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U653 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U654 ( .A(KEYINPUT82), .B(KEYINPUT48), .Z(n578) );
  XNOR2_X1 U655 ( .A(n579), .B(n578), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n580), .A2(n674), .ZN(n581) );
  XOR2_X1 U657 ( .A(KEYINPUT100), .B(n581), .Z(n583) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT43), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n585), .A2(n563), .ZN(n621) );
  OR2_X1 U661 ( .A1(n586), .A2(n712), .ZN(n719) );
  NAND2_X1 U662 ( .A1(n621), .A2(n719), .ZN(n587) );
  OR2_X2 U663 ( .A1(n588), .A2(n587), .ZN(n723) );
  NOR2_X1 U664 ( .A1(n723), .A2(KEYINPUT81), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n612), .A2(n589), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n351), .A2(G472), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT62), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n727), .A2(G952), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n599), .B(n598), .ZN(G57) );
  XOR2_X1 U670 ( .A(KEYINPUT27), .B(KEYINPUT107), .Z(n601) );
  XNOR2_X1 U671 ( .A(G107), .B(KEYINPUT26), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n601), .B(n600), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT106), .B(n602), .Z(n604) );
  NOR2_X1 U674 ( .A1(n699), .A2(n712), .ZN(n603) );
  XOR2_X1 U675 ( .A(n604), .B(n603), .Z(G9) );
  XNOR2_X1 U676 ( .A(n605), .B(G101), .ZN(G3) );
  INV_X1 U677 ( .A(n607), .ZN(n709) );
  NOR2_X1 U678 ( .A1(n606), .A2(n709), .ZN(n608) );
  XOR2_X1 U679 ( .A(G113), .B(n608), .Z(G15) );
  XNOR2_X1 U680 ( .A(n609), .B(G110), .ZN(G12) );
  NOR2_X1 U681 ( .A1(n610), .A2(n611), .ZN(n620) );
  INV_X1 U682 ( .A(n612), .ZN(n613) );
  NOR2_X1 U683 ( .A1(n613), .A2(G953), .ZN(n618) );
  NAND2_X1 U684 ( .A1(G953), .A2(G224), .ZN(n614) );
  XNOR2_X1 U685 ( .A(KEYINPUT61), .B(n614), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n615), .A2(G898), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT123), .ZN(n617) );
  NOR2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U689 ( .A(n620), .B(n619), .Z(G69) );
  XNOR2_X1 U690 ( .A(n621), .B(G140), .ZN(G42) );
  XNOR2_X1 U691 ( .A(n622), .B(G137), .ZN(G39) );
  NOR2_X1 U692 ( .A1(n352), .A2(n623), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n626), .A2(n654), .ZN(n627) );
  XNOR2_X1 U695 ( .A(n627), .B(KEYINPUT122), .ZN(G63) );
  XNOR2_X1 U696 ( .A(n629), .B(n350), .ZN(G21) );
  XOR2_X1 U697 ( .A(n630), .B(G122), .Z(G24) );
  NAND2_X1 U698 ( .A1(n351), .A2(G217), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U700 ( .A1(n633), .A2(n654), .ZN(G66) );
  NOR2_X1 U701 ( .A1(n352), .A2(n634), .ZN(n638) );
  XOR2_X1 U702 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n635) );
  XNOR2_X1 U703 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U704 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n639), .A2(n654), .ZN(n640) );
  XNOR2_X1 U706 ( .A(n640), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U707 ( .A1(n351), .A2(G469), .ZN(n647) );
  XOR2_X1 U708 ( .A(KEYINPUT117), .B(KEYINPUT119), .Z(n643) );
  XNOR2_X1 U709 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(KEYINPUT58), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n649), .B(KEYINPUT120), .ZN(G54) );
  XOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n651) );
  XNOR2_X1 U715 ( .A(n650), .B(n651), .ZN(n652) );
  XNOR2_X1 U716 ( .A(n653), .B(n652), .ZN(n655) );
  NOR2_X2 U717 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U718 ( .A(n656), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U719 ( .A(n657), .B(KEYINPUT80), .ZN(n696) );
  NOR2_X1 U720 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U721 ( .A(KEYINPUT49), .B(n660), .Z(n661) );
  NOR2_X1 U722 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U723 ( .A(KEYINPUT113), .B(n663), .ZN(n667) );
  NOR2_X1 U724 ( .A1(n502), .A2(n353), .ZN(n665) );
  XNOR2_X1 U725 ( .A(n665), .B(KEYINPUT50), .ZN(n666) );
  OR2_X1 U726 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U727 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U728 ( .A(n670), .B(KEYINPUT51), .ZN(n671) );
  NOR2_X1 U729 ( .A1(n671), .A2(n690), .ZN(n685) );
  NOR2_X1 U730 ( .A1(n673), .A2(n672), .ZN(n681) );
  NOR2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n678) );
  INV_X1 U732 ( .A(n676), .ZN(n677) );
  NOR2_X1 U733 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U734 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  NOR2_X1 U735 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U736 ( .A1(n691), .A2(n682), .ZN(n683) );
  XOR2_X1 U737 ( .A(KEYINPUT115), .B(n683), .Z(n684) );
  NOR2_X1 U738 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U739 ( .A(n686), .B(KEYINPUT52), .Z(n689) );
  AND2_X1 U740 ( .A1(n687), .A2(G952), .ZN(n688) );
  NAND2_X1 U741 ( .A1(n689), .A2(n688), .ZN(n694) );
  NOR2_X1 U742 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U743 ( .A1(n692), .A2(G953), .ZN(n693) );
  NAND2_X1 U744 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U745 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U746 ( .A(KEYINPUT116), .B(KEYINPUT53), .ZN(n697) );
  XNOR2_X1 U747 ( .A(n698), .B(n697), .ZN(G75) );
  XOR2_X1 U748 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n701) );
  NOR2_X1 U749 ( .A1(n699), .A2(n709), .ZN(n700) );
  XOR2_X1 U750 ( .A(n701), .B(n700), .Z(n702) );
  XNOR2_X1 U751 ( .A(G104), .B(n702), .ZN(G6) );
  INV_X1 U752 ( .A(n703), .ZN(n710) );
  NOR2_X1 U753 ( .A1(n710), .A2(n712), .ZN(n707) );
  XOR2_X1 U754 ( .A(KEYINPUT108), .B(KEYINPUT29), .Z(n705) );
  XNOR2_X1 U755 ( .A(G128), .B(KEYINPUT109), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n707), .B(n706), .ZN(G30) );
  XOR2_X1 U758 ( .A(G143), .B(n708), .Z(G45) );
  NOR2_X1 U759 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U760 ( .A(G146), .B(n711), .Z(G48) );
  XOR2_X1 U761 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n714) );
  NOR2_X1 U762 ( .A1(n606), .A2(n712), .ZN(n713) );
  XOR2_X1 U763 ( .A(n714), .B(n713), .Z(n715) );
  XNOR2_X1 U764 ( .A(G116), .B(n715), .ZN(G18) );
  XNOR2_X1 U765 ( .A(n716), .B(KEYINPUT37), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n717), .B(KEYINPUT112), .ZN(n718) );
  XNOR2_X1 U767 ( .A(G125), .B(n718), .ZN(G27) );
  XNOR2_X1 U768 ( .A(G134), .B(n719), .ZN(G36) );
  XOR2_X1 U769 ( .A(KEYINPUT124), .B(n720), .Z(n721) );
  XNOR2_X1 U770 ( .A(n722), .B(n721), .ZN(n725) );
  XNOR2_X1 U771 ( .A(n723), .B(n725), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(n727), .ZN(n730) );
  XNOR2_X1 U773 ( .A(n725), .B(G227), .ZN(n726) );
  NOR2_X1 U774 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U775 ( .A1(G900), .A2(n728), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U777 ( .A(KEYINPUT125), .B(n731), .ZN(G72) );
  XNOR2_X1 U778 ( .A(G131), .B(n732), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(KEYINPUT126), .ZN(G33) );
endmodule

