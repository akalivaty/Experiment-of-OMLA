//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n208), .B2(new_n205), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n204), .B1(new_n216), .B2(KEYINPUT25), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n220), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n221), .A2(new_n212), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n229));
  INV_X1    g028(.A(new_n215), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n230), .A2(new_n211), .A3(new_n213), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT65), .B(new_n218), .C1(new_n231), .C2(new_n209), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n219), .A2(new_n233), .A3(new_n227), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n217), .A2(new_n229), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n222), .A2(new_n224), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT27), .B(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT69), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n242));
  INV_X1    g041(.A(G169gat), .ZN(new_n243));
  INV_X1    g042(.A(G176gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n205), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(KEYINPUT26), .B2(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n246), .A2(KEYINPUT26), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n247), .A2(new_n248), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n241), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n203), .B1(new_n235), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n203), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n235), .B2(new_n250), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G211gat), .ZN(new_n256));
  INV_X1    g055(.A(G218gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G197gat), .ZN(new_n259));
  INV_X1    g058(.A(G204gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262));
  OAI22_X1  g061(.A1(KEYINPUT22), .A2(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G211gat), .B(G218gat), .Z(new_n264));
  OR3_X1    g063(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT73), .B1(new_n263), .B2(new_n264), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n264), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(KEYINPUT72), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(KEYINPUT72), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n255), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n235), .A2(new_n250), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n253), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT74), .B1(new_n278), .B2(new_n251), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n254), .B2(new_n253), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n202), .B(new_n275), .C1(new_n282), .C2(new_n272), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n272), .B1(new_n279), .B2(new_n281), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT75), .B1(new_n284), .B2(new_n274), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n293));
  XOR2_X1   g092(.A(G127gat), .B(G134gat), .Z(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G141gat), .B(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n305), .B2(KEYINPUT77), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n304), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n314), .A2(KEYINPUT78), .B1(KEYINPUT2), .B2(new_n299), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n298), .A2(KEYINPUT79), .A3(new_n299), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n317));
  INV_X1    g116(.A(new_n299), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n297), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n312), .A2(new_n315), .A3(new_n316), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n296), .B(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n323), .B(KEYINPUT80), .Z(new_n324));
  AOI21_X1  g123(.A(new_n291), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n295), .B1(new_n321), .B2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n327), .A3(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n310), .A2(KEYINPUT81), .A3(new_n320), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT4), .A4(new_n295), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n296), .B2(new_n321), .ZN(new_n335));
  INV_X1    g134(.A(new_n324), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n329), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n325), .A2(new_n337), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT5), .B(new_n324), .C1(new_n326), .C2(new_n328), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n295), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT4), .B1(new_n296), .B2(new_n321), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(KEYINPUT82), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT82), .B1(new_n339), .B2(new_n342), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n346), .B2(new_n351), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n340), .A2(new_n341), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n329), .A2(new_n291), .A3(new_n336), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n358), .A2(new_n343), .B1(new_n325), .B2(new_n337), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n350), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT30), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n284), .A2(new_n274), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n288), .ZN(new_n364));
  NOR4_X1   g163(.A1(new_n284), .A2(new_n274), .A3(KEYINPUT30), .A4(new_n289), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n290), .B(new_n361), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n272), .B1(new_n277), .B2(new_n328), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n267), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n263), .A2(new_n264), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n265), .A2(KEYINPUT83), .A3(new_n266), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT3), .B1(new_n374), .B2(new_n277), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n331), .A2(new_n332), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n369), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT85), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n272), .A2(new_n382), .A3(new_n277), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n327), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n272), .B2(new_n277), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n321), .B(new_n381), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n367), .B1(new_n368), .B2(new_n379), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n378), .A2(new_n379), .B1(new_n386), .B2(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n390), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT31), .B(G50gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(KEYINPUT86), .A2(G22gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT86), .A2(G22gat), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n380), .A2(new_n388), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n397), .C1(new_n400), .C2(new_n393), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n276), .A2(new_n296), .ZN(new_n405));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n235), .A2(new_n295), .A3(new_n250), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT34), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT70), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n408), .B2(KEYINPUT70), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n415));
  XOR2_X1   g214(.A(G15gat), .B(G43gat), .Z(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n414), .B(new_n415), .C1(KEYINPUT33), .C2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n415), .B2(KEYINPUT33), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n415), .A2(new_n414), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n413), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  INV_X1    g223(.A(new_n412), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n410), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n421), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n404), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT35), .B1(new_n366), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT91), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT91), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(KEYINPUT35), .C1(new_n366), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n365), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n275), .B(new_n288), .C1(new_n282), .C2(new_n272), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT30), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n290), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT88), .B1(new_n359), .B2(new_n350), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT6), .B1(new_n359), .B2(new_n350), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n346), .A2(new_n442), .A3(new_n351), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n444), .A2(new_n352), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n399), .A2(new_n403), .ZN(new_n446));
  NOR4_X1   g245(.A1(new_n439), .A2(new_n445), .A3(new_n446), .A4(KEYINPUT35), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT71), .B1(new_n428), .B2(new_n423), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n423), .A2(KEYINPUT71), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n284), .A2(KEYINPUT37), .A3(new_n274), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n273), .B1(new_n279), .B2(new_n281), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT37), .B1(new_n255), .B2(new_n272), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OR3_X1    g256(.A1(new_n453), .A2(new_n457), .A3(new_n288), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n445), .A2(new_n458), .A3(KEYINPUT90), .A4(new_n436), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT37), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n289), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT38), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n352), .A3(new_n436), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n453), .A2(new_n457), .A3(new_n288), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n459), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n336), .B1(new_n342), .B2(new_n329), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n351), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT39), .B1(new_n322), .B2(new_n324), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n471), .B(new_n474), .C1(new_n469), .C2(new_n475), .ZN(new_n476));
  OR3_X1    g275(.A1(new_n476), .A2(new_n472), .A3(new_n473), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  AND4_X1   g277(.A1(new_n440), .A2(new_n477), .A3(new_n443), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n446), .B1(new_n439), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n450), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n428), .B2(new_n423), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n366), .A2(new_n446), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n452), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G197gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT11), .B(G169gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(KEYINPUT12), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT13), .Z(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G8gat), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT16), .ZN(new_n501));
  INV_X1    g300(.A(G22gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G15gat), .ZN(new_n503));
  INV_X1    g302(.A(G15gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G22gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n506), .B2(KEYINPUT94), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(G1gat), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI221_X1 g309(.A(new_n506), .B1(KEYINPUT94), .B2(new_n499), .C1(G1gat), .C2(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(KEYINPUT96), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT92), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G43gat), .ZN(new_n521));
  AOI21_X1  g320(.A(G50gat), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G50gat), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT93), .B1(new_n523), .B2(G43gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n518), .A3(G50gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n517), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT14), .B(G29gat), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G29gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n523), .A2(G43gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n518), .A2(G50gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n531), .B2(new_n533), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n516), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n538), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n528), .B2(new_n534), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n540), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n514), .A3(new_n515), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n498), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n539), .A2(KEYINPUT95), .A3(KEYINPUT17), .A4(new_n541), .ZN(new_n549));
  OR2_X1    g348(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g349(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n550), .B(new_n551), .C1(new_n545), .C2(new_n540), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n512), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n496), .A3(new_n547), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n548), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n512), .B1(new_n549), .B2(new_n552), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n546), .A2(new_n514), .A3(new_n515), .ZN(new_n560));
  INV_X1    g359(.A(new_n496), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT18), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n495), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n495), .A3(new_n563), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n489), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G64gat), .ZN(new_n576));
  INV_X1    g375(.A(G64gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G57gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n573), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT97), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n516), .B1(new_n584), .B2(new_n583), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n602));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT8), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n607), .A2(new_n610), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n553), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G190gat), .B(G218gat), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n542), .B2(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n626), .B2(new_n631), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n605), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n632), .A2(new_n633), .A3(new_n605), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G230gat), .ZN(new_n638));
  INV_X1    g437(.A(G233gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n583), .B1(new_n618), .B2(new_n623), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n615), .A2(new_n617), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n621), .A2(new_n616), .A3(new_n622), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n644), .A2(new_n574), .A3(new_n645), .A4(new_n582), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n624), .A2(KEYINPUT98), .A3(new_n574), .A4(new_n582), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT10), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n641), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n648), .A3(new_n640), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n600), .A2(new_n637), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n568), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n361), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n500), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n568), .A2(new_n439), .A3(new_n662), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n668), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n666), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n668), .B2(KEYINPUT42), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT99), .B(new_n672), .C1(new_n666), .C2(new_n667), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n484), .A2(new_n675), .A3(new_n486), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT36), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT100), .B1(new_n677), .B2(new_n485), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n663), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n450), .A2(new_n504), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n663), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n404), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(new_n361), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n599), .A2(new_n661), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n637), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n568), .A2(new_n532), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n488), .B1(new_n468), .B2(new_n480), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n431), .A2(new_n433), .B1(new_n447), .B2(new_n450), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT44), .B(new_n637), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n567), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n599), .A3(new_n661), .ZN(new_n696));
  INV_X1    g495(.A(new_n637), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n487), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n366), .A2(KEYINPUT101), .A3(new_n446), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n481), .A2(new_n676), .A3(new_n701), .A4(new_n678), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n697), .B1(new_n702), .B2(new_n452), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n694), .B(new_n696), .C1(new_n703), .C2(KEYINPUT44), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n361), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n691), .A2(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(new_n439), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(G36gat), .A3(new_n688), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n489), .A2(new_n567), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n704), .B2(new_n707), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT102), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  AND2_X1   g516(.A1(new_n519), .A2(new_n521), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n679), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n704), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n489), .A2(new_n567), .A3(new_n450), .A4(new_n689), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n722), .A2(new_n718), .B1(KEYINPUT103), .B2(KEYINPUT47), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n721), .B1(new_n720), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1330gat));
  OAI21_X1  g526(.A(G50gat), .B1(new_n704), .B2(new_n404), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n568), .A2(new_n523), .A3(new_n446), .A4(new_n689), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1331gat));
  NAND2_X1  g531(.A1(new_n702), .A2(new_n452), .ZN(new_n733));
  INV_X1    g532(.A(new_n661), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n600), .A2(new_n567), .A3(new_n637), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n361), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n575), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n707), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n736), .B2(new_n679), .ZN(new_n744));
  INV_X1    g543(.A(G71gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n450), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n736), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g547(.A1(new_n736), .A2(new_n404), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g549(.A1(new_n599), .A2(new_n567), .A3(new_n734), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n694), .B(new_n751), .C1(new_n703), .C2(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n361), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n686), .A2(new_n611), .A3(new_n661), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n599), .A2(new_n567), .ZN(new_n756));
  AND4_X1   g555(.A1(KEYINPUT51), .A2(new_n733), .A3(new_n637), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n703), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT104), .ZN(G1336gat));
  NOR2_X1   g560(.A1(KEYINPUT106), .A2(KEYINPUT52), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT106), .A2(KEYINPUT52), .ZN(new_n763));
  OAI21_X1  g562(.A(G92gat), .B1(new_n752), .B2(new_n707), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n439), .A2(new_n612), .A3(new_n661), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT105), .Z(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n757), .B2(new_n758), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n767), .ZN(new_n768));
  AND4_X1   g567(.A1(KEYINPUT106), .A2(new_n764), .A3(new_n767), .A4(KEYINPUT52), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n752), .B2(new_n679), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT108), .B(G99gat), .Z(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n752), .A2(new_n771), .A3(new_n679), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n757), .A2(new_n758), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n450), .A2(new_n661), .A3(new_n773), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(G1338gat));
  OAI21_X1  g578(.A(G106gat), .B1(new_n752), .B2(new_n404), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n404), .A2(G106gat), .A3(new_n734), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n757), .B2(new_n758), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g583(.A1(new_n662), .A2(new_n695), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n647), .A2(new_n648), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n650), .ZN(new_n787));
  INV_X1    g586(.A(new_n651), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n640), .A3(new_n788), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n652), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n641), .B(new_n791), .C1(new_n649), .C2(new_n651), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n658), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(KEYINPUT110), .A3(new_n658), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT111), .B1(new_n797), .B2(KEYINPUT55), .ZN(new_n798));
  INV_X1    g597(.A(new_n660), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n797), .B2(KEYINPUT55), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n652), .ZN(new_n801));
  INV_X1    g600(.A(new_n796), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT110), .B1(new_n792), .B2(new_n658), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n798), .A2(new_n800), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT112), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n798), .A2(new_n800), .A3(new_n810), .A4(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n567), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n561), .B1(new_n559), .B2(new_n560), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n543), .A2(new_n547), .A3(new_n498), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n493), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT113), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n813), .B2(new_n814), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n817), .A2(new_n566), .A3(new_n661), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n637), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n818), .B(KEYINPUT113), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n637), .A2(new_n566), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n824), .A3(new_n811), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n827), .A3(new_n824), .A4(new_n811), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n822), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n785), .B1(new_n829), .B2(new_n599), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n686), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n439), .A2(new_n429), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n567), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n830), .A2(new_n404), .A3(new_n450), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n439), .A2(new_n361), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(G113gat), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n695), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n835), .A2(new_n840), .ZN(G1340gat));
  AOI21_X1  g640(.A(G120gat), .B1(new_n834), .B2(new_n661), .ZN(new_n842));
  INV_X1    g641(.A(G120gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n843), .A3(new_n734), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(G1341gat));
  OAI21_X1  g644(.A(G127gat), .B1(new_n838), .B2(new_n600), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n600), .A2(G127gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n833), .B2(new_n847), .ZN(G1342gat));
  OAI21_X1  g647(.A(G134gat), .B1(new_n838), .B2(new_n697), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n697), .A2(G134gat), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT56), .B1(new_n833), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n831), .A2(new_n853), .A3(new_n832), .A4(new_n850), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT115), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1343gat));
  XNOR2_X1  g658(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n679), .A2(new_n837), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n404), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n785), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n826), .A2(new_n828), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT55), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n558), .A2(new_n495), .A3(new_n563), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n868), .B(new_n660), .C1(new_n869), .C2(new_n564), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n797), .A2(KEYINPUT117), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(new_n804), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n821), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n823), .A2(KEYINPUT116), .A3(new_n566), .A4(new_n661), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n697), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT118), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n881), .B(new_n697), .C1(new_n874), .C2(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n600), .B1(new_n867), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n866), .B1(new_n884), .B2(KEYINPUT119), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n826), .A2(new_n828), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n599), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n865), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n830), .B2(new_n446), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n567), .B(new_n862), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G141gat), .ZN(new_n894));
  AND4_X1   g693(.A1(new_n707), .A2(new_n676), .A3(new_n446), .A4(new_n678), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n830), .A2(new_n686), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n695), .A2(G141gat), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT120), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n860), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n860), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n899), .B(new_n902), .C1(new_n893), .C2(G141gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(new_n896), .ZN(new_n905));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n661), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n785), .B1(new_n888), .B2(new_n889), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n884), .A2(KEYINPUT119), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n864), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n892), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n861), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT59), .B(new_n906), .C1(new_n912), .C2(new_n661), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n830), .A2(KEYINPUT57), .A3(new_n446), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n824), .A2(new_n807), .A3(new_n800), .A4(new_n798), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n599), .B1(new_n879), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n446), .B1(new_n917), .B2(new_n866), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n863), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n661), .A3(new_n862), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n914), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n907), .B1(new_n913), .B2(new_n922), .ZN(G1345gat));
  INV_X1    g722(.A(G155gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n924), .A3(new_n599), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n912), .A2(new_n599), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n924), .ZN(G1346gat));
  OR3_X1    g726(.A1(new_n896), .A2(G162gat), .A3(new_n697), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n697), .B(new_n861), .C1(new_n910), .C2(new_n911), .ZN(new_n929));
  OAI21_X1  g728(.A(G162gat), .B1(new_n929), .B2(KEYINPUT122), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n912), .A2(KEYINPUT122), .A3(new_n637), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n707), .A2(new_n686), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n836), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(G169gat), .A3(new_n567), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n830), .A2(new_n361), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n707), .A2(new_n429), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n243), .B1(new_n940), .B2(new_n695), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n936), .A2(KEYINPUT124), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1348gat));
  INV_X1    g745(.A(new_n940), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n244), .A3(new_n661), .ZN(new_n948));
  OAI21_X1  g747(.A(G176gat), .B1(new_n934), .B2(new_n734), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n947), .A2(new_n237), .A3(new_n599), .ZN(new_n951));
  OAI21_X1  g750(.A(G183gat), .B1(new_n934), .B2(new_n600), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1350gat));
  NAND3_X1  g756(.A1(new_n947), .A2(new_n236), .A3(new_n637), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n935), .A2(new_n637), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(G190gat), .ZN(new_n961));
  INV_X1    g760(.A(G190gat), .ZN(new_n962));
  AOI211_X1 g761(.A(KEYINPUT61), .B(new_n962), .C1(new_n935), .C2(new_n637), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n958), .B1(new_n961), .B2(new_n963), .ZN(G1351gat));
  NAND3_X1  g763(.A1(new_n676), .A2(new_n678), .A3(new_n933), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n920), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n967), .A2(new_n259), .A3(new_n695), .ZN(new_n968));
  AND4_X1   g767(.A1(new_n439), .A2(new_n676), .A3(new_n446), .A4(new_n678), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n937), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n567), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n973), .B2(new_n259), .ZN(G1352gat));
  AND2_X1   g773(.A1(new_n920), .A2(new_n966), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n260), .B1(new_n975), .B2(new_n661), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n734), .A2(G204gat), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n830), .A2(new_n361), .A3(new_n969), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT62), .ZN(new_n979));
  OAI21_X1  g778(.A(KEYINPUT127), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n979), .ZN(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n967), .B2(new_n734), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n980), .A2(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n972), .A2(new_n256), .A3(new_n599), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n920), .A2(new_n599), .A3(new_n679), .A4(new_n933), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n257), .A3(new_n637), .ZN(new_n991));
  OAI21_X1  g790(.A(G218gat), .B1(new_n967), .B2(new_n697), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1355gat));
endmodule


