//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI22_X1  g0024(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n220), .B(new_n225), .C1(G58), .C2(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT66), .B(G238), .Z(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n226), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n215), .B(new_n234), .C1(new_n211), .C2(new_n214), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n252), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n258), .B2(G226), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n262), .B(new_n264), .C1(new_n265), .C2(new_n263), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n206), .B1(G33), .B2(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n267), .C1(G77), .C2(new_n262), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(new_n260), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n261), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G190), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G13), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n273), .A2(new_n207), .A3(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n206), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G1), .B2(new_n207), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n278), .B2(G50), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT69), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n203), .A2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G58), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n281), .B1(new_n282), .B2(new_n284), .C1(new_n290), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n276), .A2(new_n206), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n280), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n272), .B1(new_n297), .B2(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n270), .A2(G200), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n298), .B(new_n299), .C1(KEYINPUT9), .C2(new_n297), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n305));
  INV_X1    g0105(.A(G232), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G226), .B2(G1698), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT3), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n304), .B(new_n305), .C1(new_n308), .C2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(new_n267), .B1(G238), .B2(new_n258), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n254), .B(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(G179), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT14), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT12), .ZN(new_n328));
  INV_X1    g0128(.A(new_n274), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(G68), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n227), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(new_n278), .C2(new_n227), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT74), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n292), .A2(G77), .B1(G20), .B2(new_n227), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n283), .A2(G50), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n277), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g0136(.A(new_n336), .B(KEYINPUT11), .Z(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n320), .B2(G190), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n320), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n312), .B1(new_n228), .B2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n306), .B2(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n267), .C1(G107), .C2(new_n262), .ZN(new_n345));
  INV_X1    g0145(.A(G41), .ZN(new_n346));
  INV_X1    g0146(.A(G45), .ZN(new_n347));
  AOI21_X1  g0147(.A(G1), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G274), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n345), .B(new_n349), .C1(new_n217), .C2(new_n257), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT70), .B(G179), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n325), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT15), .B(G87), .Z(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n292), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n283), .B(KEYINPUT71), .Z(new_n356));
  OAI221_X1 g0156(.A(new_n355), .B1(new_n207), .B2(new_n216), .C1(new_n356), .C2(new_n285), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n295), .B1(new_n216), .B2(new_n274), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n216), .B2(new_n278), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n301), .A2(new_n339), .A3(new_n342), .A4(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(KEYINPUT3), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n310), .A2(KEYINPUT76), .ZN(new_n364));
  OAI21_X1  g0164(.A(G33), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n310), .B2(G33), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n291), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n263), .A2(G226), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n265), .A2(new_n263), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n365), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  XOR2_X1   g0173(.A(new_n373), .B(KEYINPUT80), .Z(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n267), .ZN(new_n376));
  INV_X1    g0176(.A(new_n351), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n349), .B1(new_n257), .B2(new_n306), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT81), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT81), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n349), .C1(new_n257), .C2(new_n306), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT82), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n256), .B1(new_n372), .B2(new_n374), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n325), .B1(new_n385), .B2(new_n378), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n384), .B1(new_n383), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n310), .A2(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n362), .A2(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G33), .B1(new_n367), .B2(new_n368), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n390), .B(new_n393), .C1(new_n397), .C2(G20), .ZN(new_n398));
  XNOR2_X1  g0198(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n291), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT75), .B1(new_n291), .B2(KEYINPUT3), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n399), .A2(new_n291), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n402), .A2(new_n391), .A3(new_n392), .A4(new_n207), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(G68), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(G58), .B(G68), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n394), .A2(new_n395), .A3(new_n291), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n311), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT7), .B1(new_n312), .B2(new_n207), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n227), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n406), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n295), .A3(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n278), .A2(new_n289), .A3(new_n287), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n274), .B1(new_n287), .B2(new_n289), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT78), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n418), .A2(KEYINPUT78), .A3(new_n419), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT79), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n417), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n417), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n389), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT18), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n376), .A2(new_n271), .A3(new_n382), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n341), .B1(new_n385), .B2(new_n378), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n417), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT17), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n389), .C1(new_n426), .C2(new_n427), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n297), .B1(new_n325), .B2(new_n270), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n270), .B2(new_n351), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n359), .B1(G200), .B2(new_n350), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n271), .B2(new_n350), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n361), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT91), .ZN(new_n444));
  INV_X1    g0244(.A(G303), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n262), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n222), .A2(G1698), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n397), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n224), .A2(new_n263), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n369), .B(new_n449), .C1(new_n291), .C2(new_n399), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT88), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n397), .A2(KEYINPUT88), .A3(new_n449), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT89), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT89), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n448), .A2(new_n452), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n267), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT90), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n251), .B(G45), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n464), .A2(new_n253), .ZN(new_n465));
  INV_X1    g0265(.A(G270), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n256), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n458), .A2(KEYINPUT90), .A3(new_n267), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n461), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(new_n207), .C1(G33), .C2(new_n221), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(new_n295), .C1(new_n207), .C2(G116), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT20), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n274), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n329), .B(new_n277), .C1(G1), .C2(new_n291), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G169), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT21), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n444), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(KEYINPUT91), .B(KEYINPUT21), .C1(new_n471), .C2(new_n481), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(KEYINPUT21), .A3(new_n481), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT90), .B1(new_n458), .B2(new_n267), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n460), .B(new_n256), .C1(new_n455), .C2(new_n457), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(G179), .A3(new_n479), .A4(new_n469), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n484), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n479), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n471), .B2(new_n271), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n487), .A2(new_n488), .A3(new_n468), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n341), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT92), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n479), .B1(new_n495), .B2(G190), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT92), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n471), .A2(G200), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT25), .B1(new_n329), .B2(G107), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n329), .A2(KEYINPUT25), .A3(G107), .ZN(new_n504));
  INV_X1    g0304(.A(new_n478), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G107), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n218), .A2(G20), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n365), .A2(KEYINPUT22), .A3(new_n369), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n309), .A3(new_n311), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n207), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n223), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n509), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n292), .A2(G116), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT24), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n508), .A2(new_n514), .A3(new_n518), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT93), .B1(new_n520), .B2(new_n295), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT93), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n522), .B(new_n277), .C1(new_n517), .C2(new_n519), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n503), .B(new_n506), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n397), .B1(G250), .B2(G1698), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n263), .A2(G257), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT94), .B(G294), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n525), .A2(new_n526), .B1(new_n291), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n267), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n467), .A2(new_n224), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n530), .A2(G179), .A3(new_n465), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT95), .ZN(new_n534));
  INV_X1    g0334(.A(new_n465), .ZN(new_n535));
  AOI211_X1 g0335(.A(new_n535), .B(new_n531), .C1(new_n529), .C2(new_n267), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n533), .B(new_n534), .C1(new_n536), .C2(new_n325), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(KEYINPUT95), .A3(G179), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n524), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n531), .B1(new_n529), .B2(new_n267), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n465), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n271), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n536), .A2(new_n341), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n524), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n217), .B2(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n365), .A2(new_n369), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n256), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(G274), .B1(KEYINPUT84), .B2(G250), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n251), .A2(G45), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT84), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n554), .A3(G250), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n267), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT85), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  INV_X1    g0358(.A(new_n556), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n397), .A2(new_n547), .B1(G33), .B2(G116), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n256), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n271), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n365), .A2(new_n207), .A3(G68), .A4(new_n369), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n304), .B2(new_n305), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n566), .B2(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n302), .A2(new_n565), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n295), .ZN(new_n570));
  INV_X1    g0370(.A(new_n354), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n274), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n572), .C1(new_n218), .C2(new_n478), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n562), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n557), .A2(new_n561), .A3(G200), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n557), .A2(new_n561), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n377), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n505), .A2(new_n354), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT86), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n557), .A2(new_n561), .A3(new_n325), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n570), .A2(new_n583), .A3(new_n572), .A4(new_n579), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n578), .A2(new_n581), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n283), .A2(G77), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n221), .A2(new_n223), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G97), .A2(G107), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n591), .B2(KEYINPUT6), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G20), .ZN(new_n593));
  AOI21_X1  g0393(.A(G20), .B1(new_n409), .B2(new_n311), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n412), .B1(new_n594), .B2(KEYINPUT7), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n587), .B(new_n593), .C1(new_n595), .C2(new_n223), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n295), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n274), .A2(new_n221), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n478), .B2(new_n221), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT4), .B1(new_n312), .B2(new_n219), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT4), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n402), .B2(new_n217), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n535), .B1(new_n607), .B2(new_n267), .ZN(new_n608));
  INV_X1    g0408(.A(new_n467), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G257), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n325), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n262), .B2(G250), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n472), .B(new_n606), .C1(new_n612), .C2(new_n263), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT4), .B1(new_n397), .B2(G244), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n267), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n465), .A3(new_n610), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n377), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n601), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT83), .B1(new_n597), .B2(new_n600), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  AOI211_X1 g0420(.A(new_n620), .B(new_n599), .C1(new_n596), .C2(new_n295), .ZN(new_n621));
  AOI21_X1  g0421(.A(G200), .B1(new_n608), .B2(new_n610), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n271), .A2(new_n615), .A3(new_n465), .A4(new_n610), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n619), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n586), .A2(KEYINPUT87), .A3(new_n618), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n618), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n576), .A2(new_n585), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n545), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n443), .A2(new_n492), .A3(new_n502), .A4(new_n630), .ZN(G372));
  XNOR2_X1  g0431(.A(new_n301), .B(KEYINPUT97), .ZN(new_n632));
  INV_X1    g0432(.A(new_n339), .ZN(new_n633));
  INV_X1    g0433(.A(new_n360), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n342), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n434), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n417), .A2(new_n424), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n383), .A2(new_n386), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT82), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n637), .B1(new_n389), .B2(new_n638), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n435), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n417), .A2(new_n424), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n639), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT96), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n389), .A2(new_n637), .A3(new_n638), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n636), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n632), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n439), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT98), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n653), .B(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n480), .B1(new_n489), .B2(new_n469), .ZN(new_n656));
  INV_X1    g0456(.A(G179), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n487), .A2(new_n488), .A3(new_n657), .A4(new_n468), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n656), .A2(KEYINPUT21), .B1(new_n658), .B2(new_n479), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT91), .B1(new_n656), .B2(KEYINPUT21), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n482), .A2(new_n444), .A3(new_n483), .ZN(new_n661));
  INV_X1    g0461(.A(new_n539), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n544), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n559), .B1(new_n560), .B2(new_n256), .ZN(new_n665));
  AOI211_X1 g0465(.A(new_n573), .B(new_n562), .C1(G200), .C2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n627), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n325), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n578), .A2(new_n580), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n666), .A2(new_n670), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n619), .A2(new_n621), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n611), .A2(new_n617), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n628), .A2(new_n618), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(KEYINPUT26), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n668), .A2(new_n671), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n443), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n655), .A2(new_n681), .ZN(G369));
  NAND3_X1  g0482(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n251), .A2(new_n207), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n493), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n492), .A2(new_n502), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  INV_X1    g0494(.A(new_n524), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n545), .B1(new_n695), .B2(new_n690), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n662), .B2(new_n690), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(G330), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n663), .A2(new_n664), .A3(new_n690), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n213), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n564), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n210), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(KEYINPUT26), .B2(new_n676), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n668), .A2(new_n671), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n690), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n492), .A2(new_n630), .A3(new_n502), .A4(new_n690), .ZN(new_n713));
  INV_X1    g0513(.A(new_n616), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n540), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n658), .A2(new_n577), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n714), .A2(new_n351), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n471), .A2(new_n665), .A3(new_n541), .A4(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n658), .A2(KEYINPUT30), .A3(new_n577), .A4(new_n716), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n689), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n726), .A3(new_n689), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(G330), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n680), .A2(new_n729), .A3(new_n690), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n712), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT99), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT99), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n712), .A2(new_n733), .A3(new_n728), .A4(new_n730), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n707), .B1(new_n735), .B2(G1), .ZN(G364));
  AND2_X1   g0536(.A1(new_n694), .A2(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n207), .A2(G13), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT100), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n347), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n740), .A2(new_n251), .A3(new_n702), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n694), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n262), .A2(new_n213), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT101), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n745), .A2(G355), .B1(new_n476), .B2(new_n701), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT102), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n397), .A2(new_n701), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n210), .A2(G45), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n748), .B(new_n749), .C1(new_n246), .C2(new_n347), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n206), .B1(G20), .B2(new_n325), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n741), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n351), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(new_n271), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n351), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G200), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G311), .A2(new_n761), .B1(new_n764), .B2(G322), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n760), .A2(new_n341), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(KEYINPUT33), .B(G317), .Z(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G179), .A2(G200), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n207), .B1(new_n770), .B2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n341), .A2(G179), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n312), .B1(new_n528), .B2(new_n771), .C1(new_n776), .C2(new_n445), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n759), .A2(new_n770), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n769), .B(new_n777), .C1(G329), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT103), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n763), .B2(new_n341), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n351), .A2(KEYINPUT103), .A3(G200), .A4(new_n762), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G326), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n772), .A2(new_n759), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT105), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n780), .B(new_n785), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT106), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(new_n223), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G68), .B2(new_n766), .ZN(new_n792));
  INV_X1    g0592(.A(new_n764), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n288), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n779), .A2(G159), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(new_n761), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n776), .A2(new_n218), .B1(new_n216), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n794), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n771), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G97), .ZN(new_n801));
  INV_X1    g0601(.A(new_n784), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n799), .B(new_n801), .C1(new_n202), .C2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n790), .B1(new_n312), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n758), .B1(new_n804), .B2(new_n755), .ZN(new_n805));
  INV_X1    g0605(.A(new_n754), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n757), .B(new_n805), .C1(new_n694), .C2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n743), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n680), .A2(new_n690), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n359), .A2(new_n689), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n441), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n360), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n634), .A2(new_n690), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n680), .A2(new_n690), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(new_n728), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n758), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n817), .A2(new_n753), .ZN(new_n822));
  INV_X1    g0622(.A(new_n755), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n776), .A2(new_n202), .B1(new_n227), .B2(new_n788), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n397), .B1(new_n288), .B2(new_n771), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT109), .B(G143), .Z(new_n826));
  AOI22_X1  g0626(.A1(G159), .A2(new_n761), .B1(new_n764), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n282), .B2(new_n767), .C1(new_n802), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n824), .B(new_n825), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n830), .B2(new_n829), .C1(new_n832), .C2(new_n778), .ZN(new_n833));
  INV_X1    g0633(.A(new_n788), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(G87), .B1(G311), .B2(new_n779), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT108), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n312), .B1(new_n776), .B2(new_n223), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT107), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n766), .A2(G283), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n801), .B1(new_n793), .B2(new_n840), .C1(new_n476), .C2(new_n797), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G303), .B2(new_n784), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n823), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n755), .A2(new_n752), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(G77), .ZN(new_n847));
  OR4_X1    g0647(.A1(new_n758), .A2(new_n822), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n821), .A2(new_n848), .ZN(G384));
  AND2_X1   g0649(.A1(new_n592), .A2(KEYINPUT35), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n592), .A2(KEYINPUT35), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n850), .A2(new_n851), .A3(new_n476), .A4(new_n209), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI21_X1  g0653(.A(G77), .B1(new_n288), .B2(new_n227), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n854), .A2(new_n210), .B1(G50), .B2(new_n227), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(G1), .A3(new_n273), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n739), .A2(G1), .ZN(new_n857));
  INV_X1    g0657(.A(new_n687), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n407), .A2(new_n295), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n404), .B2(new_n406), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n424), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n437), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n646), .A2(new_n687), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n861), .ZN(new_n864));
  INV_X1    g0664(.A(new_n433), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n863), .B1(new_n427), .B2(new_n426), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n433), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n338), .A2(new_n689), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n339), .A2(new_n342), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT110), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n339), .A2(KEYINPUT110), .A3(new_n342), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n633), .A2(new_n689), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n815), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n875), .A2(new_n725), .A3(new_n727), .A4(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n644), .A2(new_n434), .A3(new_n649), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n858), .B1(new_n426), .B2(new_n427), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n888), .A2(new_n647), .A3(new_n433), .A4(new_n648), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n869), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n872), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n885), .B1(new_n895), .B2(new_n874), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n896), .A2(new_n725), .A3(new_n727), .A4(new_n883), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n725), .A2(new_n727), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n443), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n898), .B(new_n900), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(G330), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n818), .A2(new_n814), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n881), .A2(new_n882), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n875), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n650), .A2(new_n858), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n890), .B2(new_n893), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n339), .A2(new_n689), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n905), .A2(new_n907), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n730), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n729), .B1(new_n710), .B2(new_n690), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n443), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n655), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n915), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n857), .B1(new_n902), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT111), .Z(new_n922));
  AND2_X1   g0722(.A1(new_n902), .A2(new_n920), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n853), .B(new_n856), .C1(new_n922), .C2(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n683), .A2(new_n690), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n675), .A2(new_n689), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n624), .B(new_n618), .C1(new_n673), .C2(new_n690), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n545), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n925), .A2(new_n539), .A3(new_n544), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT42), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n933), .A3(new_n929), .ZN(new_n934));
  INV_X1    g0734(.A(new_n929), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n618), .B1(new_n935), .B2(new_n662), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n690), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n931), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n573), .A2(new_n689), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n672), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n671), .B2(new_n939), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n698), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n944), .A3(new_n929), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n938), .B(new_n942), .C1(new_n698), .C2(new_n935), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n702), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n663), .A2(new_n627), .A3(new_n664), .A4(new_n690), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(KEYINPUT44), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT45), .B1(new_n699), .B2(new_n929), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n953), .B(new_n954), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT112), .ZN(new_n958));
  AND4_X1   g0758(.A1(new_n958), .A2(new_n694), .A3(G330), .A4(new_n697), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n926), .A2(new_n697), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n932), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n698), .B1(new_n737), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n957), .A2(new_n959), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n735), .A2(new_n960), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n951), .B1(new_n967), .B2(new_n735), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n740), .A2(new_n251), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n949), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n748), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n756), .B1(new_n213), .B2(new_n571), .C1(new_n972), .C2(new_n242), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n741), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT113), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n784), .A2(G311), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n786), .B2(new_n797), .C1(new_n445), .C2(new_n793), .ZN(new_n977));
  INV_X1    g0777(.A(new_n776), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT46), .B1(new_n978), .B2(G116), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n402), .B1(new_n223), .B2(new_n771), .C1(new_n980), .C2(new_n778), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n221), .C2(new_n787), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n977), .B(new_n984), .C1(new_n527), .C2(new_n766), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n978), .A2(G58), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G137), .A2(new_n779), .B1(new_n800), .B2(G68), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n262), .C1(new_n216), .C2(new_n787), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G150), .A2(new_n764), .B1(new_n766), .B2(G159), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n202), .B2(new_n797), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(new_n784), .C2(new_n826), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n985), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n975), .B1(new_n806), .B2(new_n941), .C1(new_n993), .C2(new_n823), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n971), .A2(new_n994), .ZN(G387));
  NAND2_X1  g0795(.A1(new_n735), .A2(new_n964), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n732), .A2(new_n734), .A3(new_n963), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n702), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n779), .A2(G326), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G303), .A2(new_n761), .B1(new_n766), .B2(G311), .ZN(new_n1000));
  INV_X1    g0800(.A(G322), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n980), .B2(new_n793), .C1(new_n802), .C2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT48), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n786), .B2(new_n771), .C1(new_n528), .C2(new_n776), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n397), .B(new_n999), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .C1(new_n476), .C2(new_n787), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n571), .A2(new_n771), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n978), .A2(G77), .B1(G68), .B2(new_n761), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n282), .B2(new_n778), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G159), .C2(new_n784), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n202), .A2(new_n793), .B1(new_n767), .B2(new_n290), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G97), .B2(new_n834), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n397), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT114), .Z(new_n1015));
  AOI21_X1  g0815(.A(new_n823), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n285), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT50), .B1(new_n285), .B2(G50), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1017), .A2(new_n1018), .A3(new_n347), .A4(new_n704), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G68), .B2(G77), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n748), .B1(new_n239), .B2(new_n347), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n745), .B1(G116), .B2(new_n564), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n223), .B2(new_n701), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1024), .A2(new_n754), .A3(new_n755), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n697), .A2(new_n806), .ZN(new_n1026));
  NOR4_X1   g0826(.A1(new_n1016), .A2(new_n758), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n964), .B2(new_n970), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n998), .A2(new_n1028), .ZN(G393));
  OAI21_X1  g0829(.A(new_n397), .B1(new_n216), .B2(new_n771), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n978), .A2(G68), .B1(new_n834), .B2(G87), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n285), .B2(new_n797), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(new_n779), .C2(new_n826), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n784), .A2(G150), .B1(G159), .B2(new_n764), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT51), .Z(new_n1035));
  OAI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(new_n202), .C2(new_n767), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n784), .A2(G317), .B1(G311), .B2(new_n764), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  OAI22_X1  g0838(.A1(new_n840), .A2(new_n797), .B1(new_n767), .B2(new_n445), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n312), .B1(new_n778), .B2(new_n1001), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n771), .A2(new_n476), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1039), .A2(new_n791), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1038), .B(new_n1042), .C1(new_n786), .C2(new_n776), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n758), .B1(new_n1044), .B2(new_n755), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n756), .B1(new_n221), .B2(new_n213), .C1(new_n972), .C2(new_n249), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n806), .C2(new_n929), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n957), .B(new_n944), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n969), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n963), .B(new_n965), .C1(new_n732), .C2(new_n734), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n703), .B1(new_n1050), .B2(new_n960), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n996), .A2(new_n1048), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G390));
  NAND2_X1  g0854(.A1(new_n911), .A2(new_n912), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n752), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n764), .A2(G116), .B1(G77), .B2(new_n800), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n802), .A2(new_n786), .B1(new_n1057), .B2(KEYINPUT117), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n767), .A2(new_n223), .B1(new_n788), .B2(new_n227), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n312), .B1(new_n776), .B2(new_n218), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G294), .C2(new_n779), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n221), .B2(new_n797), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1058), .B(new_n1062), .C1(KEYINPUT117), .C2(new_n1057), .ZN(new_n1063));
  INV_X1    g0863(.A(G159), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n262), .B1(new_n771), .B2(new_n1064), .C1(new_n202), .C2(new_n787), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G125), .B2(new_n779), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT54), .B(G143), .Z(new_n1067));
  AOI22_X1  g0867(.A1(G132), .A2(new_n764), .B1(new_n761), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(new_n828), .C2(new_n767), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n978), .A2(G150), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT53), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(G128), .C2(new_n784), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1063), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1073), .A2(new_n755), .B1(new_n290), .B2(new_n845), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1056), .A2(new_n741), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n725), .A2(G330), .A3(new_n727), .A4(new_n883), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT115), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n913), .B1(new_n895), .B2(new_n874), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n710), .A2(new_n690), .A3(new_n813), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(new_n814), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n904), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n818), .B2(new_n814), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1055), .B1(new_n1083), .B2(new_n913), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1077), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1076), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1075), .B1(new_n1088), .B2(new_n969), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n725), .A2(G330), .A3(new_n727), .A4(new_n817), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT116), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n1091), .A3(new_n1081), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1090), .A2(new_n1081), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1076), .A2(KEYINPUT116), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n903), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1081), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1080), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n899), .A2(new_n443), .A3(G330), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n655), .A2(new_n918), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1088), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1077), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1078), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1079), .A2(new_n814), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n904), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n903), .A2(new_n904), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n913), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1112), .B2(new_n1055), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1106), .B1(new_n1113), .B2(new_n1086), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1102), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n703), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1089), .B1(new_n1105), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(G378));
  INV_X1    g0918(.A(KEYINPUT57), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n886), .A2(G330), .A3(new_n897), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n915), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n875), .B2(new_n1083), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n886), .A2(G330), .A3(new_n897), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n907), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n297), .A2(new_n687), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT97), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n301), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n301), .A2(new_n1130), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n439), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT119), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT119), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n632), .A2(new_n1135), .A3(new_n439), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1129), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1129), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1127), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1127), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1141), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1126), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1121), .A2(new_n1125), .A3(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1102), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1119), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1103), .B1(new_n1088), .B2(new_n1104), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1121), .A2(new_n1144), .A3(new_n1125), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1144), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1154), .A3(KEYINPUT57), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n1155), .A3(new_n702), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n846), .A2(G50), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n397), .A2(G33), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G50), .B1(new_n1158), .B2(new_n346), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n978), .A2(G77), .B1(G97), .B2(new_n766), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n223), .B2(new_n793), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n346), .B1(new_n787), .B2(new_n288), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n402), .B1(new_n227), .B2(new_n771), .C1(new_n786), .C2(new_n778), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n476), .B2(new_n802), .C1(new_n571), .C2(new_n797), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT58), .Z(new_n1166));
  AOI22_X1  g0966(.A1(new_n978), .A2(new_n1067), .B1(G128), .B2(new_n764), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT118), .Z(new_n1168));
  OAI22_X1  g0968(.A1(new_n797), .A2(new_n828), .B1(new_n282), .B2(new_n771), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n784), .B2(G125), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n832), .C2(new_n767), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT59), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n291), .B1(new_n787), .B2(new_n1064), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n779), .B2(G124), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1159), .B(new_n1166), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n741), .B1(new_n1176), .B2(new_n823), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1157), .B(new_n1177), .C1(new_n1145), .C2(new_n752), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1154), .B2(new_n970), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1156), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT120), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1156), .A2(new_n1182), .A3(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(G375));
  NOR2_X1   g0984(.A1(new_n904), .A2(new_n753), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT121), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT121), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n776), .A2(new_n221), .B1(new_n476), .B2(new_n767), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G77), .B2(new_n834), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n312), .B1(new_n778), .B2(new_n445), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1190), .B(new_n1008), .C1(G107), .C2(new_n761), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n786), .B2(new_n793), .C1(new_n840), .C2(new_n802), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n978), .A2(G159), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n787), .A2(new_n288), .B1(new_n771), .B2(new_n202), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n402), .B(new_n1195), .C1(G128), .C2(new_n779), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G150), .A2(new_n761), .B1(new_n766), .B2(new_n1067), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n832), .B2(new_n802), .C1(new_n828), .C2(new_n793), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n823), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n227), .B2(new_n845), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1186), .A2(new_n1187), .A3(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1100), .A2(new_n970), .B1(new_n741), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1095), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n950), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1203), .B1(new_n1205), .B2(new_n1115), .ZN(G381));
  AND3_X1   g1006(.A1(new_n1156), .A2(new_n1182), .A3(new_n1179), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1182), .B1(new_n1156), .B2(new_n1179), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1207), .A2(new_n1208), .A3(G378), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n998), .A2(new_n808), .A3(new_n1028), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G384), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT122), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n971), .A2(new_n1053), .A3(new_n994), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(G381), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1209), .A2(new_n1214), .A3(new_n1216), .ZN(G407));
  NAND3_X1  g1017(.A1(new_n1181), .A2(new_n1117), .A3(new_n1183), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G407), .B(G213), .C1(G343), .C2(new_n1218), .ZN(G409));
  NAND3_X1  g1019(.A1(new_n688), .A2(G213), .A3(G2897), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT60), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1204), .A2(KEYINPUT123), .A3(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1223), .A2(new_n702), .A3(new_n1104), .A4(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1226), .A2(G384), .A3(new_n1203), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G384), .B1(new_n1226), .B2(new_n1203), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1203), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1212), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(G384), .A3(new_n1203), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1220), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1180), .A2(G378), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1151), .A2(new_n1154), .A3(new_n950), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1117), .A2(new_n1179), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n688), .A2(G213), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT61), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n1239), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT62), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1117), .B1(new_n1156), .B2(new_n1179), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1244), .A2(KEYINPUT62), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1244), .A2(KEYINPUT62), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1248), .A2(new_n1242), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1241), .A2(new_n1245), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n808), .B1(new_n998), .B2(new_n1028), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1211), .A2(new_n1253), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n971), .A2(new_n1053), .A3(new_n994), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1053), .B1(new_n971), .B2(new_n994), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(G390), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1254), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1215), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1252), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1257), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1257), .A2(new_n1260), .A3(KEYINPUT124), .A4(new_n1263), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1266), .A2(new_n1267), .B1(new_n1240), .B2(new_n1234), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT125), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(KEYINPUT125), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1243), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1243), .A2(new_n1271), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1268), .A2(new_n1270), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1262), .A2(new_n1274), .ZN(G405));
  AND3_X1   g1075(.A1(new_n1218), .A2(new_n1261), .A3(new_n1235), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1261), .B1(new_n1218), .B2(new_n1235), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1242), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1261), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1209), .B2(new_n1246), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1218), .A2(new_n1261), .A3(new_n1235), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1242), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1279), .A2(new_n1283), .ZN(G402));
endmodule


