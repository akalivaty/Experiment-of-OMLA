//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G227), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n192), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT3), .B1(new_n197), .B2(G107), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G101), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT81), .B(G101), .Z(new_n205));
  OAI211_X1 g019(.A(new_n204), .B(KEYINPUT4), .C1(new_n205), .C2(new_n203), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(new_n207), .A3(G101), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT0), .A4(G128), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT0), .B(G128), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(G104), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n202), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n203), .B2(new_n205), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n215), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n215), .A3(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n212), .A2(KEYINPUT1), .A3(G146), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n227), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT10), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n209), .A2(new_n218), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n233), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n211), .A2(new_n229), .A3(new_n231), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n211), .A2(new_n229), .A3(new_n231), .A4(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(G128), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n244), .B2(new_n225), .ZN(new_n245));
  NOR4_X1   g059(.A1(new_n245), .A2(KEYINPUT82), .A3(new_n237), .A4(new_n223), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(G128), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n242), .B1(new_n249), .B2(new_n211), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n225), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n237), .B1(new_n251), .B2(new_n233), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n247), .B1(new_n252), .B2(new_n224), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n238), .B1(new_n246), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT64), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n260), .A3(new_n263), .A4(new_n258), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(G131), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n257), .A2(new_n260), .A3(new_n266), .A4(new_n258), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n262), .A2(new_n268), .A3(G131), .A4(new_n264), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n254), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n251), .A2(new_n233), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n236), .B1(new_n274), .B2(new_n224), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT12), .B1(new_n275), .B2(new_n272), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n196), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n272), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n254), .A2(KEYINPUT83), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n274), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT82), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n252), .A2(new_n247), .A3(new_n224), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT83), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n238), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n280), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n280), .A3(new_n238), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n195), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n191), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI211_X1 g109(.A(KEYINPUT84), .B(new_n191), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n286), .B1(new_n285), .B2(new_n238), .ZN(new_n298));
  INV_X1    g112(.A(new_n204), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT4), .B1(new_n203), .B2(new_n205), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n218), .B(new_n208), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n233), .A2(new_n234), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n223), .B1(new_n302), .B2(new_n227), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(KEYINPUT10), .ZN(new_n304));
  AOI211_X1 g118(.A(KEYINPUT83), .B(new_n304), .C1(new_n283), .C2(new_n284), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n272), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n195), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  INV_X1    g121(.A(new_n277), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT85), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n276), .B2(new_n277), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n310), .A2(new_n312), .A3(new_n289), .A4(new_n195), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n191), .B(new_n292), .C1(new_n307), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n196), .B1(new_n288), .B2(new_n273), .ZN(new_n318));
  AOI21_X1  g132(.A(G902), .B1(new_n318), .B2(new_n313), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT86), .A3(new_n191), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n190), .B1(new_n297), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT98), .ZN(new_n323));
  INV_X1    g137(.A(G478), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT15), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n212), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n226), .A2(G143), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n256), .ZN(new_n328));
  INV_X1    g142(.A(G122), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT92), .B1(new_n329), .B2(G116), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n331));
  INV_X1    g145(.A(G116), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G122), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n330), .A2(new_n333), .B1(G116), .B2(new_n329), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n200), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n226), .A2(G143), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT94), .A3(KEYINPUT13), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n327), .B1(new_n336), .B2(KEYINPUT13), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT93), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT93), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n340), .B(new_n327), .C1(new_n336), .C2(KEYINPUT13), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT13), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n326), .B2(new_n343), .ZN(new_n344));
  AND4_X1   g158(.A1(new_n337), .A2(new_n339), .A3(new_n341), .A4(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n328), .B(new_n335), .C1(new_n345), .C2(new_n256), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n256), .B1(new_n326), .B2(new_n327), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT95), .A3(new_n328), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT95), .ZN(new_n350));
  INV_X1    g164(.A(new_n328), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(new_n347), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n329), .A2(G116), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n200), .B1(new_n354), .B2(KEYINPUT14), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n334), .B(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT96), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT96), .B1(new_n353), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n346), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G217), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n188), .A2(new_n360), .A3(G953), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n346), .B(new_n361), .C1(new_n357), .C2(new_n358), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT97), .B1(new_n365), .B2(new_n292), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n367), .B(G902), .C1(new_n363), .C2(new_n364), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n325), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n292), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n367), .ZN(new_n371));
  INV_X1    g185(.A(new_n325), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n323), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(new_n373), .A3(new_n323), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n378));
  INV_X1    g192(.A(G125), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT75), .A2(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n382), .A2(KEYINPUT16), .A3(G140), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(G140), .A3(new_n381), .ZN(new_n385));
  NOR2_X1   g199(.A1(G125), .A2(G140), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT76), .B1(new_n388), .B2(KEYINPUT16), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT16), .ZN(new_n391));
  AOI211_X1 g205(.A(new_n390), .B(new_n391), .C1(new_n385), .C2(new_n387), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n384), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n210), .ZN(new_n394));
  OAI211_X1 g208(.A(G146), .B(new_n384), .C1(new_n389), .C2(new_n392), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  INV_X1    g210(.A(G237), .ZN(new_n397));
  INV_X1    g211(.A(G953), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G214), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n212), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n396), .B1(new_n400), .B2(G131), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n399), .B(G143), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT90), .A3(new_n266), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(G131), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n401), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(KEYINPUT17), .A3(G131), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n394), .A2(new_n395), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n197), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n402), .B1(new_n411), .B2(new_n266), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n400), .A2(KEYINPUT18), .A3(G131), .ZN(new_n413));
  XNOR2_X1  g227(.A(G125), .B(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n210), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n388), .B2(new_n210), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT89), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n408), .A2(new_n410), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n410), .B1(new_n408), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n292), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G475), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n401), .A2(new_n405), .A3(new_n403), .ZN(new_n427));
  AND2_X1   g241(.A1(KEYINPUT75), .A2(G125), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT75), .A2(G125), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n386), .B1(new_n430), .B2(G140), .ZN(new_n431));
  MUX2_X1   g245(.A(new_n414), .B(new_n431), .S(KEYINPUT19), .Z(new_n432));
  OAI211_X1 g246(.A(new_n427), .B(new_n395), .C1(G146), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n421), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n410), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(G475), .B1(new_n436), .B2(new_n422), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n292), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT91), .B1(new_n436), .B2(new_n422), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(KEYINPUT20), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n439), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n441), .A2(new_n442), .B1(new_n437), .B2(new_n292), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n426), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n377), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G234), .A2(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G952), .A3(new_n398), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT21), .B(G898), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(G902), .A3(G953), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G210), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT2), .B(G113), .Z(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G119), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT69), .A3(G116), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n332), .B2(G119), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n332), .A2(G119), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n458), .B(new_n461), .C1(new_n464), .C2(new_n463), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n206), .A2(new_n468), .A3(new_n208), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(G113), .B(new_n471), .C1(new_n465), .C2(new_n470), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n224), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(G110), .B(G122), .Z(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT6), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n469), .B2(new_n473), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n218), .A2(new_n430), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n245), .B2(new_n430), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT87), .B(G224), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G953), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n482), .B(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n477), .A2(new_n478), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n480), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT7), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT88), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n474), .B(KEYINPUT8), .Z(new_n493));
  INV_X1    g307(.A(new_n473), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n224), .B1(new_n467), .B2(new_n472), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n274), .A2(new_n382), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n481), .A4(new_n490), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n482), .A2(new_n491), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n492), .A2(new_n496), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n476), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n292), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n457), .B1(new_n488), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  INV_X1    g319(.A(new_n486), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n477), .A2(new_n478), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n479), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n505), .A2(new_n508), .A3(new_n292), .A4(new_n456), .ZN(new_n509));
  AOI211_X1 g323(.A(new_n447), .B(new_n455), .C1(new_n504), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n322), .A2(new_n445), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n226), .A2(G119), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n226), .A2(G119), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n514), .B2(new_n512), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT24), .B(G110), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT79), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(KEYINPUT79), .A3(new_n517), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n512), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n526));
  OAI22_X1  g340(.A1(new_n523), .A2(new_n525), .B1(new_n512), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT78), .B(G110), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n520), .B(new_n521), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n395), .A3(new_n415), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n394), .A2(new_n395), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(G110), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n516), .A2(new_n517), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND4_X1   g348(.A1(KEYINPUT77), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n394), .B2(new_n395), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT77), .B1(new_n536), .B2(new_n532), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n530), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n398), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n390), .B1(new_n431), .B2(new_n391), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n388), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G146), .B1(new_n546), .B2(new_n384), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n210), .B(new_n383), .C1(new_n544), .C2(new_n545), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n532), .B(new_n534), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n536), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n530), .A3(new_n541), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n292), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n543), .A2(new_n554), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n360), .B1(G234), .B2(new_n292), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT80), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT80), .ZN(new_n562));
  INV_X1    g376(.A(new_n560), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n562), .B(new_n563), .C1(new_n557), .C2(new_n558), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n541), .B1(new_n553), .B2(new_n530), .ZN(new_n565));
  INV_X1    g379(.A(new_n530), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n566), .B(new_n542), .C1(new_n551), .C2(new_n552), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n560), .A2(G902), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n561), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n259), .A2(G134), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n256), .A2(G137), .ZN(new_n575));
  OAI21_X1  g389(.A(G131), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n267), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT66), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n274), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n217), .B1(new_n270), .B2(new_n271), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n573), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n245), .A2(new_n577), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n272), .A2(new_n218), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT30), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n587), .A3(new_n468), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT70), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n466), .A2(new_n467), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n466), .B2(new_n467), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n585), .A2(new_n593), .A3(new_n586), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n397), .A2(new_n398), .A3(G210), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT27), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT26), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n219), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n582), .A2(new_n584), .A3(new_n592), .ZN(new_n603));
  INV_X1    g417(.A(new_n468), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n586), .B2(new_n580), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT28), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT71), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n603), .B2(KEYINPUT28), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT28), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n594), .A2(KEYINPUT71), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n600), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n602), .A2(new_n612), .A3(KEYINPUT29), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n593), .B1(new_n586), .B2(new_n585), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n603), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n608), .B(new_n610), .C1(new_n615), .C2(new_n609), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n599), .A2(KEYINPUT29), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n292), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n611), .A2(new_n600), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n588), .A2(new_n594), .A3(new_n599), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT31), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT31), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n588), .A2(new_n623), .A3(new_n594), .A4(new_n599), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n620), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(G472), .A2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT72), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT32), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT32), .ZN(new_n630));
  AOI211_X1 g444(.A(KEYINPUT72), .B(new_n630), .C1(new_n625), .C2(new_n626), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n619), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n572), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n511), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(new_n205), .Z(G3));
  INV_X1    g449(.A(new_n322), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT25), .B1(new_n568), .B2(new_n292), .ZN(new_n637));
  INV_X1    g451(.A(new_n558), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n560), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n562), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n559), .A2(KEYINPUT80), .A3(new_n560), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n570), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n625), .A2(new_n292), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(G472), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n627), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n636), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n504), .A2(new_n509), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(KEYINPUT99), .B(new_n457), .C1(new_n488), .C2(new_n503), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n446), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n455), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n324), .A2(new_n292), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n370), .A2(G478), .ZN(new_n655));
  NAND2_X1  g469(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n365), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n658));
  OAI21_X1  g472(.A(new_n657), .B1(new_n365), .B2(new_n658), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n654), .B(new_n655), .C1(new_n659), .C2(G478), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n444), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n646), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  AND2_X1   g479(.A1(KEYINPUT101), .A2(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g480(.A1(KEYINPUT101), .A2(KEYINPUT20), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n438), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n438), .A2(new_n667), .ZN(new_n669));
  INV_X1    g483(.A(new_n426), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n377), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n653), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n646), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n538), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n569), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n640), .A2(new_n641), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n511), .A2(new_n645), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT37), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G110), .ZN(G12));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n454), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n449), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n377), .A2(new_n651), .A3(new_n671), .A4(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n322), .A3(new_n680), .A4(new_n632), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(new_n687), .B(KEYINPUT39), .Z(new_n691));
  NOR2_X1   g505(.A1(new_n636), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT40), .ZN(new_n693));
  INV_X1    g507(.A(new_n376), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n444), .B1(new_n694), .B2(new_n374), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n680), .A2(new_n447), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n504), .A2(new_n509), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n629), .A2(new_n631), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n621), .B(G472), .C1(new_n599), .C2(new_n615), .ZN(new_n704));
  NAND2_X1  g518(.A1(G472), .A2(G902), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT102), .Z(new_n707));
  NOR2_X1   g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n702), .B(new_n708), .C1(new_n696), .C2(new_n697), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n693), .A2(new_n699), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n212), .ZN(G45));
  NAND2_X1  g525(.A1(new_n297), .A2(new_n321), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n632), .A3(new_n189), .ZN(new_n713));
  INV_X1    g527(.A(new_n687), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n661), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n713), .A2(new_n651), .A3(new_n680), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OR2_X1    g531(.A1(new_n319), .A2(new_n191), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n315), .A2(new_n316), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT86), .B1(new_n319), .B2(new_n191), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n189), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT104), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n321), .A2(new_n723), .A3(new_n189), .A4(new_n718), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n632), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n642), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n662), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n673), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AND2_X1   g547(.A1(new_n321), .A2(new_n718), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n189), .A3(new_n652), .A4(new_n651), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n680), .A2(new_n632), .A3(new_n445), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n460), .ZN(G21));
  NAND2_X1  g552(.A1(new_n616), .A2(new_n600), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n622), .A3(new_n624), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n626), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n644), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n642), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT105), .B1(new_n695), .B2(new_n650), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n377), .A2(new_n651), .A3(new_n746), .A4(new_n444), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n725), .A2(new_n744), .A3(new_n652), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  AND4_X1   g564(.A1(new_n189), .A2(new_n321), .A3(new_n651), .A4(new_n718), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n680), .A3(new_n715), .A4(new_n742), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NOR2_X1   g567(.A1(new_n700), .A2(new_n447), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n293), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n190), .B(new_n755), .C1(new_n321), .C2(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(new_n632), .A3(new_n572), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n661), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n627), .B(KEYINPUT32), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n619), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n757), .A2(new_n572), .A3(new_n715), .A4(new_n761), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n758), .A2(new_n759), .B1(new_n762), .B2(KEYINPUT42), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NOR2_X1   g578(.A1(new_n672), .A2(new_n714), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n727), .A2(new_n765), .A3(new_n757), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  XNOR2_X1  g581(.A(new_n291), .B(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(G469), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n191), .A2(new_n292), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n321), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(KEYINPUT106), .B(new_n321), .C1(new_n772), .C2(new_n773), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n775), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n189), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n691), .ZN(new_n783));
  INV_X1    g597(.A(new_n444), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n660), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n645), .A4(new_n680), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT108), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n645), .A3(new_n680), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n755), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n783), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT109), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  NAND2_X1  g609(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n726), .A2(new_n642), .A3(new_n715), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n781), .A2(new_n798), .A3(new_n189), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n754), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  AND3_X1   g615(.A1(new_n744), .A2(new_n787), .A3(new_n450), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n796), .A2(new_n799), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n734), .A2(new_n190), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n754), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n721), .A2(new_n449), .A3(new_n755), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n787), .A3(new_n680), .A4(new_n742), .ZN(new_n807));
  INV_X1    g621(.A(new_n708), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n642), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n444), .A3(new_n660), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n721), .A2(new_n446), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n701), .B1(new_n813), .B2(KEYINPUT116), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n802), .B(new_n814), .C1(KEYINPUT116), .C2(new_n813), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n812), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n805), .A2(new_n807), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  OAI211_X1 g637(.A(G952), .B(new_n398), .C1(new_n811), .C2(new_n661), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n806), .A2(new_n787), .A3(new_n572), .A4(new_n761), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT48), .Z(new_n826));
  OR2_X1    g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n822), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n802), .A2(new_n751), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n725), .B(new_n727), .C1(new_n662), .C2(new_n673), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n749), .ZN(new_n831));
  INV_X1    g645(.A(new_n645), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n572), .A2(new_n322), .A3(new_n510), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n369), .A2(new_n373), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n784), .A2(new_n834), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n833), .A2(new_n835), .B1(new_n735), .B2(new_n736), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n682), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n833), .A2(new_n661), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT110), .B1(new_n838), .B2(new_n634), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  OAI221_X1 g654(.A(new_n840), .B1(new_n511), .B2(new_n633), .C1(new_n661), .C2(new_n833), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n831), .A2(new_n837), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n757), .A2(new_n680), .A3(new_n715), .A4(new_n742), .ZN(new_n843));
  INV_X1    g657(.A(new_n834), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n844), .A2(new_n671), .A3(new_n687), .A4(new_n754), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n322), .A2(new_n680), .A3(new_n632), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n766), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n763), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n842), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n680), .A2(new_n714), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n190), .B1(new_n321), .B2(new_n756), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n808), .A3(new_n748), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n716), .A2(new_n855), .A3(new_n689), .A4(new_n752), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT52), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n748), .A2(new_n854), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n708), .A2(new_n680), .A3(new_n714), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n752), .A2(KEYINPUT112), .A3(new_n689), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT112), .B1(new_n752), .B2(new_n689), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n716), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n865), .A2(KEYINPUT114), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT114), .B1(new_n865), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n851), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n858), .A2(new_n872), .A3(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n867), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(KEYINPUT114), .A3(new_n867), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n851), .A2(KEYINPUT53), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n871), .B1(new_n852), .B2(new_n857), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT53), .A4(new_n851), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n879), .A2(new_n880), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n828), .A2(new_n829), .A3(new_n873), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n785), .A2(new_n701), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT49), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n887), .B1(new_n734), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n888), .B2(new_n734), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n189), .A3(new_n446), .A4(new_n809), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(G75));
  OR2_X1    g706(.A1(new_n398), .A2(G952), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT119), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(G210), .A3(G902), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n486), .B1(new_n480), .B2(new_n487), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n508), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n895), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n896), .A2(KEYINPUT117), .A3(G210), .A4(G902), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n903), .A2(new_n909), .ZN(G51));
  NAND2_X1  g724(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n884), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n770), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n318), .A2(new_n313), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n896), .A2(G902), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(G469), .A3(new_n768), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n895), .B1(new_n917), .B2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n436), .A2(new_n422), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n922), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n895), .B1(new_n923), .B2(new_n925), .ZN(G60));
  XNOR2_X1  g740(.A(new_n654), .B(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n884), .B2(new_n873), .ZN(new_n928));
  INV_X1    g742(.A(new_n659), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n894), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n659), .A2(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n912), .B2(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(KEYINPUT121), .ZN(new_n934));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT60), .Z(new_n936));
  NAND3_X1  g750(.A1(new_n896), .A2(new_n678), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n895), .B1(KEYINPUT121), .B2(new_n933), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n568), .B1(new_n896), .B2(new_n936), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  INV_X1    g756(.A(new_n934), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n937), .A4(new_n938), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n941), .A2(new_n944), .ZN(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n452), .B2(new_n484), .ZN(new_n946));
  INV_X1    g760(.A(new_n842), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n480), .A2(new_n487), .B1(G898), .B2(new_n398), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  OR2_X1    g764(.A1(new_n863), .A2(new_n864), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n716), .ZN(new_n952));
  AND2_X1   g766(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n952), .A2(new_n710), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n793), .A2(new_n800), .ZN(new_n955));
  NOR2_X1   g769(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n956));
  OAI22_X1  g770(.A1(new_n952), .A2(new_n710), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n835), .A2(new_n661), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n692), .A2(new_n727), .A3(new_n754), .A4(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n954), .A2(new_n955), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n583), .A2(new_n587), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n432), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n951), .A2(new_n716), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n763), .A2(new_n766), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n748), .A2(new_n572), .A3(new_n761), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n783), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n965), .A2(new_n968), .A3(new_n793), .A4(new_n800), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n398), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n970), .B(new_n962), .C1(G900), .C2(new_n398), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n964), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n193), .B2(new_n685), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G72));
  XOR2_X1   g793(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n705), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n969), .B2(new_n842), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n595), .B(KEYINPUT125), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n600), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(new_n894), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n984), .B2(new_n894), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n960), .B2(new_n842), .ZN(new_n989));
  INV_X1    g803(.A(new_n983), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n599), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n601), .A2(new_n621), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n858), .A2(new_n872), .A3(new_n981), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT127), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n984), .A2(new_n894), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT126), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n984), .A2(new_n985), .A3(new_n894), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n999), .A2(new_n1000), .A3(new_n993), .A4(new_n991), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n995), .A2(new_n1001), .ZN(G57));
endmodule


