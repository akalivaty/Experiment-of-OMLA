//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(G77), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT66), .B(G244), .Z(new_n225));
  OAI211_X1 g0025(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G13), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n248), .A2(new_n207), .A3(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n207), .A2(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(KEYINPUT74), .B2(new_n256), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(KEYINPUT74), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n257), .A2(new_n258), .B1(new_n254), .B2(new_n249), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n219), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n262), .B2(new_n201), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G159), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT68), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n207), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n275), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n268), .A2(new_n269), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT73), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n277), .A2(new_n279), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n267), .B1(new_n285), .B2(new_n219), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT16), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n251), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n279), .A2(new_n207), .A3(new_n282), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n274), .A2(new_n207), .A3(new_n275), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n219), .B1(new_n291), .B2(KEYINPUT7), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n266), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n289), .B1(new_n293), .B2(KEYINPUT16), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n260), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(G1), .A2(G13), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n274), .A2(new_n275), .ZN(new_n299));
  INV_X1    g0099(.A(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G1698), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n299), .B(new_n301), .C1(G223), .C2(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G87), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT75), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n298), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  AOI21_X1  g0108(.A(G1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n298), .A2(G274), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n298), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G232), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n305), .A2(new_n306), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n305), .A2(new_n314), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(G169), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT18), .B1(new_n295), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n275), .ZN(new_n322));
  AOI21_X1  g0122(.A(G20), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n319), .A2(new_n320), .B1(new_n323), .B2(new_n278), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n266), .B1(new_n324), .B2(G68), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n294), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n317), .B1(new_n326), .B2(new_n259), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n305), .B2(new_n314), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n316), .B2(G190), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n259), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n318), .B(new_n329), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n224), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G20), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n207), .A2(G33), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  INV_X1    g0143(.A(new_n264), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n341), .B1(new_n342), .B2(new_n343), .C1(new_n254), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(new_n251), .ZN(new_n346));
  INV_X1    g0146(.A(G77), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n255), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n252), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n248), .A2(G1), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G20), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n340), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n310), .B1(new_n312), .B2(new_n225), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n271), .A2(new_n276), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(G232), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(G238), .A3(G1698), .ZN(new_n358));
  INV_X1    g0158(.A(G107), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n355), .ZN(new_n360));
  INV_X1    g0160(.A(new_n298), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n353), .B1(new_n362), .B2(G190), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n361), .ZN(new_n364));
  INV_X1    g0164(.A(new_n354), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G200), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n346), .A2(new_n352), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(new_n306), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n339), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n321), .A2(new_n322), .A3(G232), .A4(G1698), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n321), .A2(new_n322), .A3(G226), .A4(new_n356), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G97), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n361), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n310), .B1(new_n312), .B2(new_n220), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT13), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n379), .B2(new_n361), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT13), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT71), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n249), .A2(new_n219), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT12), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n347), .B2(new_n342), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n396));
  INV_X1    g0196(.A(new_n255), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n252), .A2(G68), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT11), .B1(new_n395), .B2(new_n251), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n387), .B1(new_n380), .B2(new_n382), .ZN(new_n402));
  AOI211_X1 g0202(.A(KEYINPUT13), .B(new_n381), .C1(new_n379), .C2(new_n361), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n391), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G169), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT14), .B(G169), .C1(new_n402), .C2(new_n403), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n385), .A2(new_n388), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n403), .A2(new_n306), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n405), .B1(new_n412), .B2(new_n401), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n255), .A2(new_n202), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n252), .A2(new_n415), .B1(new_n202), .B2(new_n249), .ZN(new_n416));
  INV_X1    g0216(.A(G150), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n254), .A2(new_n342), .B1(new_n417), .B2(new_n344), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(G20), .B2(new_n203), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(new_n289), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT9), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT9), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(new_n416), .C1(new_n419), .C2(new_n289), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n424), .A2(KEYINPUT69), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT10), .B1(new_n424), .B2(KEYINPUT69), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n310), .B1(new_n312), .B2(new_n300), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n355), .A2(G222), .A3(new_n356), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n355), .A2(G223), .A3(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n429), .C1(new_n224), .C2(new_n355), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n430), .B2(new_n361), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n361), .ZN(new_n434));
  INV_X1    g0234(.A(new_n427), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(G190), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n425), .A2(new_n426), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n424), .C1(new_n330), .C2(new_n431), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT70), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT10), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n438), .B2(KEYINPUT10), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n306), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n420), .C1(G169), .C2(new_n431), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n375), .A2(new_n414), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G87), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n447), .A2(KEYINPUT22), .A3(G20), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n321), .A2(new_n322), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT83), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT83), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n321), .A2(new_n322), .A3(new_n451), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(new_n274), .B2(new_n275), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G87), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n359), .A2(KEYINPUT23), .A3(G20), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT23), .B1(new_n359), .B2(G20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G116), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n460), .A2(new_n461), .B1(G20), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(KEYINPUT24), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n456), .B1(new_n450), .B2(new_n452), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(new_n463), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n251), .A3(new_n468), .ZN(new_n469));
  OR3_X1    g0269(.A1(new_n351), .A2(KEYINPUT25), .A3(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT25), .B1(new_n351), .B2(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n273), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n289), .A2(new_n351), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n470), .B(new_n471), .C1(new_n359), .C2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n308), .A2(G1), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(new_n298), .A3(G274), .A4(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n478), .B2(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G264), .A3(new_n298), .ZN(new_n484));
  NOR2_X1   g0284(.A1(G250), .A2(G1698), .ZN(new_n485));
  INV_X1    g0285(.A(G257), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(G1698), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n299), .B1(G33), .B2(G294), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n482), .B(new_n484), .C1(new_n488), .C2(new_n298), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n370), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(G179), .B2(new_n489), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT85), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n494), .B(new_n491), .C1(new_n469), .C2(new_n476), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n489), .A2(new_n330), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G190), .B2(new_n489), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n469), .A2(new_n476), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n281), .A2(new_n284), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n321), .A2(new_n322), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n278), .B1(new_n502), .B2(new_n207), .ZN(new_n503));
  OAI21_X1  g0303(.A(G107), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n505), .A2(new_n506), .A3(G107), .ZN(new_n507));
  XNOR2_X1  g0307(.A(G97), .B(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n509), .A2(new_n207), .B1(new_n347), .B2(new_n344), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n289), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n351), .A2(G97), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n249), .A2(new_n251), .A3(new_n472), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(G97), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT77), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n356), .C1(new_n268), .C2(new_n269), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n518), .A2(new_n519), .B1(G33), .B2(G283), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n321), .A2(new_n322), .A3(G250), .A4(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G244), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n321), .A2(new_n322), .A3(new_n356), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n361), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n483), .A2(new_n298), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n482), .B1(new_n527), .B2(new_n486), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n525), .B2(new_n361), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G179), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n510), .B1(new_n324), .B2(G107), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n515), .C1(new_n536), .C2(new_n289), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n517), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n511), .B1(new_n285), .B2(new_n359), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n516), .B1(new_n539), .B2(new_n251), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n532), .A2(G190), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n330), .C2(new_n532), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  INV_X1    g0344(.A(G270), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n482), .B1(new_n527), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(G303), .B1(new_n271), .B2(new_n276), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n299), .A2(G264), .A3(G1698), .ZN(new_n548));
  OAI211_X1 g0348(.A(G257), .B(new_n356), .C1(new_n268), .C2(new_n269), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n299), .A2(KEYINPUT81), .A3(G257), .A4(new_n356), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(new_n548), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n546), .B1(new_n553), .B2(new_n361), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n250), .A2(new_n215), .B1(G20), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(G20), .B1(G33), .B2(G283), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G33), .B2(new_n506), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT20), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT20), .B1(new_n556), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n249), .A2(G116), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n474), .B2(G116), .ZN(new_n563));
  OAI21_X1  g0363(.A(G169), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n544), .B1(new_n554), .B2(new_n564), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n306), .B(new_n546), .C1(new_n553), .C2(new_n361), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n561), .A2(new_n563), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n565), .A2(KEYINPUT21), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G250), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n296), .B2(new_n297), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT79), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n206), .A2(KEYINPUT78), .A3(G45), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT78), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n308), .B2(G1), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n298), .A2(G274), .A3(new_n481), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n220), .A2(new_n356), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n522), .A2(G1698), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n268), .C2(new_n269), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n298), .B1(new_n581), .B2(new_n462), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n575), .A2(new_n573), .ZN(new_n584));
  AND2_X1   g0384(.A1(G33), .A2(G41), .ZN(new_n585));
  OAI21_X1  g0385(.A(G250), .B1(new_n585), .B2(new_n215), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT79), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n578), .A2(new_n306), .A3(new_n583), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n577), .A3(new_n576), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n370), .B1(new_n589), .B2(new_n582), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n207), .B1(new_n378), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n447), .A2(new_n506), .A3(new_n359), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n207), .B(G68), .C1(new_n268), .C2(new_n269), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n342), .B2(new_n506), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n251), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n343), .A2(new_n249), .ZN(new_n600));
  INV_X1    g0400(.A(new_n343), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n514), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n598), .A2(new_n251), .B1(new_n249), .B2(new_n343), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT80), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n514), .A2(G87), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n599), .A2(new_n600), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n589), .A2(new_n582), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(G190), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n589), .B2(new_n582), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n591), .A2(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT21), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n544), .B(new_n615), .C1(new_n554), .C2(new_n564), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n554), .A2(G190), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n567), .C1(new_n330), .C2(new_n554), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n569), .A2(new_n614), .A3(new_n616), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n543), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n446), .A2(new_n500), .A3(new_n620), .ZN(G372));
  NAND3_X1  g0421(.A1(new_n295), .A2(new_n332), .A3(new_n336), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n333), .A2(new_n334), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n371), .A2(new_n372), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n625), .A2(new_n405), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n412), .A2(new_n401), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n318), .A2(new_n329), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n442), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n444), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n582), .A2(KEYINPUT86), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT86), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n635), .B(new_n298), .C1(new_n581), .C2(new_n462), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n587), .B(new_n578), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n370), .B1(new_n306), .B2(new_n611), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(G200), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n608), .B1(new_n612), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n499), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT87), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(new_n538), .A4(new_n542), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n538), .A2(new_n499), .A3(new_n542), .A4(new_n640), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n569), .A2(new_n616), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n491), .B1(new_n469), .B2(new_n476), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n614), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT26), .B1(new_n538), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n515), .B1(new_n536), .B2(new_n289), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n640), .A2(new_n652), .A3(new_n653), .A4(new_n534), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n638), .A2(KEYINPUT88), .A3(new_n608), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT88), .B1(new_n638), .B2(new_n608), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n651), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n446), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n633), .A2(new_n661), .ZN(G369));
  NAND2_X1  g0462(.A1(new_n350), .A2(new_n207), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT89), .ZN(new_n665));
  INV_X1    g0465(.A(G213), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n663), .B2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n477), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n500), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n647), .A2(new_n671), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n646), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n677), .B(new_n618), .C1(new_n567), .C2(new_n670), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n646), .A2(new_n568), .A3(new_n671), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n677), .A2(new_n671), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n500), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n647), .A2(new_n670), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n210), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n594), .A2(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n213), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n644), .B1(new_n496), .B2(new_n677), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n653), .A2(KEYINPUT77), .B1(new_n531), .B2(new_n533), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n652), .A3(new_n537), .A4(new_n614), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n639), .A2(new_n612), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n583), .A2(new_n635), .ZN(new_n701));
  INV_X1    g0501(.A(new_n636), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n589), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n588), .B1(new_n703), .B2(G169), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n606), .B1(new_n605), .B2(new_n602), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n700), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n530), .A2(new_n306), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n532), .A2(new_n370), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n653), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT26), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT88), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n704), .B2(new_n707), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n655), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(new_n714), .B2(new_n655), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n699), .B(new_n712), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n696), .B(new_n670), .C1(new_n697), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT90), .B1(new_n656), .B2(new_n657), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n716), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n712), .A2(new_n699), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n493), .A2(new_n495), .A3(new_n646), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n644), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n696), .B1(new_n726), .B2(new_n670), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT29), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n671), .B1(new_n649), .B2(new_n659), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(KEYINPUT29), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n620), .A2(new_n496), .A3(new_n499), .A4(new_n670), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n484), .B1(new_n488), .B2(new_n298), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n732), .A2(new_n589), .A3(new_n582), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n554), .A3(new_n532), .A4(G179), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n566), .A2(KEYINPUT30), .A3(new_n532), .A4(new_n733), .ZN(new_n737));
  INV_X1    g0537(.A(new_n554), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n489), .A2(new_n306), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n530), .A3(new_n637), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n741), .B2(new_n671), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n730), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n695), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n248), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n690), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n215), .B1(G20), .B2(new_n370), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n306), .A2(new_n330), .A3(G190), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n506), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n207), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n355), .B1(new_n447), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(new_n389), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n759), .B(new_n762), .C1(G107), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n766), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n771), .A2(new_n389), .A3(G200), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n774), .A2(new_n340), .B1(G58), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(new_n389), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n771), .A2(new_n389), .A3(new_n330), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n778), .A2(G68), .B1(new_n779), .B2(G50), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n765), .A2(new_n770), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G317), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n778), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  INV_X1    g0586(.A(new_n775), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n767), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G329), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n763), .B1(new_n761), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G294), .B2(new_n757), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n774), .A2(G311), .B1(new_n779), .B2(G326), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n790), .A2(new_n502), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n755), .B1(new_n781), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n754), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n355), .A2(G355), .A3(new_n210), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n689), .A2(new_n299), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n213), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n246), .A2(new_n308), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n802), .B1(G116), .B2(new_n210), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n753), .B(new_n797), .C1(new_n801), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT92), .ZN(new_n808));
  INV_X1    g0608(.A(new_n800), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n680), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n680), .A2(G330), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n681), .A2(new_n753), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n660), .A2(new_n670), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n625), .A2(new_n670), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n363), .A2(new_n367), .B1(new_n353), .B2(new_n671), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n625), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n660), .A2(new_n670), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n752), .B1(new_n823), .B2(new_n746), .ZN(new_n824));
  INV_X1    g0624(.A(G330), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n731), .B2(new_n744), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n820), .A2(new_n826), .A3(new_n822), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G137), .A2(new_n779), .B1(new_n775), .B2(G143), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n417), .B2(new_n777), .C1(new_n768), .C2(new_n773), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n763), .A2(new_n219), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n282), .B(new_n834), .C1(G132), .C2(new_n789), .ZN(new_n835));
  INV_X1    g0635(.A(new_n761), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G50), .B1(new_n757), .B2(G58), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n763), .A2(new_n447), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n839), .B(new_n759), .C1(G107), .C2(new_n836), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n777), .A2(new_n791), .B1(new_n767), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G303), .B2(new_n779), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n774), .A2(G116), .B1(G294), .B2(new_n775), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n502), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n755), .B1(new_n838), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n754), .A2(new_n798), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n753), .B1(new_n347), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n846), .B(new_n849), .C1(new_n819), .C2(new_n798), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n828), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n749), .A2(new_n206), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT97), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT29), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n670), .B1(new_n697), .B2(new_n719), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT91), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(new_n720), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n446), .B1(KEYINPUT29), .B2(new_n729), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n445), .B1(new_n816), .B2(new_n855), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n728), .A2(new_n861), .A3(KEYINPUT97), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n632), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT98), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n326), .A2(new_n259), .A3(new_n332), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n327), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  AOI211_X1 g0667(.A(KEYINPUT95), .B(new_n668), .C1(new_n326), .C2(new_n259), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT95), .ZN(new_n869));
  OAI21_X1  g0669(.A(G68), .B1(new_n501), .B2(new_n503), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT16), .B1(new_n870), .B2(new_n267), .ZN(new_n871));
  INV_X1    g0671(.A(new_n294), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n259), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n873), .B2(new_n669), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n317), .A2(new_n668), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n293), .A2(KEYINPUT16), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n259), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n867), .B1(new_n879), .B2(new_n333), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n669), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n622), .A2(new_n623), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n318), .A2(new_n329), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n868), .A2(new_n874), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n333), .B1(new_n295), .B2(new_n317), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(new_n875), .B1(new_n339), .B2(new_n890), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n888), .B(new_n889), .C1(new_n893), .C2(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(KEYINPUT96), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n873), .A2(new_n869), .A3(new_n669), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT95), .B1(new_n295), .B2(new_n668), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n891), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n880), .B1(new_n900), .B2(new_n867), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n883), .B1(new_n629), .B2(new_n624), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT96), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n882), .A2(new_n904), .A3(new_n887), .A4(KEYINPUT38), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n896), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n895), .B1(KEYINPUT39), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n627), .A2(new_n670), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n408), .A2(new_n409), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n410), .A2(new_n411), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n405), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n670), .A2(new_n401), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT94), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n913), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n405), .B(new_n917), .C1(new_n412), .C2(new_n401), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(KEYINPUT94), .A3(new_n913), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n822), .B2(new_n817), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n906), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n629), .B2(new_n669), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n909), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n864), .B(new_n925), .Z(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n920), .A2(new_n745), .A3(new_n821), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n906), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n893), .A2(KEYINPUT38), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n932), .B2(new_n888), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n929), .A2(new_n930), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n446), .A2(new_n745), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n446), .A3(new_n745), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(G330), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n853), .B1(new_n927), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n927), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(new_n509), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(G116), .A3(new_n216), .A4(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT36), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n224), .A2(new_n213), .A3(new_n262), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n219), .A2(G50), .ZN(new_n948));
  OAI211_X1 g0748(.A(G1), .B(new_n248), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n946), .A3(new_n949), .ZN(G367));
  INV_X1    g0750(.A(new_n803), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n801), .B1(new_n210), .B2(new_n343), .C1(new_n951), .C2(new_n239), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n752), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n671), .A2(new_n610), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n640), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n658), .B2(new_n954), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n787), .A2(new_n792), .B1(new_n767), .B2(new_n782), .ZN(new_n957));
  INV_X1    g0757(.A(G294), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n282), .B1(new_n777), .B2(new_n958), .C1(new_n506), .C2(new_n763), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n957), .B(new_n959), .C1(G311), .C2(new_n779), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n836), .A2(G116), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT46), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n758), .A2(new_n359), .B1(new_n773), .B2(new_n791), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT105), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n757), .A2(G68), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n417), .B2(new_n787), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT106), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(G143), .ZN(new_n971));
  INV_X1    g0771(.A(new_n779), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n969), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT107), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n777), .A2(new_n768), .B1(new_n773), .B2(new_n202), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT108), .Z(new_n976));
  INV_X1    g0776(.A(G137), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n355), .B1(new_n977), .B2(new_n767), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n261), .A2(new_n761), .B1(new_n763), .B2(new_n224), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n973), .A2(KEYINPUT107), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n965), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT47), .Z(new_n984));
  OAI221_X1 g0784(.A(new_n953), .B1(new_n809), .B2(new_n956), .C1(new_n984), .C2(new_n755), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n711), .A2(new_n670), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT100), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n538), .B(new_n542), .C1(new_n540), .C2(new_n670), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n685), .A2(new_n686), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT45), .Z(new_n991));
  INV_X1    g0791(.A(KEYINPUT102), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n989), .B1(new_n685), .B2(new_n686), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n993), .B2(new_n995), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n992), .B(new_n994), .C1(new_n687), .C2(new_n989), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n991), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n682), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT103), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n682), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n685), .B1(new_n675), .B2(new_n684), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(new_n681), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n747), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n747), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT104), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n690), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n747), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT104), .B1(new_n1014), .B2(new_n1010), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n751), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n989), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n685), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n538), .B1(new_n1017), .B2(new_n496), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(KEYINPUT42), .B1(new_n1021), .B2(new_n670), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1020), .A2(new_n1022), .B1(KEYINPUT43), .B2(new_n956), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n683), .A2(new_n1017), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n985), .B1(new_n1016), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(G387));
  INV_X1    g0830(.A(new_n692), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n355), .A2(new_n210), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(G107), .B2(new_n210), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n236), .A2(new_n308), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(G45), .B(new_n1031), .C1(G68), .C2(G77), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n254), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n951), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1033), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT111), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n801), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n774), .A2(G68), .B1(G50), .B2(new_n775), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n417), .B2(new_n767), .C1(new_n768), .C2(new_n972), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n299), .B1(new_n777), .B2(new_n254), .C1(new_n506), .C2(new_n763), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n758), .A2(new_n343), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n761), .A2(new_n224), .ZN(new_n1049));
  NOR4_X1   g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n836), .A2(G294), .B1(new_n757), .B2(G283), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G322), .A2(new_n779), .B1(new_n775), .B2(G317), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n792), .B2(new_n773), .C1(new_n841), .C2(new_n777), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT49), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n763), .A2(new_n555), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n299), .B(new_n1060), .C1(G326), .C2(new_n789), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1050), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n752), .B1(new_n1043), .B2(new_n1044), .C1(new_n1062), .C2(new_n755), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT113), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n676), .B2(new_n800), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1004), .B2(new_n751), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1005), .A2(new_n690), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n747), .A2(new_n1004), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  AND2_X1   g0869(.A1(new_n999), .A2(new_n682), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(new_n1002), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n691), .B1(new_n1071), .B2(new_n1005), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1007), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1071), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1017), .A2(new_n800), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n801), .B1(new_n506), .B2(new_n210), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n803), .B2(new_n243), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G150), .A2(new_n779), .B1(new_n775), .B2(G159), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n761), .A2(new_n219), .B1(new_n767), .B2(new_n971), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT114), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n299), .B1(new_n773), .B2(new_n254), .C1(new_n202), .C2(new_n777), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n758), .A2(new_n347), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1082), .A2(new_n839), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G317), .A2(new_n779), .B1(new_n775), .B2(G311), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  AOI22_X1  g0887(.A1(new_n778), .A2(G303), .B1(new_n774), .B2(G294), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n764), .A2(G107), .B1(new_n757), .B2(G116), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1087), .A2(new_n502), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n761), .A2(new_n791), .B1(new_n767), .B2(new_n786), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT115), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1085), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n753), .B(new_n1077), .C1(new_n1093), .C2(new_n754), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1074), .A2(new_n751), .B1(new_n1075), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1073), .A2(new_n1095), .ZN(G390));
  NAND2_X1  g0896(.A1(new_n446), .A2(new_n826), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n858), .A2(new_n859), .A3(new_n854), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT97), .B1(new_n728), .B2(new_n861), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n633), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n921), .B1(new_n746), .B2(new_n819), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n825), .B(new_n819), .C1(new_n731), .C2(new_n744), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n920), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n826), .A2(new_n920), .A3(new_n1102), .A4(new_n821), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1101), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n818), .A2(new_n625), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n729), .A2(new_n1109), .B1(new_n625), .B2(new_n670), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n826), .A2(new_n821), .A3(new_n920), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n857), .A2(new_n720), .A3(new_n817), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1109), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1107), .A2(new_n1111), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1100), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT118), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1109), .A3(new_n920), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n908), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n932), .B2(new_n888), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n903), .A2(new_n905), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n881), .A2(new_n875), .B1(new_n339), .B2(new_n884), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n904), .B1(new_n1124), .B2(KEYINPUT38), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT39), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n894), .C1(new_n922), .C2(new_n1120), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1122), .A2(new_n1127), .A3(new_n1112), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n908), .B1(new_n1110), .B2(new_n921), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n907), .A2(new_n1129), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1112), .A2(KEYINPUT116), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1105), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1128), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1118), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1122), .A2(new_n1127), .A3(new_n1112), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1132), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT117), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1117), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n920), .B1(new_n826), .B2(new_n821), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1131), .B2(new_n1105), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n721), .A2(new_n727), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1108), .B1(new_n1142), .B2(new_n817), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1141), .A2(new_n1110), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n863), .A3(new_n1097), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT117), .B1(new_n1133), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1139), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1134), .A2(new_n690), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1137), .A2(new_n751), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n907), .A2(new_n798), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n753), .B1(new_n254), .B2(new_n847), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n834), .B(new_n1083), .C1(G87), .C2(new_n836), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n787), .A2(new_n555), .B1(new_n767), .B2(new_n958), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G283), .B2(new_n779), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n778), .A2(G107), .B1(new_n774), .B2(G97), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n502), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G132), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n787), .A2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n502), .B(new_n1159), .C1(G125), .C2(new_n789), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n761), .A2(new_n417), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n972), .A2(new_n1163), .B1(new_n777), .B2(new_n977), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n774), .B2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n764), .A2(G50), .B1(new_n757), .B2(G159), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1160), .A2(new_n1162), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1151), .B(new_n1152), .C1(new_n755), .C2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1149), .A2(new_n1150), .A3(new_n1171), .ZN(G378));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n925), .B1(new_n825), .B2(new_n935), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n934), .B(G330), .C1(new_n909), .C2(new_n924), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n442), .A2(new_n444), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n669), .A2(new_n420), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT55), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1178), .B(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1176), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1177), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1174), .A2(new_n1185), .A3(new_n1175), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1173), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1100), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT122), .B1(new_n1148), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT122), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1190), .B(new_n1100), .C1(new_n1139), .C2(new_n1147), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1187), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1176), .B(new_n1185), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1138), .B1(new_n1137), .B2(new_n1117), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1133), .A2(new_n1146), .A3(KEYINPUT117), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1190), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1148), .A2(KEYINPUT122), .A3(new_n1188), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1193), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n690), .B(new_n1192), .C1(new_n1199), .C2(KEYINPUT57), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT123), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1183), .A2(new_n799), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n847), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n752), .B1(G50), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n282), .B2(new_n307), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n972), .A2(new_n555), .B1(new_n777), .B2(new_n506), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n787), .A2(new_n359), .B1(new_n767), .B2(new_n791), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G41), .B(new_n299), .C1(new_n774), .C2(new_n601), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1049), .B1(G58), .B2(new_n764), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n966), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n774), .A2(G137), .B1(new_n779), .B2(G125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1158), .B2(new_n777), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n787), .A2(new_n1163), .B1(new_n761), .B2(new_n1165), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT119), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G150), .C2(new_n757), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT59), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1216), .B1(new_n768), .B2(new_n763), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1215), .B1(new_n1214), .B2(new_n1213), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1205), .B1(new_n1225), .B2(new_n754), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1202), .A2(new_n751), .B1(new_n1203), .B2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1200), .A2(new_n1201), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1201), .B1(new_n1200), .B2(new_n1227), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1100), .A2(new_n1116), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1118), .A2(new_n1011), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT124), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n921), .B2(new_n798), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n920), .A2(KEYINPUT124), .A3(new_n799), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1048), .B1(G97), .B2(new_n836), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n347), .B2(new_n763), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n502), .B1(new_n359), .B2(new_n773), .C1(new_n792), .C2(new_n767), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n778), .A2(G116), .B1(new_n779), .B2(G294), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n791), .B2(new_n787), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n299), .B1(new_n773), .B2(new_n417), .C1(new_n763), .C2(new_n261), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n758), .A2(new_n202), .B1(new_n761), .B2(new_n768), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n972), .A2(new_n1158), .B1(new_n777), .B2(new_n1165), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n787), .A2(new_n977), .B1(new_n767), .B2(new_n1163), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n754), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n752), .C1(G68), .C2(new_n1204), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT125), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1234), .A2(new_n1235), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1145), .B2(new_n751), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1232), .A2(new_n1251), .ZN(G381));
  OAI211_X1 g1052(.A(new_n1066), .B(new_n814), .C1(new_n1068), .C2(new_n1067), .ZN(new_n1253));
  OR4_X1    g1053(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1253), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1254), .ZN(G407));
  NAND2_X1  g1055(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1256), .B2(new_n1202), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1192), .A2(new_n690), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1227), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT123), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1200), .A2(new_n1201), .A3(new_n1227), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G378), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n666), .A2(G343), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(new_n1264), .A3(G213), .ZN(G409));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1227), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1011), .B(new_n1202), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1203), .A2(new_n1226), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1202), .A2(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n751), .B1(new_n1193), .B2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1268), .B(new_n1269), .C1(new_n1270), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G378), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1267), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1263), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1231), .B1(new_n1117), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1100), .A2(new_n1116), .A3(KEYINPUT60), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n690), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1251), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n851), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1283), .A2(new_n851), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1266), .B1(new_n1278), .B2(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1263), .A2(G2897), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1287), .B(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1253), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1029), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1073), .A2(new_n1095), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1073), .A2(new_n1095), .B1(new_n1298), .B2(new_n1253), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1301), .B(new_n985), .C1(new_n1016), .C2(new_n1027), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1296), .B2(new_n1295), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1028), .A2(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1263), .B1(new_n1267), .B2(new_n1275), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1289), .A2(new_n1292), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1306), .A2(new_n1309), .A3(new_n1287), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1291), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1311), .B1(new_n1306), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1309), .B1(new_n1306), .B2(new_n1287), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1310), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1308), .B1(new_n1315), .B2(new_n1305), .ZN(G405));
  NAND2_X1  g1116(.A1(new_n1259), .A2(G378), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT127), .B1(new_n1262), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1274), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1317), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1302), .A2(new_n1288), .A3(new_n1304), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1288), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1319), .A2(new_n1322), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1319), .B2(new_n1322), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


