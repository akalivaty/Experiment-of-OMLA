

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(n955), .ZN(n780) );
  AND2_X1 U550 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U551 ( .A1(n595), .A2(G1384), .ZN(n710) );
  XNOR2_X2 U552 ( .A(G2104), .B(KEYINPUT65), .ZN(n570) );
  BUF_X1 U553 ( .A(n633), .Z(n647) );
  NOR2_X1 U554 ( .A1(n627), .A2(n626), .ZN(n632) );
  INV_X1 U555 ( .A(KEYINPUT97), .ZN(n674) );
  NOR2_X1 U556 ( .A1(n687), .A2(n689), .ZN(n690) );
  OR2_X1 U557 ( .A1(n696), .A2(n695), .ZN(n516) );
  BUF_X1 U558 ( .A(n652), .Z(n633) );
  INV_X1 U559 ( .A(KEYINPUT30), .ZN(n657) );
  INV_X1 U560 ( .A(KEYINPUT29), .ZN(n645) );
  INV_X1 U561 ( .A(KEYINPUT31), .ZN(n663) );
  AND2_X1 U562 ( .A1(n653), .A2(n652), .ZN(n654) );
  INV_X1 U563 ( .A(n961), .ZN(n689) );
  INV_X1 U564 ( .A(n949), .ZN(n695) );
  NAND2_X1 U565 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U566 ( .A(KEYINPUT101), .ZN(n748) );
  NOR2_X1 U567 ( .A1(G651), .A2(n554), .ZN(n600) );
  XNOR2_X1 U568 ( .A(n586), .B(KEYINPUT23), .ZN(n587) );
  XNOR2_X1 U569 ( .A(n749), .B(n748), .ZN(n763) );
  XNOR2_X1 U570 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n764) );
  XOR2_X1 U571 ( .A(KEYINPUT71), .B(n535), .Z(G301) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U573 ( .A1(G91), .A2(n793), .ZN(n518) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n554) );
  INV_X1 U575 ( .A(G651), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n554), .A2(n519), .ZN(n797) );
  NAND2_X1 U577 ( .A1(G78), .A2(n797), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n518), .A2(n517), .ZN(n523) );
  NOR2_X1 U579 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n520), .Z(n597) );
  BUF_X1 U581 ( .A(n597), .Z(n794) );
  NAND2_X1 U582 ( .A1(G65), .A2(n794), .ZN(n521) );
  XNOR2_X1 U583 ( .A(KEYINPUT73), .B(n521), .ZN(n522) );
  NOR2_X1 U584 ( .A1(n523), .A2(n522), .ZN(n525) );
  BUF_X1 U585 ( .A(n600), .Z(n798) );
  NAND2_X1 U586 ( .A1(n798), .A2(G53), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(G299) );
  NAND2_X1 U588 ( .A1(G64), .A2(n794), .ZN(n527) );
  NAND2_X1 U589 ( .A1(G52), .A2(n798), .ZN(n526) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT69), .ZN(n534) );
  XNOR2_X1 U592 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n532) );
  NAND2_X1 U593 ( .A1(G90), .A2(n793), .ZN(n530) );
  NAND2_X1 U594 ( .A1(G77), .A2(n797), .ZN(n529) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X1 U598 ( .A(G301), .ZN(G171) );
  NAND2_X1 U599 ( .A1(n793), .A2(G89), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT4), .ZN(n538) );
  NAND2_X1 U601 ( .A1(G76), .A2(n797), .ZN(n537) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT5), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G63), .A2(n794), .ZN(n541) );
  NAND2_X1 U605 ( .A1(G51), .A2(n798), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G88), .A2(n793), .ZN(n547) );
  NAND2_X1 U612 ( .A1(G62), .A2(n794), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U614 ( .A1(G50), .A2(n798), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT83), .B(n548), .ZN(n549) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n797), .A2(G75), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(G303) );
  NAND2_X1 U619 ( .A1(G74), .A2(G651), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT80), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G49), .A2(n798), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G87), .A2(n554), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U624 ( .A1(n794), .A2(n557), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(G288) );
  NAND2_X1 U626 ( .A1(G48), .A2(n798), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT82), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n797), .A2(G73), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT2), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G61), .A2(n794), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G86), .A2(n793), .ZN(n564) );
  XNOR2_X1 U633 ( .A(KEYINPUT81), .B(n564), .ZN(n565) );
  NOR2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(G305) );
  AND2_X2 U636 ( .A1(n570), .A2(G2105), .ZN(n890) );
  NAND2_X1 U637 ( .A1(G126), .A2(n890), .ZN(n569) );
  XNOR2_X1 U638 ( .A(KEYINPUT87), .B(n569), .ZN(n577) );
  NOR2_X2 U639 ( .A1(G2105), .A2(n570), .ZN(n585) );
  NAND2_X1 U640 ( .A1(G102), .A2(n585), .ZN(n572) );
  AND2_X1 U641 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U642 ( .A1(G114), .A2(n891), .ZN(n571) );
  AND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n575) );
  NOR2_X1 U644 ( .A1(G2105), .A2(G2104), .ZN(n573) );
  XOR2_X1 U645 ( .A(KEYINPUT17), .B(n573), .Z(n588) );
  NAND2_X1 U646 ( .A1(n588), .A2(G138), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n595) );
  BUF_X1 U649 ( .A(n595), .Z(G164) );
  NAND2_X1 U650 ( .A1(G85), .A2(n793), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G72), .A2(n797), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U653 ( .A(KEYINPUT68), .B(n580), .Z(n584) );
  NAND2_X1 U654 ( .A1(G60), .A2(n794), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G47), .A2(n798), .ZN(n581) );
  AND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(G290) );
  NAND2_X1 U658 ( .A1(G101), .A2(n585), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT67), .ZN(n590) );
  BUF_X1 U660 ( .A(n588), .Z(n887) );
  NAND2_X1 U661 ( .A1(G137), .A2(n887), .ZN(n589) );
  AND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n767) );
  NAND2_X1 U663 ( .A1(n890), .A2(G125), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT66), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G113), .A2(n891), .ZN(n592) );
  AND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n766) );
  AND2_X1 U667 ( .A1(n766), .A2(G40), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n767), .A2(n594), .ZN(n711) );
  INV_X1 U669 ( .A(n710), .ZN(n596) );
  NOR2_X2 U670 ( .A1(n711), .A2(n596), .ZN(n652) );
  NAND2_X1 U671 ( .A1(n797), .A2(G79), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G92), .A2(n793), .ZN(n599) );
  NAND2_X1 U673 ( .A1(G66), .A2(n597), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G54), .A2(n600), .ZN(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT75), .B(n601), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X2 U678 ( .A(KEYINPUT15), .B(n606), .ZN(n955) );
  NAND2_X1 U679 ( .A1(G1348), .A2(n780), .ZN(n607) );
  XNOR2_X1 U680 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n620) );
  NAND2_X1 U681 ( .A1(n607), .A2(n620), .ZN(n608) );
  NOR2_X1 U682 ( .A1(G1341), .A2(n608), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n647), .A2(n609), .ZN(n627) );
  NOR2_X1 U684 ( .A1(G1996), .A2(n620), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G56), .A2(n794), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT14), .B(n610), .Z(n616) );
  NAND2_X1 U687 ( .A1(n793), .A2(G81), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT12), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G68), .A2(n797), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT13), .B(n614), .Z(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n798), .A2(G43), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n957) );
  NOR2_X1 U695 ( .A1(n619), .A2(n957), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n780), .A2(G2067), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G1996), .A2(n620), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n623), .A2(n647), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U701 ( .A(n652), .ZN(n667) );
  NAND2_X1 U702 ( .A1(G1348), .A2(n667), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G2067), .A2(n647), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n780), .A2(n630), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n639) );
  NAND2_X1 U707 ( .A1(n633), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(n634), .ZN(n637) );
  NAND2_X1 U709 ( .A1(G1956), .A2(n667), .ZN(n635) );
  XNOR2_X1 U710 ( .A(KEYINPUT95), .B(n635), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n641) );
  INV_X1 U712 ( .A(G299), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n644) );
  OR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n642), .B(KEYINPUT28), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n651) );
  INV_X1 U719 ( .A(G1961), .ZN(n967) );
  NAND2_X1 U720 ( .A1(n667), .A2(n967), .ZN(n649) );
  XNOR2_X1 U721 ( .A(G2078), .B(KEYINPUT25), .ZN(n1014) );
  NAND2_X1 U722 ( .A1(n647), .A2(n1014), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n660) );
  NAND2_X1 U724 ( .A1(n660), .A2(G171), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n666) );
  NAND2_X1 U726 ( .A1(G8), .A2(n667), .ZN(n687) );
  NOR2_X1 U727 ( .A1(G1966), .A2(n687), .ZN(n681) );
  INV_X1 U728 ( .A(G2084), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT94), .ZN(n678) );
  INV_X1 U730 ( .A(n678), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n655), .A2(G8), .ZN(n656) );
  NOR2_X1 U732 ( .A1(n681), .A2(n656), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U734 ( .A1(G168), .A2(n659), .ZN(n662) );
  NOR2_X1 U735 ( .A1(G171), .A2(n660), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n679) );
  NAND2_X1 U739 ( .A1(n679), .A2(G286), .ZN(n673) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n687), .ZN(n669) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G303), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT96), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n676), .A2(G8), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT32), .ZN(n685) );
  NAND2_X1 U749 ( .A1(n678), .A2(G8), .ZN(n683) );
  INV_X1 U750 ( .A(n679), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n698) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n693) );
  NOR2_X1 U755 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n693), .A2(n686), .ZN(n960) );
  NAND2_X1 U757 ( .A1(n698), .A2(n960), .ZN(n691) );
  NAND2_X1 U758 ( .A1(G288), .A2(G1976), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT98), .ZN(n961) );
  NOR2_X1 U760 ( .A1(KEYINPUT33), .A2(n692), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n693), .A2(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n687), .A2(n694), .ZN(n696) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n949) );
  NOR2_X1 U764 ( .A1(n697), .A2(n516), .ZN(n707) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U766 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n698), .A2(n700), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n701), .A2(n687), .ZN(n705) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XOR2_X1 U770 ( .A(n702), .B(KEYINPUT24), .Z(n703) );
  OR2_X1 U771 ( .A1(n687), .A2(n703), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U774 ( .A(KEYINPUT99), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n709), .B(n708), .ZN(n744) );
  NOR2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n760) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n758) );
  XNOR2_X1 U778 ( .A(KEYINPUT34), .B(KEYINPUT88), .ZN(n715) );
  NAND2_X1 U779 ( .A1(G104), .A2(n585), .ZN(n713) );
  NAND2_X1 U780 ( .A1(G140), .A2(n887), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U782 ( .A(n715), .B(n714), .ZN(n721) );
  XNOR2_X1 U783 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n719) );
  NAND2_X1 U784 ( .A1(G128), .A2(n890), .ZN(n717) );
  NAND2_X1 U785 ( .A1(G116), .A2(n891), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U787 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U789 ( .A(n722), .B(KEYINPUT36), .ZN(n866) );
  NOR2_X1 U790 ( .A1(n758), .A2(n866), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n723), .B(KEYINPUT90), .ZN(n936) );
  NAND2_X1 U792 ( .A1(n760), .A2(n936), .ZN(n756) );
  BUF_X1 U793 ( .A(n585), .Z(n886) );
  NAND2_X1 U794 ( .A1(G95), .A2(n886), .ZN(n725) );
  NAND2_X1 U795 ( .A1(G131), .A2(n887), .ZN(n724) );
  NAND2_X1 U796 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U797 ( .A(KEYINPUT92), .B(n726), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G119), .A2(n890), .ZN(n727) );
  XNOR2_X1 U799 ( .A(KEYINPUT91), .B(n727), .ZN(n728) );
  NOR2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n891), .A2(G107), .ZN(n730) );
  NAND2_X1 U802 ( .A1(n731), .A2(n730), .ZN(n881) );
  AND2_X1 U803 ( .A1(n881), .A2(G1991), .ZN(n741) );
  NAND2_X1 U804 ( .A1(G105), .A2(n886), .ZN(n732) );
  XNOR2_X1 U805 ( .A(n732), .B(KEYINPUT38), .ZN(n739) );
  NAND2_X1 U806 ( .A1(G117), .A2(n891), .ZN(n734) );
  NAND2_X1 U807 ( .A1(G141), .A2(n887), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n737) );
  NAND2_X1 U809 ( .A1(G129), .A2(n890), .ZN(n735) );
  XNOR2_X1 U810 ( .A(KEYINPUT93), .B(n735), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n867) );
  AND2_X1 U813 ( .A1(n867), .A2(G1996), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n934) );
  INV_X1 U815 ( .A(n934), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n742), .A2(n760), .ZN(n750) );
  NAND2_X1 U817 ( .A1(n756), .A2(n750), .ZN(n743) );
  NOR2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U819 ( .A(n745), .B(KEYINPUT100), .ZN(n747) );
  XNOR2_X1 U820 ( .A(G1986), .B(G290), .ZN(n953) );
  NAND2_X1 U821 ( .A1(n760), .A2(n953), .ZN(n746) );
  NAND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n749) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n867), .ZN(n929) );
  INV_X1 U824 ( .A(n750), .ZN(n753) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U826 ( .A1(G1991), .A2(n881), .ZN(n940) );
  NOR2_X1 U827 ( .A1(n751), .A2(n940), .ZN(n752) );
  NOR2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U829 ( .A1(n929), .A2(n754), .ZN(n755) );
  XNOR2_X1 U830 ( .A(n755), .B(KEYINPUT39), .ZN(n757) );
  NAND2_X1 U831 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U832 ( .A1(n866), .A2(n758), .ZN(n933) );
  NAND2_X1 U833 ( .A1(n759), .A2(n933), .ZN(n761) );
  NAND2_X1 U834 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U835 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n765), .B(n764), .ZN(G329) );
  AND2_X1 U837 ( .A1(n767), .A2(n766), .ZN(G160) );
  NAND2_X1 U838 ( .A1(G99), .A2(n585), .ZN(n769) );
  NAND2_X1 U839 ( .A1(G111), .A2(n891), .ZN(n768) );
  NAND2_X1 U840 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U841 ( .A(KEYINPUT78), .B(n770), .ZN(n773) );
  NAND2_X1 U842 ( .A1(n890), .A2(G123), .ZN(n771) );
  XOR2_X1 U843 ( .A(KEYINPUT18), .B(n771), .Z(n772) );
  NOR2_X1 U844 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U845 ( .A1(n887), .A2(G135), .ZN(n774) );
  NAND2_X1 U846 ( .A1(n775), .A2(n774), .ZN(n937) );
  XNOR2_X1 U847 ( .A(G2096), .B(n937), .ZN(n776) );
  OR2_X1 U848 ( .A1(G2100), .A2(n776), .ZN(G156) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  INV_X1 U851 ( .A(G120), .ZN(G236) );
  NAND2_X1 U852 ( .A1(G94), .A2(G452), .ZN(n777) );
  XOR2_X1 U853 ( .A(KEYINPUT72), .B(n777), .Z(G173) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U855 ( .A(n778), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U856 ( .A(G223), .B(KEYINPUT74), .Z(n829) );
  NAND2_X1 U857 ( .A1(n829), .A2(G567), .ZN(n779) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n785) );
  OR2_X1 U860 ( .A1(n957), .A2(n785), .ZN(G153) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n782) );
  INV_X1 U862 ( .A(G868), .ZN(n811) );
  NAND2_X1 U863 ( .A1(n780), .A2(n811), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n782), .A2(n781), .ZN(G284) );
  NOR2_X1 U865 ( .A1(G286), .A2(n811), .ZN(n784) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U867 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n785), .A2(G559), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n786), .A2(n955), .ZN(n787) );
  XNOR2_X1 U870 ( .A(n787), .B(KEYINPUT76), .ZN(n788) );
  XNOR2_X1 U871 ( .A(KEYINPUT16), .B(n788), .ZN(G148) );
  NOR2_X1 U872 ( .A1(G868), .A2(n957), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G868), .A2(n955), .ZN(n789) );
  NOR2_X1 U874 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U876 ( .A(KEYINPUT77), .B(n792), .Z(G282) );
  INV_X1 U877 ( .A(G303), .ZN(G166) );
  NAND2_X1 U878 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G67), .A2(n794), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n802) );
  NAND2_X1 U881 ( .A1(G80), .A2(n797), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U884 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U885 ( .A(KEYINPUT79), .B(n803), .Z(n836) );
  XNOR2_X1 U886 ( .A(G305), .B(n836), .ZN(n805) );
  XOR2_X1 U887 ( .A(G299), .B(G166), .Z(n804) );
  XNOR2_X1 U888 ( .A(n805), .B(n804), .ZN(n808) );
  XOR2_X1 U889 ( .A(KEYINPUT19), .B(G290), .Z(n806) );
  XNOR2_X1 U890 ( .A(G288), .B(n806), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n808), .B(n807), .ZN(n901) );
  NAND2_X1 U892 ( .A1(G559), .A2(n955), .ZN(n809) );
  XNOR2_X1 U893 ( .A(n957), .B(n809), .ZN(n835) );
  XNOR2_X1 U894 ( .A(n901), .B(n835), .ZN(n810) );
  NOR2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n813) );
  NOR2_X1 U896 ( .A1(n836), .A2(G868), .ZN(n812) );
  NOR2_X1 U897 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U898 ( .A(KEYINPUT84), .B(n814), .Z(G295) );
  NAND2_X1 U899 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XNOR2_X1 U900 ( .A(n815), .B(KEYINPUT20), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n816), .B(KEYINPUT85), .ZN(n817) );
  NAND2_X1 U902 ( .A1(n817), .A2(G2090), .ZN(n818) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U906 ( .A1(G69), .A2(G57), .ZN(n820) );
  NOR2_X1 U907 ( .A1(G236), .A2(n820), .ZN(n821) );
  XNOR2_X1 U908 ( .A(KEYINPUT86), .B(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n822), .A2(G108), .ZN(n833) );
  NAND2_X1 U910 ( .A1(n833), .A2(G567), .ZN(n827) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U913 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U914 ( .A1(G96), .A2(n825), .ZN(n834) );
  NAND2_X1 U915 ( .A1(n834), .A2(G2106), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n827), .A2(n826), .ZN(n838) );
  NAND2_X1 U917 ( .A1(G483), .A2(G661), .ZN(n828) );
  NOR2_X1 U918 ( .A1(n838), .A2(n828), .ZN(n832) );
  NAND2_X1 U919 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U922 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U925 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  NOR2_X1 U926 ( .A1(n834), .A2(n833), .ZN(G325) );
  XNOR2_X1 U927 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G57), .ZN(G237) );
  NOR2_X1 U932 ( .A1(n835), .A2(G860), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(G145) );
  INV_X1 U934 ( .A(n838), .ZN(G319) );
  XOR2_X1 U935 ( .A(G2096), .B(KEYINPUT106), .Z(n840) );
  XNOR2_X1 U936 ( .A(G2090), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U938 ( .A(n841), .B(KEYINPUT42), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U941 ( .A(G2678), .B(G2100), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n849) );
  XOR2_X1 U946 ( .A(G1991), .B(n967), .Z(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(G1981), .B(G1956), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT107), .B(G2474), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(KEYINPUT41), .B(n856), .ZN(n857) );
  XOR2_X1 U955 ( .A(n857), .B(G1996), .Z(G229) );
  NAND2_X1 U956 ( .A1(G112), .A2(n891), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G136), .A2(n887), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G100), .A2(n585), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT108), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(G162) );
  XNOR2_X1 U965 ( .A(G160), .B(n866), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n885) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT110), .B(KEYINPUT48), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n879) );
  NAND2_X1 U970 ( .A1(G130), .A2(n890), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G118), .A2(n891), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G106), .A2(n886), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G142), .A2(n887), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(n879), .B(n878), .Z(n880) );
  XOR2_X1 U979 ( .A(n880), .B(G162), .Z(n883) );
  XOR2_X1 U980 ( .A(G164), .B(n881), .Z(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n898) );
  NAND2_X1 U983 ( .A1(G103), .A2(n886), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U986 ( .A1(G127), .A2(n890), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n924) );
  XNOR2_X1 U991 ( .A(n937), .B(n924), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G37), .A2(n899), .ZN(n900) );
  XOR2_X1 U994 ( .A(KEYINPUT111), .B(n900), .Z(G395) );
  XNOR2_X1 U995 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n957), .B(n901), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(n904), .B(G171), .Z(n905) );
  XOR2_X1 U999 ( .A(n905), .B(n955), .Z(n906) );
  XOR2_X1 U1000 ( .A(G286), .B(n906), .Z(n907) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1002 ( .A(G2454), .B(G2435), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G2438), .B(G2427), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n916) );
  XOR2_X1 U1005 ( .A(KEYINPUT103), .B(G2446), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G2443), .B(G2430), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n912), .B(G2451), .Z(n914) );
  XNOR2_X1 U1009 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1021 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT50), .B(n927), .ZN(n932) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n945) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n943) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT114), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(KEYINPUT115), .ZN(n1024) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n1024), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n948), .A2(G29), .ZN(n1031) );
  INV_X1 U1041 ( .A(G16), .ZN(n1001) );
  XOR2_X1 U1042 ( .A(n1001), .B(KEYINPUT56), .Z(n976) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT57), .B(n951), .ZN(n974) );
  XOR2_X1 U1046 ( .A(G299), .B(G1956), .Z(n952) );
  XNOR2_X1 U1047 ( .A(n952), .B(KEYINPUT121), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n971) );
  XNOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT120), .ZN(n956) );
  XOR2_X1 U1050 ( .A(n956), .B(n955), .Z(n959) );
  XNOR2_X1 U1051 ( .A(G1341), .B(n957), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n966) );
  AND2_X1 U1053 ( .A1(G303), .A2(G1971), .ZN(n963) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n964), .B(KEYINPUT122), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1058 ( .A(n967), .B(G301), .Z(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(KEYINPUT123), .B(n972), .ZN(n973) );
  NAND2_X1 U1062 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1063 ( .A1(n976), .A2(n975), .ZN(n1003) );
  XOR2_X1 U1064 ( .A(G1966), .B(G21), .Z(n984) );
  XNOR2_X1 U1065 ( .A(G1986), .B(G24), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G22), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G1976), .B(G23), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(KEYINPUT125), .B(n979), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT58), .B(n982), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n997) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n985), .B(G4), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G20), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G1981), .B(G6), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(G1341), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(G19), .B(n990), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(KEYINPUT60), .ZN(n995) );
  XOR2_X1 U1083 ( .A(G1961), .B(G5), .Z(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n999), .B(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1029) );
  XNOR2_X1 U1090 ( .A(KEYINPUT54), .B(G34), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1004), .B(KEYINPUT117), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G2084), .B(n1005), .ZN(n1021) );
  XNOR2_X1 U1093 ( .A(G2090), .B(G35), .ZN(n1019) );
  XNOR2_X1 U1094 ( .A(G2067), .B(G26), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G33), .B(G2072), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(G32), .B(G1996), .Z(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(G28), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G25), .B(G1991), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT116), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G27), .B(n1014), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT53), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT118), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(n1024), .B(n1023), .Z(n1025) );
  OR2_X1 U1110 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(G11), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT119), .B(n1027), .Z(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

