

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  INV_X1 U323 ( .A(n523), .ZN(n509) );
  INV_X1 U324 ( .A(n547), .ZN(n584) );
  XNOR2_X1 U325 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U326 ( .A(n420), .B(n419), .ZN(n423) );
  XNOR2_X1 U327 ( .A(n418), .B(n291), .ZN(n419) );
  XOR2_X1 U328 ( .A(n417), .B(n416), .Z(n291) );
  INV_X1 U329 ( .A(KEYINPUT45), .ZN(n428) );
  XOR2_X1 U330 ( .A(G169GAT), .B(G8GAT), .Z(n444) );
  XNOR2_X1 U331 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U332 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U333 ( .A(n404), .B(n403), .ZN(n427) );
  XNOR2_X1 U334 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U335 ( .A(KEYINPUT83), .B(KEYINPUT65), .Z(n293) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U338 ( .A(G120GAT), .B(G71GAT), .Z(n398) );
  XOR2_X1 U339 ( .A(n294), .B(n398), .Z(n296) );
  XNOR2_X1 U340 ( .A(G169GAT), .B(G15GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n302) );
  XOR2_X1 U342 ( .A(G127GAT), .B(KEYINPUT0), .Z(n298) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G134GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n329) );
  XOR2_X1 U345 ( .A(G176GAT), .B(n329), .Z(n300) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U348 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U349 ( .A(KEYINPUT18), .B(G190GAT), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT17), .B(n305), .ZN(n447) );
  XOR2_X1 U353 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n307) );
  XNOR2_X1 U354 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n447), .B(n308), .Z(n309) );
  XOR2_X1 U357 ( .A(n310), .B(n309), .Z(n525) );
  INV_X1 U358 ( .A(n525), .ZN(n533) );
  XOR2_X1 U359 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n312) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U362 ( .A(n313), .B(KEYINPUT85), .Z(n317) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(G78GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n314), .B(G148GAT), .ZN(n389) );
  XNOR2_X1 U365 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n315), .B(KEYINPUT3), .ZN(n336) );
  XNOR2_X1 U367 ( .A(n389), .B(n336), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U369 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n319) );
  XOR2_X1 U370 ( .A(G141GAT), .B(G22GAT), .Z(n372) );
  XOR2_X1 U371 ( .A(KEYINPUT76), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U372 ( .A(n372), .B(n409), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n323) );
  XNOR2_X1 U375 ( .A(G50GAT), .B(KEYINPUT84), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n328) );
  XOR2_X1 U377 ( .A(KEYINPUT21), .B(G204GAT), .Z(n325) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G211GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U380 ( .A(G218GAT), .B(KEYINPUT86), .Z(n326) );
  XOR2_X1 U381 ( .A(n327), .B(n326), .Z(n442) );
  XOR2_X1 U382 ( .A(n328), .B(n442), .Z(n471) );
  XOR2_X1 U383 ( .A(G162GAT), .B(n329), .Z(n331) );
  NAND2_X1 U384 ( .A1(G225GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U386 ( .A(G29GAT), .B(n332), .ZN(n348) );
  XOR2_X1 U387 ( .A(KEYINPUT6), .B(KEYINPUT88), .Z(n338) );
  XOR2_X1 U388 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n334) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U393 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n340) );
  XNOR2_X1 U394 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U396 ( .A(G85GAT), .B(G148GAT), .Z(n342) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(G120GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U399 ( .A(n344), .B(n343), .Z(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U401 ( .A(n348), .B(n347), .Z(n521) );
  INV_X1 U402 ( .A(n521), .ZN(n505) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G1GAT), .Z(n379) );
  XOR2_X1 U404 ( .A(G155GAT), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U405 ( .A(G22GAT), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n379), .B(n351), .Z(n353) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n354), .B(KEYINPUT79), .Z(n357) );
  XNOR2_X1 U411 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n355), .B(KEYINPUT13), .ZN(n396) );
  XNOR2_X1 U413 ( .A(n396), .B(KEYINPUT14), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U415 ( .A(G71GAT), .B(G127GAT), .Z(n359) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(G183GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n361) );
  XNOR2_X1 U419 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U421 ( .A(n363), .B(n362), .Z(n364) );
  XOR2_X1 U422 ( .A(n365), .B(n364), .Z(n547) );
  XNOR2_X1 U423 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n366), .B(G29GAT), .ZN(n367) );
  XOR2_X1 U425 ( .A(n367), .B(KEYINPUT7), .Z(n369) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(G50GAT), .ZN(n368) );
  XOR2_X1 U427 ( .A(n369), .B(n368), .Z(n421) );
  XOR2_X1 U428 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n371) );
  XNOR2_X1 U429 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U431 ( .A(n373), .B(n372), .Z(n377) );
  XOR2_X1 U432 ( .A(n444), .B(KEYINPUT30), .Z(n375) );
  NAND2_X1 U433 ( .A1(G229GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n381) );
  XNOR2_X1 U436 ( .A(G197GAT), .B(G113GAT), .ZN(n378) );
  XOR2_X1 U437 ( .A(n421), .B(n382), .Z(n578) );
  INV_X1 U438 ( .A(G92GAT), .ZN(n383) );
  NAND2_X1 U439 ( .A1(n383), .A2(KEYINPUT74), .ZN(n386) );
  INV_X1 U440 ( .A(KEYINPUT74), .ZN(n384) );
  NAND2_X1 U441 ( .A1(n384), .A2(G92GAT), .ZN(n385) );
  NAND2_X1 U442 ( .A1(n386), .A2(n385), .ZN(n388) );
  XNOR2_X1 U443 ( .A(G99GAT), .B(G85GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n410) );
  XNOR2_X1 U445 ( .A(n389), .B(n410), .ZN(n395) );
  XNOR2_X1 U446 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n391) );
  NAND2_X1 U447 ( .A1(G230GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n393) );
  INV_X1 U449 ( .A(KEYINPUT32), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n404) );
  XOR2_X1 U453 ( .A(G176GAT), .B(G64GAT), .Z(n435) );
  XNOR2_X1 U454 ( .A(n398), .B(n435), .ZN(n402) );
  XOR2_X1 U455 ( .A(KEYINPUT75), .B(KEYINPUT73), .Z(n400) );
  XNOR2_X1 U456 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U458 ( .A(KEYINPUT41), .B(n427), .Z(n559) );
  AND2_X1 U459 ( .A1(n578), .A2(n559), .ZN(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n407) );
  NOR2_X1 U462 ( .A1(n584), .A2(n407), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n408), .B(KEYINPUT110), .ZN(n424) );
  XOR2_X1 U464 ( .A(n410), .B(n409), .Z(n412) );
  XNOR2_X1 U465 ( .A(G190GAT), .B(G218GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n420) );
  XOR2_X1 U467 ( .A(KEYINPUT77), .B(KEYINPUT66), .Z(n414) );
  XNOR2_X1 U468 ( .A(G134GAT), .B(G106GAT), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n415), .B(KEYINPUT10), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n417) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n416) );
  INV_X1 U473 ( .A(n421), .ZN(n422) );
  XOR2_X1 U474 ( .A(n423), .B(n422), .Z(n551) );
  NAND2_X1 U475 ( .A1(n424), .A2(n551), .ZN(n425) );
  XNOR2_X1 U476 ( .A(n425), .B(KEYINPUT47), .ZN(n426) );
  XNOR2_X1 U477 ( .A(n426), .B(KEYINPUT111), .ZN(n433) );
  BUF_X1 U478 ( .A(n427), .Z(n581) );
  INV_X1 U479 ( .A(n551), .ZN(n570) );
  XOR2_X1 U480 ( .A(n570), .B(KEYINPUT36), .Z(n589) );
  NOR2_X1 U481 ( .A1(n589), .A2(n547), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  NOR2_X1 U483 ( .A1(n581), .A2(n430), .ZN(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT70), .B(n578), .Z(n539) );
  NAND2_X1 U485 ( .A1(n431), .A2(n539), .ZN(n432) );
  NAND2_X1 U486 ( .A1(n433), .A2(n432), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n434), .B(KEYINPUT48), .ZN(n534) );
  XOR2_X1 U488 ( .A(n435), .B(KEYINPUT94), .Z(n437) );
  NAND2_X1 U489 ( .A1(G226GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U491 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n439) );
  XNOR2_X1 U492 ( .A(G36GAT), .B(G92GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U494 ( .A(n441), .B(n440), .Z(n446) );
  INV_X1 U495 ( .A(n442), .ZN(n443) );
  XOR2_X1 U496 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n449) );
  INV_X1 U498 ( .A(n447), .ZN(n448) );
  XOR2_X1 U499 ( .A(n449), .B(n448), .Z(n523) );
  NAND2_X1 U500 ( .A1(n534), .A2(n523), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U503 ( .A1(n505), .A2(n452), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT64), .ZN(n577) );
  NOR2_X1 U505 ( .A1(n471), .A2(n577), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NOR2_X2 U507 ( .A1(n533), .A2(n455), .ZN(n456) );
  XOR2_X2 U508 ( .A(KEYINPUT121), .B(n456), .Z(n571) );
  INV_X1 U509 ( .A(n539), .ZN(n457) );
  NAND2_X1 U510 ( .A1(n571), .A2(n457), .ZN(n459) );
  XNOR2_X1 U511 ( .A(KEYINPUT122), .B(G169GAT), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(G1348GAT) );
  NAND2_X1 U513 ( .A1(n571), .A2(n559), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n461) );
  XOR2_X1 U515 ( .A(G176GAT), .B(KEYINPUT56), .Z(n460) );
  XNOR2_X1 U516 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NOR2_X1 U517 ( .A1(n539), .A2(n581), .ZN(n495) );
  XOR2_X1 U518 ( .A(n471), .B(KEYINPUT28), .Z(n515) );
  INV_X1 U519 ( .A(n515), .ZN(n532) );
  XOR2_X1 U520 ( .A(n509), .B(KEYINPUT95), .Z(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT27), .ZN(n473) );
  NOR2_X1 U522 ( .A1(n505), .A2(n473), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT96), .ZN(n535) );
  NAND2_X1 U524 ( .A1(n533), .A2(n535), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n532), .A2(n466), .ZN(n478) );
  NAND2_X1 U526 ( .A1(n523), .A2(n525), .ZN(n467) );
  XNOR2_X1 U527 ( .A(KEYINPUT97), .B(n467), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n471), .A2(n468), .ZN(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n469), .Z(n470) );
  XNOR2_X1 U530 ( .A(KEYINPUT98), .B(n470), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n471), .A2(n533), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT26), .ZN(n576) );
  NOR2_X1 U533 ( .A1(n576), .A2(n473), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n521), .A2(n476), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n492) );
  NOR2_X1 U537 ( .A1(n547), .A2(n570), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U539 ( .A1(n492), .A2(n480), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n495), .A2(n504), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n505), .A2(n489), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT99), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U545 ( .A1(n509), .A2(n489), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(n484), .Z(n485) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n485), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n533), .A2(n489), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT35), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NOR2_X1 U552 ( .A1(n515), .A2(n489), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(n490), .Z(n491) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  NOR2_X1 U555 ( .A1(n492), .A2(n589), .ZN(n493) );
  NAND2_X1 U556 ( .A1(n493), .A2(n547), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(KEYINPUT37), .ZN(n518) );
  NAND2_X1 U558 ( .A1(n495), .A2(n518), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT38), .ZN(n502) );
  NOR2_X1 U560 ( .A1(n502), .A2(n505), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n502), .A2(n509), .ZN(n499) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U565 ( .A1(n533), .A2(n502), .ZN(n500) );
  XOR2_X1 U566 ( .A(KEYINPUT40), .B(n500), .Z(n501) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U568 ( .A1(n515), .A2(n502), .ZN(n503) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  INV_X1 U570 ( .A(n559), .ZN(n542) );
  NOR2_X1 U571 ( .A1(n542), .A2(n578), .ZN(n519) );
  NAND2_X1 U572 ( .A1(n519), .A2(n504), .ZN(n514) );
  NOR2_X1 U573 ( .A1(n505), .A2(n514), .ZN(n507) );
  XNOR2_X1 U574 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n509), .A2(n514), .ZN(n510) );
  XOR2_X1 U578 ( .A(KEYINPUT104), .B(n510), .Z(n511) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n533), .A2(n514), .ZN(n513) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n515), .A2(n514), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U587 ( .A(KEYINPUT106), .B(n520), .Z(n528) );
  NAND2_X1 U588 ( .A1(n521), .A2(n528), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT107), .Z(n527) );
  NAND2_X1 U593 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n530) );
  NAND2_X1 U596 ( .A1(n528), .A2(n532), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n531), .Z(G1339GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT112), .B(n536), .ZN(n554) );
  INV_X1 U602 ( .A(n554), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n539), .A2(n550), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  NOR2_X1 U607 ( .A1(n542), .A2(n550), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n546) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n549) );
  NOR2_X1 U613 ( .A1(n547), .A2(n550), .ZN(n548) );
  XOR2_X1 U614 ( .A(n549), .B(n548), .Z(G1342GAT) );
  NOR2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n576), .A2(n554), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n565), .A2(n578), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n557) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT116), .B(n558), .Z(n561) );
  NAND2_X1 U625 ( .A1(n565), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U628 ( .A1(n565), .A2(n584), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n570), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n584), .A2(n571), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT124), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(n569), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1351GAT) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT60), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n575), .Z(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

