//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT66), .B(G77), .Z(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT67), .B(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G87), .B(G97), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND2_X1  g0041(.A1(new_n210), .A2(G33), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT8), .B(G58), .Z(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n211), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n250), .ZN(new_n252));
  OR2_X1    g0052(.A1(KEYINPUT68), .A2(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT68), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G20), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n253), .A2(G13), .A3(G20), .A4(new_n254), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n251), .B(new_n259), .C1(G50), .C2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT9), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G222), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G223), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n269), .B(new_n270), .C1(new_n216), .C2(new_n265), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G41), .A2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  INV_X1    g0076(.A(new_n211), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n255), .B2(new_n272), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n271), .B(new_n275), .C1(new_n276), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  INV_X1    g0083(.A(G190), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n262), .B(new_n283), .C1(new_n284), .C2(new_n282), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT10), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n261), .B(new_n288), .C1(G179), .C2(new_n282), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1698), .B1(new_n263), .B2(new_n264), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n270), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  INV_X1    g0096(.A(new_n275), .ZN(new_n297));
  INV_X1    g0097(.A(new_n281), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(G238), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n280), .B1(new_n292), .B2(new_n293), .ZN(new_n301));
  INV_X1    g0101(.A(G238), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n275), .B1(new_n281), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT13), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT70), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n295), .A2(new_n299), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(G169), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT14), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n306), .A2(new_n308), .A3(new_n311), .A4(G169), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n300), .A2(new_n304), .A3(G179), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n258), .A2(G68), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT71), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT72), .B1(new_n260), .B2(G68), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n317), .B(KEYINPUT12), .Z(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n246), .A2(G50), .B1(G20), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G77), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n242), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n250), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n316), .B(new_n318), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n284), .B1(new_n307), .B2(KEYINPUT13), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n300), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n306), .A2(G200), .A3(new_n308), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n260), .A2(new_n244), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n258), .B2(new_n244), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n256), .A2(new_n278), .ZN(new_n336));
  INV_X1    g0136(.A(G159), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT73), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT73), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n246), .A2(new_n339), .A3(G159), .ZN(new_n340));
  XNOR2_X1  g0140(.A(G58), .B(G68), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n338), .A2(new_n340), .B1(G20), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(G20), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  OAI21_X1  g0146(.A(G68), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n343), .A2(new_n344), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n348), .A2(new_n210), .A3(new_n346), .ZN(new_n349));
  OAI211_X1 g0149(.A(KEYINPUT16), .B(new_n342), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n250), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n256), .A2(KEYINPUT64), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT64), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT7), .B1(new_n265), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n345), .A2(new_n346), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT16), .B1(new_n358), .B2(new_n342), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n335), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n280), .B(G232), .C1(new_n255), .C2(new_n272), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n275), .ZN(new_n363));
  OR2_X1    g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n276), .A2(G1698), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n265), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n280), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n361), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n364), .A2(new_n365), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n370), .B2(new_n348), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n270), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(new_n284), .A3(new_n275), .A4(new_n362), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n333), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(G58), .A2(G68), .ZN(new_n376));
  OAI21_X1  g0176(.A(G20), .B1(new_n376), .B2(new_n201), .ZN(new_n377));
  NOR4_X1   g0177(.A1(new_n337), .A2(KEYINPUT73), .A3(G20), .A4(G33), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n339), .B1(new_n246), .B2(G159), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n348), .A2(new_n210), .A3(new_n346), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n263), .A2(new_n256), .A3(new_n264), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n319), .B1(new_n382), .B2(KEYINPUT7), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n252), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n346), .B1(new_n348), .B2(new_n210), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT7), .A4(G20), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n387), .A2(new_n388), .A3(new_n319), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n389), .B2(new_n380), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n369), .A2(new_n373), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n335), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT74), .B1(new_n375), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n335), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n385), .B2(new_n390), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n363), .B2(new_n368), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n372), .A2(G179), .A3(new_n275), .A4(new_n362), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT18), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n360), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n375), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n395), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT15), .B(G87), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n243), .A2(new_n409), .B1(new_n216), .B2(new_n355), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n244), .B(KEYINPUT69), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(new_n336), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n250), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n413), .B1(new_n321), .B2(new_n257), .C1(new_n216), .C2(new_n260), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n298), .A2(new_n217), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n265), .A2(G232), .A3(new_n267), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n265), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n297), .B(new_n415), .C1(new_n270), .C2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n414), .B1(G190), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n361), .B2(new_n420), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n420), .A2(G169), .ZN(new_n423));
  INV_X1    g0223(.A(G179), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n414), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n290), .A2(new_n332), .A3(new_n407), .A4(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(G257), .B(G1698), .C1(new_n343), .C2(new_n344), .ZN(new_n429));
  OAI211_X1 g0229(.A(G250), .B(new_n267), .C1(new_n343), .C2(new_n344), .ZN(new_n430));
  INV_X1    g0230(.A(G294), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(new_n430), .C1(new_n278), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n270), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n253), .A2(G45), .A3(new_n254), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT5), .B(G41), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(G274), .A3(new_n280), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n436), .ZN(new_n438));
  OAI211_X1 g0238(.A(G264), .B(new_n280), .C1(new_n438), .C2(new_n434), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n433), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G169), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(KEYINPUT77), .A3(G169), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n433), .A2(G179), .A3(new_n437), .A4(new_n439), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n265), .A2(new_n210), .A3(G87), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT22), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT22), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n265), .A2(new_n210), .A3(new_n449), .A4(G87), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n256), .A2(G33), .A3(G116), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT23), .B1(new_n256), .B2(G107), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(KEYINPUT76), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n452), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n451), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n451), .B2(new_n457), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n250), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n260), .A2(G107), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n462), .A2(KEYINPUT25), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(KEYINPUT25), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n253), .A2(G33), .A3(new_n254), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n260), .A2(new_n252), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n463), .A2(new_n464), .B1(G107), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT78), .B1(new_n446), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n440), .A2(new_n361), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(G190), .B2(new_n440), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n461), .A2(new_n468), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n470), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G264), .B(G1698), .C1(new_n343), .C2(new_n344), .ZN(new_n481));
  OAI211_X1 g0281(.A(G257), .B(new_n267), .C1(new_n343), .C2(new_n344), .ZN(new_n482));
  INV_X1    g0282(.A(G303), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(new_n265), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n270), .ZN(new_n485));
  OAI211_X1 g0285(.A(G270), .B(new_n280), .C1(new_n438), .C2(new_n434), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n437), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G200), .ZN(new_n488));
  INV_X1    g0288(.A(new_n260), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n260), .A2(new_n252), .A3(new_n465), .A4(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n210), .B(new_n494), .C1(G33), .C2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n249), .A2(new_n211), .B1(G20), .B2(new_n490), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT20), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT20), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n493), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n488), .B(new_n501), .C1(new_n284), .C2(new_n487), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT21), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n487), .A2(G169), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n501), .ZN(new_n505));
  INV_X1    g0305(.A(new_n500), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n491), .B(new_n492), .C1(new_n506), .C2(new_n498), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(new_n487), .A3(KEYINPUT21), .A4(G169), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n487), .A2(new_n424), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n507), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n502), .A2(new_n505), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  XOR2_X1   g0312(.A(G97), .B(G107), .Z(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n495), .A2(G107), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n355), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n356), .A2(new_n357), .A3(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n246), .A2(G77), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n250), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n489), .A2(new_n495), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n467), .A2(G97), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(new_n267), .C1(new_n343), .C2(new_n344), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n494), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n270), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(new_n280), .C1(new_n438), .C2(new_n434), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n437), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n534), .A3(new_n424), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n287), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n525), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n524), .A2(new_n523), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n521), .B2(new_n250), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n541), .C1(new_n284), .C2(new_n536), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n242), .B2(new_n495), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  INV_X1    g0345(.A(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n543), .A2(new_n278), .A3(new_n495), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n355), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n265), .A2(new_n210), .A3(G68), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n250), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n489), .A2(new_n408), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n467), .A2(new_n409), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n291), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n265), .A2(G244), .A3(G1698), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n280), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n435), .A2(G274), .A3(new_n280), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n280), .A2(new_n434), .A3(G250), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n287), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n270), .ZN(new_n564));
  INV_X1    g0364(.A(new_n561), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n424), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(G190), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n551), .A2(new_n250), .B1(new_n489), .B2(new_n408), .ZN(new_n569));
  OAI21_X1  g0369(.A(G200), .B1(new_n558), .B2(new_n561), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n467), .A2(G87), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n512), .A2(new_n538), .A3(new_n542), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n480), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n428), .A2(new_n576), .ZN(G372));
  NOR2_X1   g0377(.A1(new_n573), .A2(new_n538), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT26), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n538), .A2(new_n542), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n573), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n475), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n446), .A2(new_n469), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n505), .A2(new_n510), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n508), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n579), .B(new_n567), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n428), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n426), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n331), .B1(new_n314), .B2(new_n326), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n375), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(new_n394), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n405), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n286), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n595), .A2(new_n289), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n588), .A2(new_n596), .ZN(G369));
  AND3_X1   g0397(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n478), .B1(new_n476), .B2(new_n477), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n210), .A2(G13), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n601), .A2(KEYINPUT27), .A3(new_n255), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT27), .B1(new_n601), .B2(new_n255), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(G213), .ZN(new_n604));
  INV_X1    g0404(.A(G343), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n584), .B2(new_n508), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(new_n475), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n606), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n583), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(KEYINPUT81), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n609), .A2(new_n501), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n585), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n511), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g0417(.A(KEYINPUT80), .B(G330), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n583), .A2(new_n606), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n469), .A2(new_n609), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n480), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n612), .A2(new_n624), .ZN(G399));
  NOR2_X1   g0425(.A1(new_n547), .A2(G116), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n626), .B(KEYINPUT82), .Z(new_n627));
  INV_X1    g0427(.A(new_n207), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n628), .A2(G41), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n627), .A2(new_n274), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n214), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT28), .Z(new_n633));
  AND2_X1   g0433(.A1(new_n587), .A2(new_n609), .ZN(new_n634));
  INV_X1    g0434(.A(new_n600), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n585), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n579), .B(new_n567), .C1(new_n636), .C2(new_n582), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n609), .ZN(new_n638));
  MUX2_X1   g0438(.A(new_n634), .B(new_n638), .S(KEYINPUT29), .Z(new_n639));
  AND4_X1   g0439(.A1(new_n433), .A2(new_n564), .A3(new_n565), .A4(new_n439), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n509), .A3(new_n532), .A4(new_n534), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT30), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n536), .A2(new_n440), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n487), .B(new_n424), .C1(new_n558), .C2(new_n561), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT83), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n606), .B1(new_n643), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT31), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT31), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n652), .B(new_n606), .C1(new_n643), .C2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT84), .B1(new_n576), .B2(new_n609), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n580), .A2(new_n511), .A3(new_n573), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n600), .A2(new_n656), .A3(new_n475), .A4(new_n609), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT84), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n654), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n618), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n639), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n633), .B1(new_n663), .B2(G1), .ZN(G364));
  INV_X1    g0464(.A(new_n601), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n274), .B1(new_n665), .B2(G45), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n629), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n628), .A2(new_n348), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(G355), .B1(new_n490), .B2(new_n628), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n240), .A2(G45), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n628), .A2(new_n265), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n215), .B2(G45), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n671), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n277), .B1(new_n256), .B2(G169), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT86), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(G13), .A2(G33), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G20), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n669), .B1(new_n676), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n683), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n210), .B2(G190), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n355), .A2(KEYINPUT88), .A3(new_n284), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n424), .A4(G200), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT89), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT89), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(G179), .A2(G200), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n688), .A2(new_n689), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n695), .A2(G283), .B1(G329), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n256), .A2(new_n284), .A3(new_n361), .A4(G179), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n210), .B1(G190), .B2(new_n696), .ZN(new_n703));
  OAI221_X1 g0503(.A(new_n348), .B1(new_n702), .B2(new_n483), .C1(new_n431), .C2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n210), .A2(new_n424), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G190), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n361), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n704), .B1(G326), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G322), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n706), .A2(G200), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n284), .A3(G200), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT33), .B(G317), .Z(new_n713));
  OAI221_X1 g0513(.A(new_n708), .B1(new_n709), .B2(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n705), .A2(new_n284), .A3(new_n361), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT87), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(KEYINPUT87), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n714), .B1(G311), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n700), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n695), .A2(G107), .ZN(new_n723));
  INV_X1    g0523(.A(new_n707), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n724), .A2(new_n202), .B1(new_n319), .B2(new_n712), .ZN(new_n725));
  INV_X1    g0525(.A(G58), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n711), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n703), .A2(new_n495), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n265), .B1(new_n702), .B2(new_n546), .ZN(new_n729));
  NOR4_X1   g0529(.A1(new_n725), .A2(new_n727), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n698), .A2(G159), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT32), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n720), .A2(new_n216), .B1(KEYINPUT32), .B2(new_n731), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n723), .A2(new_n730), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n722), .A2(KEYINPUT91), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n680), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT91), .B1(new_n722), .B2(new_n734), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n685), .B1(new_n616), .B2(new_n686), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n619), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n617), .A2(new_n618), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(new_n669), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(G396));
  INV_X1    g0542(.A(new_n662), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n414), .A2(new_n606), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n589), .B1(new_n422), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n426), .A2(new_n606), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n587), .A3(new_n609), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n747), .B(KEYINPUT93), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(new_n634), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n668), .B1(new_n743), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n743), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n680), .A2(new_n681), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n668), .B1(new_n754), .B2(G77), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n265), .B(new_n728), .C1(G107), .C2(new_n701), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n756), .B1(new_n431), .B2(new_n711), .C1(new_n483), .C2(new_n724), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(G311), .B2(new_n698), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n712), .A2(KEYINPUT92), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n712), .A2(KEYINPUT92), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G116), .A2(new_n720), .B1(new_n762), .B2(G283), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n758), .B(new_n763), .C1(new_n546), .C2(new_n694), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G137), .A2(new_n707), .B1(new_n710), .B2(G143), .ZN(new_n765));
  INV_X1    g0565(.A(G150), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n765), .B1(new_n766), .B2(new_n712), .C1(new_n719), .C2(new_n337), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(KEYINPUT34), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n695), .A2(G68), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n265), .B1(new_n702), .B2(new_n202), .C1(new_n726), .C2(new_n703), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G132), .B2(new_n698), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT34), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n770), .B(new_n772), .C1(new_n773), .C2(new_n767), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n764), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n755), .B1(new_n775), .B2(new_n680), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n682), .B2(new_n747), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n752), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G384));
  OR2_X1    g0579(.A1(new_n515), .A2(new_n517), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n490), .B(new_n213), .C1(new_n780), .C2(KEYINPUT35), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(KEYINPUT35), .B2(new_n780), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT36), .Z(new_n783));
  INV_X1    g0583(.A(new_n255), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n216), .B(new_n631), .C1(new_n726), .C2(new_n319), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n202), .A2(G68), .ZN(new_n786));
  AOI211_X1 g0586(.A(G13), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n746), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n748), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n326), .A2(new_n606), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n327), .A2(new_n331), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT94), .ZN(new_n793));
  INV_X1    g0593(.A(new_n791), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n314), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n314), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(KEYINPUT94), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n792), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT95), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT95), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n792), .A2(new_n797), .A3(new_n800), .A4(new_n795), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n384), .A2(KEYINPUT16), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n335), .B1(new_n351), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n604), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n397), .A2(new_n392), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n360), .A2(new_n400), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n360), .A2(new_n806), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT37), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n805), .A2(new_n400), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n809), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT37), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n407), .A2(new_n808), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n813), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n402), .A2(new_n404), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n591), .A2(new_n394), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(KEYINPUT38), .B(new_n819), .C1(new_n821), .C2(new_n807), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n803), .A2(new_n824), .B1(new_n405), .B2(new_n806), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT98), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n817), .A2(new_n827), .A3(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT96), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n375), .A2(new_n830), .A3(new_n393), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n405), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n375), .B2(new_n393), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n360), .B(new_n806), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n813), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT38), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n828), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(KEYINPUT99), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT99), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n826), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n839), .A2(new_n840), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n848), .A2(KEYINPUT100), .A3(new_n841), .A4(new_n842), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n327), .A2(new_n606), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n825), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT101), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n639), .A2(new_n853), .A3(new_n428), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n639), .B2(new_n428), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n596), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n852), .B(new_n856), .Z(new_n857));
  NAND3_X1  g0657(.A1(new_n802), .A2(new_n660), .A3(new_n747), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n824), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n747), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n576), .A2(KEYINPUT84), .A3(new_n609), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n657), .A2(new_n658), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n864), .B2(new_n654), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n802), .C1(KEYINPUT102), .C2(KEYINPUT40), .ZN(new_n866));
  INV_X1    g0666(.A(new_n839), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n865), .A3(new_n802), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n860), .A2(new_n866), .B1(KEYINPUT40), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n428), .A2(new_n660), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(new_n618), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n857), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n784), .B2(new_n665), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n857), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n788), .B1(new_n874), .B2(new_n875), .ZN(G367));
  OAI211_X1 g0676(.A(new_n538), .B(new_n542), .C1(new_n541), .C2(new_n609), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n538), .B1(new_n600), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n609), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n538), .A2(new_n609), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n877), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n608), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT42), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT103), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n884), .A2(new_n885), .B1(new_n883), .B2(new_n882), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n569), .A2(new_n571), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n606), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n574), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n889), .A2(new_n567), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n886), .A2(new_n887), .B1(KEYINPUT43), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n893), .B(new_n894), .Z(new_n895));
  INV_X1    g0695(.A(new_n881), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n624), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n899), .A2(KEYINPUT105), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(KEYINPUT105), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n895), .A2(new_n898), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n629), .B(KEYINPUT41), .Z(new_n904));
  NAND2_X1  g0704(.A1(new_n612), .A2(new_n881), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n612), .A2(new_n907), .A3(new_n881), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n612), .A2(new_n881), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT45), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(KEYINPUT44), .A3(new_n908), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n624), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT107), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n918), .A3(new_n624), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n608), .B1(new_n622), .B2(new_n607), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n739), .B(new_n920), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n639), .A2(new_n662), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n911), .A2(new_n913), .A3(new_n623), .A4(new_n914), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n917), .A2(new_n919), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n904), .B1(new_n925), .B2(new_n663), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n903), .B1(new_n926), .B2(new_n667), .ZN(new_n927));
  INV_X1    g0727(.A(G283), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n719), .A2(new_n928), .B1(new_n418), .B2(new_n703), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n695), .A2(G97), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n702), .A2(KEYINPUT46), .A3(new_n490), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT46), .B1(new_n702), .B2(new_n490), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n265), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT109), .B(G311), .Z(new_n935));
  OAI221_X1 g0735(.A(new_n934), .B1(new_n483), .B2(new_n711), .C1(new_n724), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G317), .B2(new_n698), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n762), .A2(G294), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n930), .A2(new_n931), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n695), .A2(new_n216), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n711), .A2(new_n766), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n707), .A2(G143), .ZN(new_n942));
  INV_X1    g0742(.A(G137), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n697), .A2(new_n943), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n265), .B1(new_n702), .B2(new_n726), .C1(new_n319), .C2(new_n703), .ZN(new_n945));
  NOR4_X1   g0745(.A1(new_n941), .A2(new_n942), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n762), .A2(G159), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n720), .A2(G50), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n940), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n939), .A2(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n950), .A2(KEYINPUT47), .B1(new_n678), .B2(new_n679), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT47), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(new_n684), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n628), .B2(new_n409), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n233), .A2(new_n674), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n669), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n952), .B(new_n956), .C1(new_n686), .C2(new_n892), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n927), .A2(new_n957), .ZN(G387));
  OAI21_X1  g0758(.A(new_n921), .B1(new_n639), .B2(new_n662), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n922), .A2(new_n629), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n622), .A2(new_n686), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n348), .B1(new_n701), .B2(new_n216), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n408), .B2(new_n703), .ZN(new_n963));
  INV_X1    g0763(.A(new_n244), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n724), .A2(new_n337), .B1(new_n964), .B2(new_n712), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(G50), .C2(new_n710), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n720), .A2(G68), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n698), .A2(G150), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n966), .A2(new_n931), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G317), .A2(new_n710), .B1(new_n707), .B2(G322), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n761), .B2(new_n935), .C1(new_n483), .C2(new_n719), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT48), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  INV_X1    g0774(.A(new_n703), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n975), .A2(G283), .B1(new_n701), .B2(G294), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT49), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n265), .B1(new_n698), .B2(G326), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n694), .B2(new_n490), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT110), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n977), .B2(new_n978), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n969), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n680), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n627), .A2(new_n670), .B1(new_n418), .B2(new_n628), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n411), .A2(G50), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT50), .Z(new_n988));
  INV_X1    g0788(.A(G45), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n319), .B2(new_n321), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n988), .A2(new_n627), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n674), .B1(new_n230), .B2(new_n989), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n669), .B1(new_n993), .B2(new_n684), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n960), .B1(new_n666), .B2(new_n921), .C1(new_n961), .C2(new_n995), .ZN(G393));
  INV_X1    g0796(.A(new_n629), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n916), .A2(new_n924), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(new_n922), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(new_n925), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n265), .B1(new_n701), .B2(G283), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n723), .B(new_n1001), .C1(new_n709), .C2(new_n697), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT111), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G311), .A2(new_n710), .B1(new_n707), .B2(G317), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT52), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n720), .A2(G294), .B1(G116), .B2(new_n975), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n761), .B2(new_n483), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G150), .A2(new_n707), .B1(new_n710), .B2(G159), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT51), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n703), .A2(new_n321), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n265), .B1(new_n702), .B2(new_n319), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G143), .C2(new_n698), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n719), .B2(new_n411), .C1(new_n761), .C2(new_n202), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1010), .B(new_n1014), .C1(G87), .C2(new_n695), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n680), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n953), .B1(G97), .B2(new_n628), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n237), .A2(new_n674), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n669), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(new_n686), .C2(new_n896), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n998), .B2(new_n666), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1000), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G390));
  INV_X1    g0823(.A(KEYINPUT115), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n803), .B1(new_n327), .B2(new_n606), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n845), .A2(new_n849), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT113), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n789), .B1(new_n638), .B2(new_n745), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n802), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n851), .B(KEYINPUT112), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n867), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1026), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n865), .A2(G330), .A3(new_n802), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1027), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1024), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT113), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1039), .A2(KEYINPUT115), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n661), .A2(new_n618), .A3(new_n861), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(new_n802), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(G330), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n661), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n428), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n596), .B(new_n1047), .C1(new_n854), .C2(new_n855), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1042), .A2(new_n1028), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT116), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n661), .B2(new_n1045), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n749), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(KEYINPUT116), .B2(new_n1046), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1049), .B1(new_n1053), .B2(new_n802), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1041), .A2(new_n802), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n790), .B1(new_n1034), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1048), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1044), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT117), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1037), .A2(new_n1040), .A3(new_n1043), .A4(new_n1057), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(new_n629), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1044), .A2(new_n1058), .A3(KEYINPUT117), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n845), .A2(new_n681), .A3(new_n849), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n668), .B1(new_n754), .B2(new_n244), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n265), .B(new_n1011), .C1(G87), .C2(new_n701), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n490), .B2(new_n711), .C1(new_n928), .C2(new_n724), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G294), .B2(new_n698), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G97), .A2(new_n720), .B1(new_n762), .B2(G107), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n770), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(KEYINPUT54), .B(G143), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n720), .A2(new_n1074), .B1(G159), .B2(new_n975), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n761), .B2(new_n943), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT118), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n710), .A2(G132), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n707), .A2(G128), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n701), .A2(G150), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT53), .Z(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(G125), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n265), .B1(new_n1083), .B2(new_n697), .C1(new_n694), .C2(new_n202), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT119), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1072), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1067), .B1(new_n1086), .B2(new_n680), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1066), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1044), .B2(new_n666), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1065), .A2(new_n1090), .ZN(G378));
  AND2_X1   g0891(.A1(new_n261), .A2(new_n806), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT55), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n290), .B(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1096));
  AND2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n681), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n668), .B1(new_n754), .B2(G50), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n724), .A2(new_n490), .B1(new_n495), .B2(new_n712), .ZN(new_n1102));
  AOI211_X1 g0902(.A(G41), .B(new_n265), .C1(new_n701), .C2(new_n216), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n319), .B2(new_n703), .C1(new_n711), .C2(new_n418), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(G283), .C2(new_n698), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n695), .A2(G58), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n408), .C2(new_n719), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT58), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n202), .B1(new_n343), .B2(G41), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n975), .A2(G150), .B1(new_n701), .B2(new_n1074), .ZN(new_n1112));
  INV_X1    g0912(.A(G132), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n712), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n710), .A2(G128), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n724), .B2(new_n1083), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(new_n720), .C2(G137), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT59), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n695), .A2(G159), .ZN(new_n1121));
  AOI211_X1 g0921(.A(G33), .B(G41), .C1(new_n698), .C2(G124), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1101), .B1(new_n1124), .B2(new_n680), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1100), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n860), .A2(new_n866), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n868), .A2(KEYINPUT40), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(G330), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1099), .B1(new_n869), .B2(new_n1045), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n850), .A2(new_n851), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n825), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n852), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1127), .B1(new_n1139), .B2(new_n667), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1048), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1062), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1139), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n852), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1136), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1138), .A2(KEYINPUT121), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n997), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(KEYINPUT122), .B(new_n1141), .C1(new_n1146), .C2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT122), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1062), .A2(new_n1142), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n629), .C1(KEYINPUT57), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1154), .B1(new_n1157), .B2(new_n1140), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1153), .A2(new_n1158), .ZN(G375));
  NAND2_X1  g0959(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n802), .A2(new_n682), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT123), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n695), .A2(G77), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n348), .B1(new_n702), .B2(new_n495), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n409), .B2(new_n975), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n724), .B2(new_n431), .C1(new_n928), .C2(new_n711), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n719), .A2(new_n418), .B1(new_n761), .B2(new_n490), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G303), .C2(new_n698), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n265), .B1(new_n702), .B2(new_n337), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G50), .B2(new_n975), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n724), .B2(new_n1113), .C1(new_n943), .C2(new_n711), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n719), .A2(new_n766), .B1(new_n761), .B2(new_n1073), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G128), .C2(new_n698), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1163), .A2(new_n1168), .B1(new_n1173), .B2(new_n1106), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n678), .B2(new_n679), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n669), .B(new_n1175), .C1(new_n319), .C2(new_n753), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1160), .A2(new_n667), .B1(new_n1162), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n904), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1058), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1160), .A2(new_n1142), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(G381));
  NAND2_X1  g0981(.A1(new_n1062), .A2(new_n629), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1089), .B1(new_n1183), .B2(new_n1064), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n927), .A2(new_n1022), .A3(new_n957), .ZN(new_n1186));
  OR4_X1    g0986(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1187));
  OR3_X1    g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(G407));
  OAI211_X1 g0988(.A(G407), .B(G213), .C1(G343), .C2(new_n1185), .ZN(G409));
  NAND2_X1  g0989(.A1(new_n605), .A2(G213), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1156), .A2(new_n1178), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n852), .A2(new_n1132), .A3(new_n1133), .A4(new_n1148), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1137), .A2(new_n1150), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT124), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n666), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1149), .A2(KEYINPUT124), .A3(new_n1150), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1127), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1065), .A2(new_n1090), .A3(new_n1191), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1141), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1190), .B(new_n1198), .C1(new_n1199), .C2(new_n1184), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1180), .B1(new_n1058), .B2(KEYINPUT60), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1054), .A2(KEYINPUT60), .A3(new_n1048), .A4(new_n1056), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n629), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1177), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n778), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G384), .B(new_n1177), .C1(new_n1201), .C2(new_n1203), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT62), .B1(new_n1200), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n605), .A2(G213), .A3(G2897), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1205), .A2(new_n1206), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT61), .B1(new_n1200), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1198), .A2(new_n1190), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT62), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1207), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1155), .A2(new_n629), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1143), .B2(new_n1139), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1140), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(G378), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1208), .A2(new_n1213), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1022), .B1(new_n927), .B2(new_n957), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(G393), .B(G396), .Z(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1186), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1186), .ZN(new_n1229));
  OAI211_X1 g1029(.A(KEYINPUT125), .B(new_n1225), .C1(new_n1229), .C2(new_n1223), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT126), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1222), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1200), .B2(new_n1207), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1214), .A2(KEYINPUT63), .A3(new_n1216), .A4(new_n1220), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1231), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n1213), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(G405));
  NAND2_X1  g1042(.A1(new_n1231), .A2(new_n1216), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1228), .A2(new_n1230), .A3(new_n1207), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1219), .A2(KEYINPUT122), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1157), .A2(new_n1154), .A3(new_n1140), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G378), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1220), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1248), .A2(KEYINPUT127), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT127), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1185), .B2(new_n1220), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT127), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1185), .A2(new_n1251), .A3(new_n1220), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1244), .A4(new_n1243), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(G402));
endmodule


