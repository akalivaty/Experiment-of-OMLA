

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761;

  AND2_X1 U376 ( .A1(n608), .A2(n607), .ZN(n623) );
  AND2_X2 U377 ( .A1(n757), .A2(n601), .ZN(n605) );
  NAND2_X1 U378 ( .A1(n614), .A2(n588), .ZN(n399) );
  XNOR2_X1 U379 ( .A(n399), .B(KEYINPUT22), .ZN(n592) );
  XNOR2_X2 U380 ( .A(n498), .B(n497), .ZN(n533) );
  XNOR2_X2 U381 ( .A(n743), .B(G146), .ZN(n374) );
  NOR2_X1 U382 ( .A1(n565), .A2(n761), .ZN(n566) );
  AND2_X1 U383 ( .A1(n386), .A2(n626), .ZN(n625) );
  XNOR2_X1 U384 ( .A(n624), .B(KEYINPUT45), .ZN(n386) );
  XNOR2_X1 U385 ( .A(n404), .B(n403), .ZN(n565) );
  XNOR2_X1 U386 ( .A(n502), .B(KEYINPUT80), .ZN(n659) );
  XNOR2_X1 U387 ( .A(n564), .B(n369), .ZN(n761) );
  AND2_X1 U388 ( .A1(n401), .A2(n370), .ZN(n551) );
  NOR2_X1 U389 ( .A1(n674), .A2(n679), .ZN(n562) );
  NAND2_X1 U390 ( .A1(n433), .A2(n432), .ZN(n431) );
  XNOR2_X2 U391 ( .A(n400), .B(n459), .ZN(n743) );
  XNOR2_X2 U392 ( .A(n491), .B(n535), .ZN(n400) );
  INV_X1 U393 ( .A(KEYINPUT84), .ZN(n384) );
  XNOR2_X1 U394 ( .A(n570), .B(n569), .ZN(n385) );
  NOR2_X1 U395 ( .A1(n690), .A2(n397), .ZN(n402) );
  INV_X1 U396 ( .A(KEYINPUT70), .ZN(n528) );
  XNOR2_X1 U397 ( .A(n690), .B(KEYINPUT6), .ZN(n597) );
  XNOR2_X1 U398 ( .A(n526), .B(n525), .ZN(n559) );
  AND2_X1 U399 ( .A1(n482), .A2(n481), .ZN(n563) );
  NOR2_X1 U400 ( .A1(n690), .A2(n363), .ZN(n423) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n505) );
  XNOR2_X1 U402 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n504) );
  OR2_X1 U403 ( .A1(n576), .A2(n384), .ZN(n379) );
  AND2_X1 U404 ( .A1(n576), .A2(n384), .ZN(n381) );
  XNOR2_X1 U405 ( .A(KEYINPUT4), .B(G131), .ZN(n459) );
  NOR2_X1 U406 ( .A1(G237), .A2(G953), .ZN(n460) );
  XNOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT72), .ZN(n439) );
  XNOR2_X1 U408 ( .A(n476), .B(G107), .ZN(n484) );
  XNOR2_X1 U409 ( .A(G110), .B(G104), .ZN(n476) );
  XOR2_X1 U410 ( .A(G137), .B(G140), .Z(n474) );
  XNOR2_X1 U411 ( .A(n372), .B(KEYINPUT94), .ZN(n371) );
  INV_X1 U412 ( .A(G101), .ZN(n372) );
  NAND2_X1 U413 ( .A1(n387), .A2(n396), .ZN(n395) );
  XNOR2_X1 U414 ( .A(n450), .B(n449), .ZN(n541) );
  NOR2_X1 U415 ( .A1(n721), .A2(G902), .ZN(n450) );
  XNOR2_X1 U416 ( .A(G113), .B(KEYINPUT90), .ZN(n464) );
  XNOR2_X1 U417 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n461) );
  XNOR2_X1 U418 ( .A(G119), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U419 ( .A(G116), .B(G107), .ZN(n521) );
  XNOR2_X1 U420 ( .A(G122), .B(KEYINPUT9), .ZN(n518) );
  XNOR2_X1 U421 ( .A(n438), .B(n437), .ZN(n522) );
  XNOR2_X1 U422 ( .A(n405), .B(KEYINPUT39), .ZN(n536) );
  XNOR2_X1 U423 ( .A(n434), .B(n361), .ZN(n433) );
  AND2_X1 U424 ( .A1(n393), .A2(n676), .ZN(n392) );
  NOR2_X1 U425 ( .A1(n679), .A2(n587), .ZN(n588) );
  INV_X1 U426 ( .A(n559), .ZN(n549) );
  OR2_X1 U427 ( .A1(n630), .A2(G902), .ZN(n473) );
  INV_X1 U428 ( .A(KEYINPUT85), .ZN(n366) );
  NAND2_X1 U429 ( .A1(n422), .A2(n421), .ZN(n538) );
  NOR2_X1 U430 ( .A1(n675), .A2(n362), .ZN(n422) );
  INV_X1 U431 ( .A(n659), .ZN(n421) );
  OR2_X1 U432 ( .A1(n659), .A2(n675), .ZN(n553) );
  INV_X1 U433 ( .A(G237), .ZN(n496) );
  INV_X1 U434 ( .A(KEYINPUT3), .ZN(n465) );
  INV_X1 U435 ( .A(G953), .ZN(n730) );
  XNOR2_X1 U436 ( .A(n503), .B(G140), .ZN(n507) );
  XOR2_X1 U437 ( .A(KEYINPUT99), .B(G143), .Z(n503) );
  XNOR2_X1 U438 ( .A(G113), .B(G104), .ZN(n511) );
  XOR2_X1 U439 ( .A(G131), .B(G122), .Z(n512) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n487) );
  XOR2_X1 U441 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n488) );
  XOR2_X1 U442 ( .A(G125), .B(G146), .Z(n490) );
  AND2_X1 U443 ( .A1(n597), .A2(n540), .ZN(n544) );
  XNOR2_X1 U444 ( .A(n574), .B(KEYINPUT38), .ZN(n677) );
  NAND2_X1 U445 ( .A1(n544), .A2(n394), .ZN(n411) );
  NAND2_X1 U446 ( .A1(n364), .A2(n458), .ZN(n363) );
  NAND2_X1 U447 ( .A1(n380), .A2(n359), .ZN(n378) );
  XOR2_X1 U448 ( .A(G122), .B(KEYINPUT16), .Z(n483) );
  XNOR2_X1 U449 ( .A(n475), .B(n478), .ZN(n435) );
  XNOR2_X1 U450 ( .A(n474), .B(n371), .ZN(n475) );
  AND2_X1 U451 ( .A1(n408), .A2(n684), .ZN(n376) );
  NOR2_X1 U452 ( .A1(n411), .A2(n407), .ZN(n406) );
  INV_X1 U453 ( .A(n545), .ZN(n407) );
  NOR2_X1 U454 ( .A1(n354), .A2(n611), .ZN(n370) );
  XNOR2_X1 U455 ( .A(n402), .B(n360), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n368), .B(G475), .ZN(n367) );
  INV_X1 U457 ( .A(KEYINPUT13), .ZN(n368) );
  NAND2_X1 U458 ( .A1(n391), .A2(n390), .ZN(n586) );
  NAND2_X1 U459 ( .A1(n394), .A2(n357), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n374), .B(n470), .ZN(n630) );
  BUF_X1 U461 ( .A(n745), .Z(n373) );
  XNOR2_X1 U462 ( .A(n424), .B(n741), .ZN(n721) );
  XNOR2_X1 U463 ( .A(n443), .B(n425), .ZN(n424) );
  XNOR2_X1 U464 ( .A(n442), .B(n426), .ZN(n425) );
  INV_X1 U465 ( .A(G217), .ZN(n419) );
  XNOR2_X1 U466 ( .A(n523), .B(n416), .ZN(n719) );
  XNOR2_X1 U467 ( .A(n418), .B(n417), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n521), .B(KEYINPUT101), .ZN(n417) );
  INV_X1 U469 ( .A(KEYINPUT42), .ZN(n369) );
  INV_X1 U470 ( .A(G134), .ZN(n535) );
  INV_X1 U471 ( .A(KEYINPUT40), .ZN(n403) );
  INV_X1 U472 ( .A(KEYINPUT35), .ZN(n430) );
  INV_X1 U473 ( .A(n600), .ZN(n432) );
  NOR2_X1 U474 ( .A1(n687), .A2(n589), .ZN(n591) );
  NAND2_X1 U475 ( .A1(n398), .A2(n358), .ZN(n589) );
  NAND2_X1 U476 ( .A1(n559), .A2(n412), .ZN(n542) );
  INV_X1 U477 ( .A(n542), .ZN(n663) );
  NAND2_X1 U478 ( .A1(n619), .A2(n687), .ZN(n650) );
  AND2_X1 U479 ( .A1(n365), .A2(n546), .ZN(n618) );
  NOR2_X1 U480 ( .A1(G953), .A2(n709), .ZN(n710) );
  XNOR2_X1 U481 ( .A(n413), .B(KEYINPUT118), .ZN(n709) );
  OR2_X1 U482 ( .A1(n532), .A2(n531), .ZN(n354) );
  XNOR2_X1 U483 ( .A(n517), .B(n367), .ZN(n560) );
  INV_X1 U484 ( .A(n560), .ZN(n412) );
  XOR2_X1 U485 ( .A(KEYINPUT74), .B(KEYINPUT24), .Z(n355) );
  NAND2_X1 U486 ( .A1(n389), .A2(n388), .ZN(n584) );
  NOR2_X1 U487 ( .A1(n629), .A2(n419), .ZN(n356) );
  BUF_X1 U488 ( .A(n533), .Z(n574) );
  BUF_X1 U489 ( .A(n541), .Z(n687) );
  INV_X1 U490 ( .A(n541), .ZN(n364) );
  AND2_X1 U491 ( .A1(n583), .A2(n392), .ZN(n357) );
  NOR2_X1 U492 ( .A1(n597), .A2(n546), .ZN(n358) );
  AND2_X1 U493 ( .A1(n379), .A2(n383), .ZN(n359) );
  XNOR2_X1 U494 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n360) );
  XNOR2_X1 U495 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n361) );
  INV_X1 U496 ( .A(n676), .ZN(n397) );
  XOR2_X1 U497 ( .A(KEYINPUT71), .B(KEYINPUT47), .Z(n362) );
  XNOR2_X1 U498 ( .A(n617), .B(n366), .ZN(n365) );
  NOR2_X2 U499 ( .A1(n378), .A2(n382), .ZN(n744) );
  XOR2_X1 U500 ( .A(KEYINPUT105), .B(n552), .Z(n756) );
  NOR2_X1 U501 ( .A1(n375), .A2(n409), .ZN(n547) );
  XNOR2_X1 U502 ( .A(n374), .B(n435), .ZN(n711) );
  XNOR2_X2 U503 ( .A(n473), .B(n472), .ZN(n690) );
  NAND2_X1 U504 ( .A1(n377), .A2(n376), .ZN(n375) );
  OR2_X1 U505 ( .A1(n410), .A2(n545), .ZN(n377) );
  NAND2_X1 U506 ( .A1(n385), .A2(n381), .ZN(n380) );
  NOR2_X1 U507 ( .A1(n385), .A2(n384), .ZN(n382) );
  INV_X1 U508 ( .A(n577), .ZN(n383) );
  NAND2_X1 U509 ( .A1(n744), .A2(n386), .ZN(n672) );
  NAND2_X1 U510 ( .A1(n386), .A2(n730), .ZN(n731) );
  NAND2_X1 U511 ( .A1(n533), .A2(n501), .ZN(n387) );
  NAND2_X1 U512 ( .A1(n394), .A2(n392), .ZN(n388) );
  INV_X1 U513 ( .A(n395), .ZN(n389) );
  NAND2_X1 U514 ( .A1(n395), .A2(n583), .ZN(n391) );
  INV_X1 U515 ( .A(n501), .ZN(n393) );
  INV_X1 U516 ( .A(n533), .ZN(n394) );
  NAND2_X1 U517 ( .A1(n397), .A2(n501), .ZN(n396) );
  NOR2_X1 U518 ( .A1(n592), .A2(n597), .ZN(n617) );
  INV_X1 U519 ( .A(n592), .ZN(n398) );
  XNOR2_X1 U520 ( .A(n400), .B(n520), .ZN(n418) );
  INV_X1 U521 ( .A(n690), .ZN(n594) );
  NAND2_X1 U522 ( .A1(n536), .A2(n663), .ZN(n404) );
  NAND2_X1 U523 ( .A1(n551), .A2(n677), .ZN(n405) );
  NOR2_X1 U524 ( .A1(n672), .A2(n415), .ZN(n629) );
  NAND2_X1 U525 ( .A1(n420), .A2(n356), .ZN(n722) );
  NOR2_X1 U526 ( .A1(n724), .A2(n723), .ZN(n725) );
  INV_X1 U527 ( .A(n411), .ZN(n410) );
  AND2_X1 U528 ( .A1(n543), .A2(n406), .ZN(n409) );
  OR2_X1 U529 ( .A1(n543), .A2(n545), .ZN(n408) );
  NAND2_X1 U530 ( .A1(n543), .A2(n544), .ZN(n571) );
  NAND2_X1 U531 ( .A1(n414), .A2(n436), .ZN(n413) );
  XNOR2_X1 U532 ( .A(n672), .B(n415), .ZN(n414) );
  INV_X1 U533 ( .A(KEYINPUT2), .ZN(n415) );
  NOR2_X2 U534 ( .A1(n428), .A2(n629), .ZN(n717) );
  INV_X1 U535 ( .A(n428), .ZN(n420) );
  NAND2_X1 U536 ( .A1(n717), .A2(G472), .ZN(n632) );
  NAND2_X1 U537 ( .A1(n717), .A2(G210), .ZN(n639) );
  NAND2_X1 U538 ( .A1(n717), .A2(G475), .ZN(n645) );
  XNOR2_X1 U539 ( .A(n423), .B(KEYINPUT28), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n427), .A2(n628), .ZN(n429) );
  NAND2_X1 U541 ( .A1(n625), .A2(n744), .ZN(n427) );
  XNOR2_X1 U542 ( .A(n429), .B(KEYINPUT65), .ZN(n428) );
  XNOR2_X2 U543 ( .A(n431), .B(n430), .ZN(n757) );
  NAND2_X1 U544 ( .A1(n682), .A2(n614), .ZN(n434) );
  XNOR2_X2 U545 ( .A(n599), .B(KEYINPUT33), .ZN(n682) );
  XNOR2_X1 U546 ( .A(n490), .B(n439), .ZN(n508) );
  XNOR2_X1 U547 ( .A(KEYINPUT117), .B(n708), .ZN(n436) );
  INV_X1 U548 ( .A(KEYINPUT48), .ZN(n569) );
  XNOR2_X1 U549 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U550 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n585) );
  XOR2_X2 U551 ( .A(KEYINPUT64), .B(G953), .Z(n745) );
  NAND2_X1 U552 ( .A1(n745), .A2(G234), .ZN(n438) );
  XNOR2_X1 U553 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n437) );
  NAND2_X1 U554 ( .A1(n522), .A2(G221), .ZN(n443) );
  INV_X1 U555 ( .A(n508), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n474), .B(n440), .ZN(n741) );
  XNOR2_X1 U557 ( .A(G128), .B(G110), .ZN(n441) );
  XNOR2_X1 U558 ( .A(n355), .B(n441), .ZN(n442) );
  XOR2_X1 U559 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n447) );
  XNOR2_X1 U560 ( .A(G902), .B(KEYINPUT89), .ZN(n445) );
  INV_X1 U561 ( .A(KEYINPUT15), .ZN(n444) );
  XNOR2_X1 U562 ( .A(n445), .B(n444), .ZN(n578) );
  NAND2_X1 U563 ( .A1(G234), .A2(n578), .ZN(n446) );
  XNOR2_X1 U564 ( .A(n447), .B(n446), .ZN(n451) );
  NAND2_X1 U565 ( .A1(n451), .A2(G217), .ZN(n448) );
  XNOR2_X1 U566 ( .A(n448), .B(KEYINPUT25), .ZN(n449) );
  NAND2_X1 U567 ( .A1(n451), .A2(G221), .ZN(n453) );
  INV_X1 U568 ( .A(KEYINPUT21), .ZN(n452) );
  XNOR2_X1 U569 ( .A(n453), .B(n452), .ZN(n688) );
  NOR2_X1 U570 ( .A1(n373), .A2(G900), .ZN(n454) );
  NAND2_X1 U571 ( .A1(G902), .A2(n454), .ZN(n455) );
  NAND2_X1 U572 ( .A1(G952), .A2(n730), .ZN(n580) );
  NAND2_X1 U573 ( .A1(n455), .A2(n580), .ZN(n457) );
  NAND2_X1 U574 ( .A1(G237), .A2(G234), .ZN(n456) );
  XNOR2_X1 U575 ( .A(n456), .B(KEYINPUT14), .ZN(n673) );
  AND2_X1 U576 ( .A1(n457), .A2(n673), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n688), .A2(n530), .ZN(n539) );
  INV_X1 U578 ( .A(n539), .ZN(n458) );
  XNOR2_X2 U579 ( .A(G143), .B(G128), .ZN(n491) );
  XNOR2_X1 U580 ( .A(n460), .B(KEYINPUT78), .ZN(n510) );
  NAND2_X1 U581 ( .A1(n510), .A2(G210), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n461), .B(G137), .ZN(n462) );
  XNOR2_X1 U583 ( .A(n463), .B(n462), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n464), .B(G101), .ZN(n468) );
  XNOR2_X1 U585 ( .A(G119), .B(G116), .ZN(n466) );
  XNOR2_X1 U586 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U587 ( .A(n468), .B(n467), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n486), .B(n469), .ZN(n470) );
  INV_X1 U589 ( .A(KEYINPUT76), .ZN(n471) );
  XNOR2_X1 U590 ( .A(n471), .B(G472), .ZN(n472) );
  NAND2_X1 U591 ( .A1(G227), .A2(n745), .ZN(n477) );
  XNOR2_X1 U592 ( .A(n484), .B(n477), .ZN(n478) );
  NOR2_X1 U593 ( .A1(n711), .A2(G902), .ZN(n480) );
  XNOR2_X1 U594 ( .A(KEYINPUT73), .B(G469), .ZN(n479) );
  XNOR2_X2 U595 ( .A(n480), .B(n479), .ZN(n609) );
  XNOR2_X1 U596 ( .A(n609), .B(KEYINPUT106), .ZN(n481) );
  XNOR2_X1 U597 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n486), .B(n485), .ZN(n726) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U600 ( .A(n490), .B(n489), .ZN(n494) );
  NAND2_X1 U601 ( .A1(G224), .A2(n745), .ZN(n492) );
  XNOR2_X1 U602 ( .A(n491), .B(n492), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U604 ( .A(n726), .B(n495), .ZN(n637) );
  NAND2_X1 U605 ( .A1(n637), .A2(n578), .ZN(n498) );
  INV_X1 U606 ( .A(G902), .ZN(n524) );
  NAND2_X1 U607 ( .A1(n524), .A2(n496), .ZN(n499) );
  NAND2_X1 U608 ( .A1(n499), .A2(G210), .ZN(n497) );
  NAND2_X1 U609 ( .A1(n499), .A2(G214), .ZN(n676) );
  INV_X1 U610 ( .A(KEYINPUT79), .ZN(n500) );
  XNOR2_X1 U611 ( .A(n500), .B(KEYINPUT19), .ZN(n501) );
  NAND2_X1 U612 ( .A1(n563), .A2(n584), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n509), .B(n440), .ZN(n516) );
  NAND2_X1 U615 ( .A1(n510), .A2(G214), .ZN(n514) );
  XNOR2_X1 U616 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n643) );
  NOR2_X1 U619 ( .A1(G902), .A2(n643), .ZN(n517) );
  XOR2_X1 U620 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n519) );
  XNOR2_X1 U621 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U622 ( .A1(n522), .A2(G217), .ZN(n523) );
  NAND2_X1 U623 ( .A1(n719), .A2(n524), .ZN(n526) );
  INV_X1 U624 ( .A(G478), .ZN(n525) );
  NOR2_X1 U625 ( .A1(n659), .A2(n542), .ZN(n527) );
  XOR2_X1 U626 ( .A(G146), .B(n527), .Z(G48) );
  NAND2_X1 U627 ( .A1(n541), .A2(n688), .ZN(n529) );
  XNOR2_X2 U628 ( .A(n529), .B(n528), .ZN(n685) );
  INV_X1 U629 ( .A(n685), .ZN(n611) );
  INV_X1 U630 ( .A(n609), .ZN(n532) );
  INV_X1 U631 ( .A(n530), .ZN(n531) );
  INV_X1 U632 ( .A(n536), .ZN(n534) );
  AND2_X1 U633 ( .A1(n560), .A2(n549), .ZN(n667) );
  INV_X1 U634 ( .A(n667), .ZN(n658) );
  NOR2_X1 U635 ( .A1(n534), .A2(n658), .ZN(n577) );
  XNOR2_X1 U636 ( .A(n577), .B(n535), .ZN(G36) );
  XOR2_X1 U637 ( .A(G131), .B(n565), .Z(G33) );
  NOR2_X1 U638 ( .A1(n663), .A2(n667), .ZN(n537) );
  XNOR2_X1 U639 ( .A(n537), .B(KEYINPUT102), .ZN(n675) );
  XNOR2_X1 U640 ( .A(n538), .B(KEYINPUT77), .ZN(n548) );
  NOR2_X1 U641 ( .A1(n539), .A2(n397), .ZN(n540) );
  NOR2_X1 U642 ( .A1(n687), .A2(n542), .ZN(n543) );
  XNOR2_X1 U643 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n545) );
  XNOR2_X2 U644 ( .A(n609), .B(KEYINPUT1), .ZN(n684) );
  INV_X1 U645 ( .A(n684), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n547), .B(KEYINPUT108), .ZN(n759) );
  NOR2_X1 U647 ( .A1(n548), .A2(n759), .ZN(n558) );
  NAND2_X1 U648 ( .A1(n412), .A2(n549), .ZN(n600) );
  NOR2_X1 U649 ( .A1(n600), .A2(n574), .ZN(n550) );
  NAND2_X1 U650 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U651 ( .A(n756), .B(KEYINPUT82), .ZN(n555) );
  NAND2_X1 U652 ( .A1(n553), .A2(KEYINPUT47), .ZN(n554) );
  NAND2_X1 U653 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U654 ( .A(n556), .B(KEYINPUT81), .ZN(n557) );
  AND2_X1 U655 ( .A1(n558), .A2(n557), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n677), .A2(n676), .ZN(n674) );
  NAND2_X1 U657 ( .A1(n560), .A2(n559), .ZN(n679) );
  XNOR2_X1 U658 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n561) );
  XNOR2_X1 U659 ( .A(n562), .B(n561), .ZN(n697) );
  NAND2_X1 U660 ( .A1(n697), .A2(n563), .ZN(n564) );
  XNOR2_X1 U661 ( .A(KEYINPUT46), .B(n566), .ZN(n567) );
  NAND2_X1 U662 ( .A1(n568), .A2(n567), .ZN(n570) );
  NOR2_X1 U663 ( .A1(n684), .A2(n571), .ZN(n573) );
  XNOR2_X1 U664 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n572) );
  XOR2_X1 U665 ( .A(n573), .B(n572), .Z(n575) );
  NOR2_X1 U666 ( .A1(n575), .A2(n394), .ZN(n671) );
  INV_X1 U667 ( .A(n671), .ZN(n576) );
  INV_X1 U668 ( .A(n578), .ZN(n626) );
  XOR2_X1 U669 ( .A(G898), .B(KEYINPUT92), .Z(n733) );
  NAND2_X1 U670 ( .A1(n733), .A2(G953), .ZN(n579) );
  XNOR2_X1 U671 ( .A(n579), .B(KEYINPUT93), .ZN(n728) );
  NAND2_X1 U672 ( .A1(n728), .A2(G902), .ZN(n581) );
  NAND2_X1 U673 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U674 ( .A1(n582), .A2(n673), .ZN(n583) );
  XNOR2_X2 U675 ( .A(n586), .B(n585), .ZN(n614) );
  INV_X1 U676 ( .A(n688), .ZN(n587) );
  XNOR2_X1 U677 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n590) );
  XNOR2_X1 U678 ( .A(n591), .B(n590), .ZN(n754) );
  NOR2_X1 U679 ( .A1(n592), .A2(n684), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n364), .A2(n593), .ZN(n595) );
  NOR2_X1 U681 ( .A1(n595), .A2(n594), .ZN(n656) );
  NOR2_X1 U682 ( .A1(n754), .A2(n656), .ZN(n604) );
  INV_X1 U683 ( .A(KEYINPUT44), .ZN(n596) );
  AND2_X1 U684 ( .A1(n604), .A2(n596), .ZN(n603) );
  INV_X1 U685 ( .A(KEYINPUT69), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n685), .A2(n684), .ZN(n613) );
  INV_X1 U687 ( .A(n613), .ZN(n598) );
  NAND2_X1 U688 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U689 ( .A(n601), .B(n757), .ZN(n602) );
  NAND2_X1 U690 ( .A1(n603), .A2(n602), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n606), .A2(KEYINPUT44), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n609), .A2(n690), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U695 ( .A1(n614), .A2(n612), .ZN(n652) );
  NOR2_X1 U696 ( .A1(n613), .A2(n690), .ZN(n695) );
  NAND2_X1 U697 ( .A1(n614), .A2(n695), .ZN(n615) );
  XNOR2_X1 U698 ( .A(KEYINPUT31), .B(n615), .ZN(n668) );
  NOR2_X1 U699 ( .A1(n652), .A2(n668), .ZN(n616) );
  NOR2_X1 U700 ( .A1(n675), .A2(n616), .ZN(n621) );
  XNOR2_X1 U701 ( .A(n618), .B(KEYINPUT86), .ZN(n619) );
  INV_X1 U702 ( .A(n650), .ZN(n620) );
  NOR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  XOR2_X1 U706 ( .A(KEYINPUT67), .B(n627), .Z(n628) );
  XOR2_X1 U707 ( .A(KEYINPUT62), .B(n630), .Z(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n373), .A2(G952), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(KEYINPUT88), .ZN(n724) );
  INV_X1 U711 ( .A(n724), .ZN(n646) );
  NAND2_X1 U712 ( .A1(n634), .A2(n646), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n635), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n636) );
  XNOR2_X1 U715 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n640), .A2(n646), .ZN(n642) );
  INV_X1 U718 ( .A(KEYINPUT56), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n642), .B(n641), .ZN(G51) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT59), .ZN(n644) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n649) );
  INV_X1 U723 ( .A(KEYINPUT60), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(G60) );
  XNOR2_X1 U725 ( .A(G101), .B(n650), .ZN(G3) );
  NAND2_X1 U726 ( .A1(n652), .A2(n663), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(G104), .ZN(G6) );
  XOR2_X1 U728 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n654) );
  NAND2_X1 U729 ( .A1(n652), .A2(n667), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(G107), .B(n655), .ZN(G9) );
  XNOR2_X1 U732 ( .A(G110), .B(n656), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT109), .ZN(G12) );
  NOR2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U735 ( .A(KEYINPUT29), .B(KEYINPUT110), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U737 ( .A(G128), .B(n662), .ZN(G30) );
  XOR2_X1 U738 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n665) );
  NAND2_X1 U739 ( .A1(n668), .A2(n663), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U741 ( .A(G113), .B(n666), .ZN(G15) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n669), .B(KEYINPUT114), .ZN(n670) );
  XNOR2_X1 U744 ( .A(G116), .B(n670), .ZN(G18) );
  XOR2_X1 U745 ( .A(G140), .B(n671), .Z(G42) );
  NAND2_X1 U746 ( .A1(n682), .A2(n697), .ZN(n707) );
  INV_X1 U747 ( .A(n673), .ZN(n704) );
  NOR2_X1 U748 ( .A1(n675), .A2(n674), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U754 ( .A(n686), .B(KEYINPUT50), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n689), .B(KEYINPUT49), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(n696), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U763 ( .A(n701), .B(KEYINPUT52), .ZN(n702) );
  XOR2_X1 U764 ( .A(KEYINPUT116), .B(n702), .Z(n703) );
  NOR2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U766 ( .A1(n705), .A2(G952), .ZN(n706) );
  NAND2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(KEYINPUT53), .B(n710), .ZN(G75) );
  NAND2_X1 U769 ( .A1(n717), .A2(G469), .ZN(n715) );
  XNOR2_X1 U770 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n713) );
  XNOR2_X1 U771 ( .A(n711), .B(KEYINPUT57), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n724), .A2(n716), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n717), .A2(G478), .ZN(n718) );
  XOR2_X1 U776 ( .A(n719), .B(n718), .Z(n720) );
  NOR2_X1 U777 ( .A1(n724), .A2(n720), .ZN(G63) );
  XNOR2_X1 U778 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U779 ( .A(KEYINPUT120), .B(n725), .ZN(G66) );
  XNOR2_X1 U780 ( .A(KEYINPUT125), .B(KEYINPUT122), .ZN(n740) );
  XOR2_X1 U781 ( .A(n726), .B(KEYINPUT123), .Z(n727) );
  XNOR2_X1 U782 ( .A(KEYINPUT124), .B(n727), .ZN(n729) );
  NOR2_X1 U783 ( .A1(n729), .A2(n728), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT121), .ZN(n736) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n732) );
  XOR2_X1 U786 ( .A(KEYINPUT61), .B(n732), .Z(n734) );
  NOR2_X1 U787 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(G69) );
  XNOR2_X1 U791 ( .A(n741), .B(KEYINPUT94), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n744), .B(n747), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(n373), .ZN(n753) );
  XOR2_X1 U795 ( .A(KEYINPUT126), .B(n747), .Z(n748) );
  XNOR2_X1 U796 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U797 ( .A1(G900), .A2(n749), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT127), .B(n750), .Z(n751) );
  NAND2_X1 U799 ( .A1(n751), .A2(G953), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U801 ( .A(G119), .B(n754), .Z(G21) );
  XOR2_X1 U802 ( .A(G143), .B(KEYINPUT111), .Z(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(G45) );
  XNOR2_X1 U804 ( .A(n757), .B(G122), .ZN(G24) );
  XOR2_X1 U805 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n758) );
  XNOR2_X1 U806 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U807 ( .A(G125), .B(n760), .ZN(G27) );
  XOR2_X1 U808 ( .A(G137), .B(n761), .Z(G39) );
endmodule

