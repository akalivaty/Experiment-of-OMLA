

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756;

  NAND2_X1 U376 ( .A1(n505), .A2(n481), .ZN(n564) );
  NOR2_X2 U377 ( .A1(n499), .A2(n667), .ZN(n500) );
  INV_X1 U378 ( .A(n493), .ZN(n667) );
  NOR2_X1 U379 ( .A1(n713), .A2(n726), .ZN(n714) );
  XNOR2_X1 U380 ( .A(KEYINPUT3), .B(G119), .ZN(n421) );
  XNOR2_X1 U381 ( .A(KEYINPUT4), .B(G101), .ZN(n419) );
  XNOR2_X2 U382 ( .A(G902), .B(KEYINPUT15), .ZN(n608) );
  OR2_X1 U383 ( .A1(n717), .A2(G902), .ZN(n448) );
  XNOR2_X1 U384 ( .A(n458), .B(n474), .ZN(n438) );
  XNOR2_X1 U385 ( .A(n384), .B(KEYINPUT10), .ZN(n372) );
  XNOR2_X1 U386 ( .A(n539), .B(KEYINPUT41), .ZN(n699) );
  XNOR2_X1 U387 ( .A(n356), .B(KEYINPUT28), .ZN(n546) );
  AND2_X1 U388 ( .A1(n560), .A2(n354), .ZN(n356) );
  XNOR2_X1 U389 ( .A(n594), .B(n593), .ZN(n357) );
  AND2_X1 U390 ( .A1(n492), .A2(n484), .ZN(n666) );
  INV_X1 U391 ( .A(n492), .ZN(n670) );
  XNOR2_X1 U392 ( .A(n486), .B(n485), .ZN(n687) );
  AND2_X2 U393 ( .A1(n357), .A2(n607), .ZN(n745) );
  XNOR2_X1 U394 ( .A(n439), .B(n367), .ZN(n368) );
  XNOR2_X1 U395 ( .A(n376), .B(G107), .ZN(n459) );
  XNOR2_X1 U396 ( .A(G122), .B(G116), .ZN(n376) );
  XNOR2_X1 U397 ( .A(n475), .B(n359), .ZN(n476) );
  INV_X1 U398 ( .A(KEYINPUT64), .ZN(n362) );
  INV_X1 U399 ( .A(KEYINPUT93), .ZN(n437) );
  XNOR2_X1 U400 ( .A(n418), .B(G125), .ZN(n384) );
  OR2_X1 U401 ( .A1(n586), .A2(n686), .ZN(n556) );
  BUF_X1 U402 ( .A(n537), .Z(n599) );
  BUF_X1 U403 ( .A(n707), .Z(n722) );
  XNOR2_X1 U404 ( .A(n548), .B(n547), .ZN(n756) );
  XNOR2_X1 U405 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U406 ( .A(KEYINPUT102), .ZN(n450) );
  NOR2_X1 U407 ( .A1(n573), .A2(n572), .ZN(n651) );
  AND2_X1 U408 ( .A1(n491), .A2(n561), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n392), .B(n391), .ZN(n537) );
  INV_X1 U410 ( .A(G146), .ZN(n418) );
  NAND2_X1 U411 ( .A1(n355), .A2(n434), .ZN(n413) );
  XNOR2_X1 U412 ( .A(n619), .B(n355), .ZN(n620) );
  XNOR2_X1 U413 ( .A(n374), .B(n375), .ZN(n355) );
  NAND2_X1 U414 ( .A1(n357), .A2(n603), .ZN(n604) );
  XNOR2_X1 U415 ( .A(n438), .B(n437), .ZN(n742) );
  XNOR2_X1 U416 ( .A(n665), .B(KEYINPUT83), .ZN(n704) );
  XNOR2_X1 U417 ( .A(n369), .B(n368), .ZN(n375) );
  XNOR2_X1 U418 ( .A(n741), .B(n469), .ZN(n477) );
  XOR2_X1 U419 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n358) );
  XOR2_X1 U420 ( .A(n474), .B(G143), .Z(n359) );
  XOR2_X1 U421 ( .A(n401), .B(n400), .Z(n360) );
  NOR2_X1 U422 ( .A1(n625), .A2(n649), .ZN(n361) );
  INV_X1 U423 ( .A(n608), .ZN(n609) );
  INV_X1 U424 ( .A(KEYINPUT11), .ZN(n467) );
  XNOR2_X1 U425 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n420) );
  XNOR2_X1 U426 ( .A(n467), .B(G122), .ZN(n468) );
  INV_X1 U427 ( .A(KEYINPUT85), .ZN(n615) );
  XNOR2_X1 U428 ( .A(n468), .B(G140), .ZN(n469) );
  XNOR2_X1 U429 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U430 ( .A(KEYINPUT104), .ZN(n463) );
  XNOR2_X1 U431 ( .A(n438), .B(n431), .ZN(n432) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n456) );
  XNOR2_X1 U433 ( .A(n500), .B(n358), .ZN(n690) );
  XNOR2_X1 U434 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U435 ( .A(n536), .B(n535), .ZN(n614) );
  XNOR2_X1 U436 ( .A(n477), .B(n476), .ZN(n634) );
  NOR2_X1 U437 ( .A1(n687), .A2(n538), .ZN(n539) );
  XNOR2_X1 U438 ( .A(n479), .B(n478), .ZN(n504) );
  XNOR2_X1 U439 ( .A(n466), .B(n465), .ZN(n505) );
  BUF_X1 U440 ( .A(n614), .Z(n730) );
  XNOR2_X1 U441 ( .A(n453), .B(n452), .ZN(n659) );
  OR2_X1 U442 ( .A1(n363), .A2(G952), .ZN(n712) );
  XNOR2_X2 U443 ( .A(n362), .B(G953), .ZN(n363) );
  NAND2_X1 U444 ( .A1(n363), .A2(G234), .ZN(n365) );
  XNOR2_X1 U445 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n364) );
  NAND2_X1 U446 ( .A1(n456), .A2(G221), .ZN(n369) );
  XNOR2_X1 U447 ( .A(G140), .B(G137), .ZN(n739) );
  INV_X1 U448 ( .A(G110), .ZN(n366) );
  XNOR2_X1 U449 ( .A(n739), .B(n366), .ZN(n439) );
  XOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n367) );
  XOR2_X1 U451 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n371) );
  XNOR2_X1 U452 ( .A(G128), .B(G119), .ZN(n370) );
  XNOR2_X1 U453 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X2 U454 ( .A(n372), .B(KEYINPUT68), .ZN(n741) );
  XNOR2_X1 U455 ( .A(n373), .B(n741), .ZN(n374) );
  INV_X1 U456 ( .A(G113), .ZN(n377) );
  XNOR2_X1 U457 ( .A(n377), .B(G104), .ZN(n470) );
  XNOR2_X1 U458 ( .A(n459), .B(n470), .ZN(n380) );
  XNOR2_X1 U459 ( .A(G110), .B(KEYINPUT16), .ZN(n378) );
  XNOR2_X1 U460 ( .A(n421), .B(n378), .ZN(n379) );
  XNOR2_X1 U461 ( .A(n380), .B(n379), .ZN(n727) );
  NAND2_X1 U462 ( .A1(n363), .A2(G224), .ZN(n383) );
  XNOR2_X1 U463 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n381) );
  XNOR2_X1 U464 ( .A(n381), .B(KEYINPUT91), .ZN(n382) );
  XNOR2_X1 U465 ( .A(n383), .B(n382), .ZN(n387) );
  XNOR2_X1 U466 ( .A(G143), .B(G128), .ZN(n428) );
  XNOR2_X1 U467 ( .A(n428), .B(n419), .ZN(n385) );
  XNOR2_X1 U468 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U469 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U470 ( .A(n727), .B(n388), .ZN(n709) );
  NAND2_X1 U471 ( .A1(n709), .A2(n608), .ZN(n392) );
  INV_X1 U472 ( .A(G902), .ZN(n434) );
  INV_X1 U473 ( .A(G237), .ZN(n389) );
  NAND2_X1 U474 ( .A1(n434), .A2(n389), .ZN(n393) );
  NAND2_X1 U475 ( .A1(n393), .A2(G210), .ZN(n390) );
  XNOR2_X1 U476 ( .A(n390), .B(KEYINPUT81), .ZN(n391) );
  NAND2_X1 U477 ( .A1(n393), .A2(G214), .ZN(n684) );
  NAND2_X1 U478 ( .A1(n537), .A2(n684), .ZN(n395) );
  XNOR2_X1 U479 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n394) );
  XNOR2_X1 U480 ( .A(n395), .B(n394), .ZN(n572) );
  INV_X1 U481 ( .A(n572), .ZN(n402) );
  XOR2_X1 U482 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n397) );
  NAND2_X1 U483 ( .A1(G234), .A2(G237), .ZN(n396) );
  XNOR2_X1 U484 ( .A(n397), .B(n396), .ZN(n398) );
  NAND2_X1 U485 ( .A1(G952), .A2(n398), .ZN(n696) );
  OR2_X1 U486 ( .A1(n696), .A2(G953), .ZN(n542) );
  NAND2_X1 U487 ( .A1(G902), .A2(n398), .ZN(n540) );
  INV_X1 U488 ( .A(G898), .ZN(n733) );
  NAND2_X1 U489 ( .A1(G953), .A2(n733), .ZN(n728) );
  OR2_X1 U490 ( .A1(n540), .A2(n728), .ZN(n399) );
  NAND2_X1 U491 ( .A1(n542), .A2(n399), .ZN(n401) );
  INV_X1 U492 ( .A(KEYINPUT92), .ZN(n400) );
  NAND2_X1 U493 ( .A1(n402), .A2(n360), .ZN(n405) );
  XNOR2_X1 U494 ( .A(KEYINPUT90), .B(KEYINPUT0), .ZN(n403) );
  XNOR2_X1 U495 ( .A(n403), .B(KEYINPUT66), .ZN(n404) );
  XNOR2_X1 U496 ( .A(n405), .B(n404), .ZN(n454) );
  INV_X1 U497 ( .A(n454), .ZN(n501) );
  XOR2_X1 U498 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n409) );
  NAND2_X1 U499 ( .A1(n608), .A2(G234), .ZN(n406) );
  XNOR2_X1 U500 ( .A(n406), .B(KEYINPUT96), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n407), .B(KEYINPUT20), .ZN(n414) );
  NAND2_X1 U502 ( .A1(n414), .A2(G217), .ZN(n408) );
  XNOR2_X1 U503 ( .A(n409), .B(n408), .ZN(n411) );
  INV_X1 U504 ( .A(KEYINPUT97), .ZN(n410) );
  XNOR2_X1 U505 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U506 ( .A(n413), .B(n412), .ZN(n492) );
  AND2_X1 U507 ( .A1(n414), .A2(G221), .ZN(n417) );
  INV_X1 U508 ( .A(KEYINPUT98), .ZN(n415) );
  XNOR2_X1 U509 ( .A(n415), .B(KEYINPUT21), .ZN(n416) );
  XNOR2_X1 U510 ( .A(n417), .B(n416), .ZN(n671) );
  INV_X1 U511 ( .A(n671), .ZN(n484) );
  XNOR2_X1 U512 ( .A(n419), .B(G146), .ZN(n441) );
  XNOR2_X1 U513 ( .A(n441), .B(n420), .ZN(n427) );
  XOR2_X1 U514 ( .A(n421), .B(KEYINPUT101), .Z(n425) );
  XOR2_X1 U515 ( .A(KEYINPUT100), .B(G116), .Z(n423) );
  XNOR2_X1 U516 ( .A(G137), .B(G113), .ZN(n422) );
  XNOR2_X1 U517 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U518 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U519 ( .A(n427), .B(n426), .Z(n433) );
  XNOR2_X1 U520 ( .A(n428), .B(G134), .ZN(n458) );
  INV_X1 U521 ( .A(KEYINPUT69), .ZN(n429) );
  XNOR2_X1 U522 ( .A(n429), .B(G131), .ZN(n474) );
  NOR2_X1 U523 ( .A1(G237), .A2(G953), .ZN(n430) );
  XNOR2_X1 U524 ( .A(n430), .B(KEYINPUT76), .ZN(n471) );
  NAND2_X1 U525 ( .A1(G210), .A2(n471), .ZN(n431) );
  XNOR2_X1 U526 ( .A(n433), .B(n432), .ZN(n627) );
  NAND2_X1 U527 ( .A1(n627), .A2(n434), .ZN(n436) );
  XNOR2_X1 U528 ( .A(G472), .B(KEYINPUT72), .ZN(n435) );
  XNOR2_X2 U529 ( .A(n436), .B(n435), .ZN(n491) );
  NAND2_X1 U530 ( .A1(n666), .A2(n491), .ZN(n449) );
  INV_X1 U531 ( .A(n439), .ZN(n440) );
  XNOR2_X1 U532 ( .A(n441), .B(n440), .ZN(n446) );
  NAND2_X1 U533 ( .A1(n363), .A2(G227), .ZN(n444) );
  XNOR2_X1 U534 ( .A(G104), .B(G107), .ZN(n442) );
  XNOR2_X1 U535 ( .A(n442), .B(KEYINPUT79), .ZN(n443) );
  XNOR2_X1 U536 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U537 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U538 ( .A(n742), .B(n447), .ZN(n717) );
  XNOR2_X2 U539 ( .A(n448), .B(G469), .ZN(n545) );
  XNOR2_X2 U540 ( .A(n545), .B(KEYINPUT1), .ZN(n493) );
  NOR2_X1 U541 ( .A1(n449), .A2(n667), .ZN(n677) );
  NAND2_X1 U542 ( .A1(n501), .A2(n677), .ZN(n453) );
  XOR2_X1 U543 ( .A(KEYINPUT103), .B(KEYINPUT31), .Z(n451) );
  NAND2_X1 U544 ( .A1(n666), .A2(n545), .ZN(n550) );
  OR2_X1 U545 ( .A1(n550), .A2(n491), .ZN(n455) );
  OR2_X1 U546 ( .A1(n455), .A2(n454), .ZN(n643) );
  NAND2_X1 U547 ( .A1(n659), .A2(n643), .ZN(n482) );
  NAND2_X1 U548 ( .A1(n456), .A2(G217), .ZN(n457) );
  XNOR2_X1 U549 ( .A(n458), .B(n457), .ZN(n462) );
  XOR2_X1 U550 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n460) );
  XOR2_X1 U551 ( .A(n460), .B(n459), .Z(n461) );
  XNOR2_X1 U552 ( .A(n462), .B(n461), .ZN(n723) );
  NOR2_X1 U553 ( .A1(G902), .A2(n723), .ZN(n466) );
  INV_X1 U554 ( .A(G478), .ZN(n464) );
  XNOR2_X1 U555 ( .A(KEYINPUT13), .B(G475), .ZN(n479) );
  XOR2_X1 U556 ( .A(n470), .B(KEYINPUT12), .Z(n473) );
  NAND2_X1 U557 ( .A1(G214), .A2(n471), .ZN(n472) );
  XNOR2_X1 U558 ( .A(n473), .B(n472), .ZN(n475) );
  OR2_X1 U559 ( .A1(G902), .A2(n634), .ZN(n478) );
  INV_X1 U560 ( .A(n504), .ZN(n481) );
  NOR2_X1 U561 ( .A1(n505), .A2(n481), .ZN(n480) );
  XNOR2_X1 U562 ( .A(n480), .B(KEYINPUT105), .ZN(n658) );
  NAND2_X1 U563 ( .A1(n658), .A2(n564), .ZN(n682) );
  NAND2_X1 U564 ( .A1(n482), .A2(n682), .ZN(n483) );
  XNOR2_X1 U565 ( .A(n483), .B(KEYINPUT106), .ZN(n497) );
  NAND2_X1 U566 ( .A1(n501), .A2(n484), .ZN(n487) );
  NAND2_X1 U567 ( .A1(n505), .A2(n504), .ZN(n486) );
  INV_X1 U568 ( .A(KEYINPUT107), .ZN(n485) );
  NOR2_X1 U569 ( .A1(n487), .A2(n687), .ZN(n490) );
  INV_X1 U570 ( .A(KEYINPUT73), .ZN(n488) );
  XNOR2_X1 U571 ( .A(n488), .B(KEYINPUT22), .ZN(n489) );
  XNOR2_X1 U572 ( .A(n490), .B(n489), .ZN(n522) );
  XNOR2_X1 U573 ( .A(n491), .B(KEYINPUT6), .ZN(n565) );
  INV_X1 U574 ( .A(n670), .ZN(n544) );
  NAND2_X1 U575 ( .A1(n565), .A2(n544), .ZN(n494) );
  NOR2_X1 U576 ( .A1(n494), .A2(n493), .ZN(n495) );
  AND2_X1 U577 ( .A1(n522), .A2(n495), .ZN(n641) );
  INV_X1 U578 ( .A(n641), .ZN(n496) );
  AND2_X1 U579 ( .A1(n497), .A2(n496), .ZN(n513) );
  INV_X1 U580 ( .A(n565), .ZN(n498) );
  NAND2_X1 U581 ( .A1(n498), .A2(n666), .ZN(n499) );
  NAND2_X1 U582 ( .A1(n690), .A2(n501), .ZN(n503) );
  INV_X1 U583 ( .A(KEYINPUT34), .ZN(n502) );
  XNOR2_X1 U584 ( .A(n503), .B(n502), .ZN(n506) );
  NOR2_X1 U585 ( .A1(n505), .A2(n504), .ZN(n584) );
  NAND2_X1 U586 ( .A1(n506), .A2(n584), .ZN(n509) );
  XNOR2_X1 U587 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n507) );
  XNOR2_X1 U588 ( .A(n507), .B(KEYINPUT80), .ZN(n508) );
  XNOR2_X2 U589 ( .A(n509), .B(n508), .ZN(n640) );
  NAND2_X1 U590 ( .A1(n640), .A2(KEYINPUT44), .ZN(n510) );
  NAND2_X1 U591 ( .A1(n513), .A2(n510), .ZN(n511) );
  NAND2_X1 U592 ( .A1(n511), .A2(KEYINPUT89), .ZN(n515) );
  INV_X1 U593 ( .A(KEYINPUT89), .ZN(n512) );
  NAND2_X1 U594 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U595 ( .A1(n515), .A2(n514), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n565), .A2(n670), .ZN(n516) );
  NOR2_X1 U597 ( .A1(n516), .A2(n667), .ZN(n517) );
  NAND2_X1 U598 ( .A1(n522), .A2(n517), .ZN(n519) );
  INV_X1 U599 ( .A(KEYINPUT32), .ZN(n518) );
  XNOR2_X1 U600 ( .A(n519), .B(n518), .ZN(n625) );
  OR2_X1 U601 ( .A1(n544), .A2(n491), .ZN(n520) );
  NOR2_X1 U602 ( .A1(n520), .A2(n493), .ZN(n521) );
  AND2_X1 U603 ( .A1(n522), .A2(n521), .ZN(n649) );
  INV_X1 U604 ( .A(n640), .ZN(n523) );
  NAND2_X1 U605 ( .A1(n361), .A2(n523), .ZN(n524) );
  INV_X1 U606 ( .A(KEYINPUT44), .ZN(n525) );
  NAND2_X1 U607 ( .A1(n524), .A2(n525), .ZN(n531) );
  NAND2_X1 U608 ( .A1(n640), .A2(n512), .ZN(n529) );
  INV_X1 U609 ( .A(n625), .ZN(n527) );
  NOR2_X1 U610 ( .A1(n649), .A2(n525), .ZN(n526) );
  AND2_X1 U611 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U612 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U613 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U614 ( .A1(n533), .A2(n532), .ZN(n536) );
  INV_X1 U615 ( .A(KEYINPUT84), .ZN(n534) );
  XNOR2_X1 U616 ( .A(n534), .B(KEYINPUT45), .ZN(n535) );
  XNOR2_X1 U617 ( .A(n599), .B(KEYINPUT38), .ZN(n686) );
  INV_X1 U618 ( .A(n686), .ZN(n681) );
  NAND2_X1 U619 ( .A1(n681), .A2(n684), .ZN(n538) );
  OR2_X1 U620 ( .A1(G900), .A2(n540), .ZN(n541) );
  OR2_X1 U621 ( .A1(n541), .A2(n363), .ZN(n543) );
  NAND2_X1 U622 ( .A1(n543), .A2(n542), .ZN(n561) );
  INV_X1 U623 ( .A(n561), .ZN(n549) );
  NOR2_X1 U624 ( .A1(n671), .A2(n544), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n546), .A2(n545), .ZN(n573) );
  NOR2_X1 U626 ( .A1(n699), .A2(n573), .ZN(n548) );
  XNOR2_X1 U627 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n547) );
  NOR2_X1 U628 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U629 ( .A1(n491), .A2(n684), .ZN(n552) );
  INV_X1 U630 ( .A(KEYINPUT30), .ZN(n551) );
  XNOR2_X1 U631 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n554), .A2(n553), .ZN(n586) );
  XNOR2_X1 U633 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n555) );
  XNOR2_X1 U634 ( .A(n556), .B(n555), .ZN(n602) );
  OR2_X1 U635 ( .A1(n602), .A2(n564), .ZN(n557) );
  XNOR2_X2 U636 ( .A(n557), .B(KEYINPUT40), .ZN(n623) );
  NAND2_X1 U637 ( .A1(n756), .A2(n623), .ZN(n559) );
  XNOR2_X1 U638 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n558) );
  XNOR2_X1 U639 ( .A(n559), .B(n558), .ZN(n592) );
  INV_X1 U640 ( .A(n560), .ZN(n563) );
  NAND2_X1 U641 ( .A1(n684), .A2(n561), .ZN(n562) );
  NOR2_X1 U642 ( .A1(n563), .A2(n562), .ZN(n567) );
  NOR2_X1 U643 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U644 ( .A1(n567), .A2(n566), .ZN(n595) );
  NAND2_X1 U645 ( .A1(n595), .A2(n599), .ZN(n569) );
  XOR2_X1 U646 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n568) );
  XNOR2_X1 U647 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U648 ( .A1(n570), .A2(n493), .ZN(n571) );
  XNOR2_X1 U649 ( .A(n571), .B(KEYINPUT111), .ZN(n753) );
  XNOR2_X1 U650 ( .A(n753), .B(KEYINPUT88), .ZN(n590) );
  NAND2_X1 U651 ( .A1(KEYINPUT74), .A2(n682), .ZN(n576) );
  INV_X1 U652 ( .A(n576), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n574), .A2(n651), .ZN(n575) );
  NAND2_X1 U654 ( .A1(n575), .A2(KEYINPUT47), .ZN(n580) );
  NOR2_X1 U655 ( .A1(KEYINPUT47), .A2(n576), .ZN(n578) );
  NOR2_X1 U656 ( .A1(KEYINPUT74), .A2(n682), .ZN(n577) );
  NOR2_X1 U657 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n580), .A2(n579), .ZN(n583) );
  INV_X1 U659 ( .A(n651), .ZN(n655) );
  INV_X1 U660 ( .A(KEYINPUT47), .ZN(n581) );
  NAND2_X1 U661 ( .A1(n655), .A2(n581), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n584), .A2(n599), .ZN(n585) );
  NOR2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n654) );
  INV_X1 U665 ( .A(n654), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U669 ( .A(KEYINPUT48), .ZN(n593) );
  XOR2_X1 U670 ( .A(KEYINPUT108), .B(n595), .Z(n596) );
  NOR2_X1 U671 ( .A1(n596), .A2(n493), .ZN(n598) );
  INV_X1 U672 ( .A(KEYINPUT43), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n598), .B(n597), .ZN(n601) );
  INV_X1 U674 ( .A(n599), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n624) );
  OR2_X1 U676 ( .A1(n602), .A2(n658), .ZN(n622) );
  AND2_X1 U677 ( .A1(n624), .A2(n622), .ZN(n607) );
  AND2_X1 U678 ( .A1(n607), .A2(KEYINPUT82), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n614), .A2(n604), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n605), .A2(KEYINPUT2), .ZN(n606) );
  NOR2_X1 U681 ( .A1(n606), .A2(n608), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n745), .A2(n609), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n614), .A2(n610), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n611), .A2(KEYINPUT82), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n745), .A2(KEYINPUT2), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n730), .A2(n617), .ZN(n663) );
  NOR2_X2 U688 ( .A1(n618), .A2(n663), .ZN(n707) );
  NAND2_X1 U689 ( .A1(n722), .A2(G217), .ZN(n619) );
  AND2_X1 U690 ( .A1(n712), .A2(n620), .ZN(G66) );
  XNOR2_X1 U691 ( .A(G134), .B(KEYINPUT116), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(G36) );
  XNOR2_X1 U693 ( .A(n623), .B(G131), .ZN(G33) );
  XNOR2_X1 U694 ( .A(n624), .B(G140), .ZN(G42) );
  XOR2_X1 U695 ( .A(G119), .B(n625), .Z(G21) );
  NAND2_X1 U696 ( .A1(n707), .A2(G472), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n630), .A2(n712), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n631), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U702 ( .A1(n707), .A2(G475), .ZN(n636) );
  XOR2_X1 U703 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT59), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U707 ( .A1(n637), .A2(n712), .ZN(n639) );
  XNOR2_X1 U708 ( .A(KEYINPUT65), .B(KEYINPUT60), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(G60) );
  XOR2_X1 U710 ( .A(n640), .B(G122), .Z(G24) );
  XOR2_X1 U711 ( .A(G101), .B(n641), .Z(G3) );
  NOR2_X1 U712 ( .A1(n564), .A2(n643), .ZN(n642) );
  XOR2_X1 U713 ( .A(G104), .B(n642), .Z(G6) );
  NOR2_X1 U714 ( .A1(n658), .A2(n643), .ZN(n648) );
  XOR2_X1 U715 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n645) );
  XNOR2_X1 U716 ( .A(G107), .B(KEYINPUT26), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(n646), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(G9) );
  XOR2_X1 U720 ( .A(G110), .B(n649), .Z(G12) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n653) );
  INV_X1 U722 ( .A(n658), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(G30) );
  XOR2_X1 U725 ( .A(G143), .B(n654), .Z(G45) );
  NOR2_X1 U726 ( .A1(n655), .A2(n564), .ZN(n656) );
  XOR2_X1 U727 ( .A(G146), .B(n656), .Z(G48) );
  NOR2_X1 U728 ( .A1(n659), .A2(n564), .ZN(n657) );
  XOR2_X1 U729 ( .A(G113), .B(n657), .Z(G15) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U731 ( .A(G116), .B(n660), .Z(G18) );
  INV_X1 U732 ( .A(n745), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n730), .A2(n661), .ZN(n662) );
  NOR2_X1 U734 ( .A1(n662), .A2(KEYINPUT2), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  INV_X1 U736 ( .A(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT50), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n672), .B(KEYINPUT117), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT49), .B(n673), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n676), .A2(n491), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U745 ( .A(KEYINPUT51), .B(n679), .Z(n680) );
  NOR2_X1 U746 ( .A1(n699), .A2(n680), .ZN(n693) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n683), .A2(n687), .ZN(n685) );
  AND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U752 ( .A(n690), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n691), .A2(n698), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U755 ( .A(n694), .B(KEYINPUT52), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(n697), .B(KEYINPUT118), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U760 ( .A(KEYINPUT119), .B(n702), .Z(n703) );
  NAND2_X1 U761 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U762 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n706), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U764 ( .A1(n707), .A2(G210), .ZN(n711) );
  XOR2_X1 U765 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n708) );
  XOR2_X1 U766 ( .A(n709), .B(n708), .Z(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n713) );
  INV_X1 U768 ( .A(n712), .ZN(n726) );
  XNOR2_X1 U769 ( .A(n714), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U770 ( .A1(n722), .A2(G469), .ZN(n720) );
  XOR2_X1 U771 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n716) );
  XNOR2_X1 U772 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n715) );
  XNOR2_X1 U773 ( .A(n716), .B(n715), .ZN(n718) );
  XOR2_X1 U774 ( .A(n718), .B(n717), .Z(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U776 ( .A1(n726), .A2(n721), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n722), .A2(G478), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(G63) );
  XNOR2_X1 U780 ( .A(n727), .B(G101), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n738) );
  NOR2_X1 U782 ( .A1(n730), .A2(G953), .ZN(n736) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n731) );
  XOR2_X1 U784 ( .A(KEYINPUT61), .B(n731), .Z(n732) );
  NOR2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n734), .B(KEYINPUT124), .ZN(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n739), .B(KEYINPUT4), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n741), .B(n740), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n743), .B(n742), .ZN(n748) );
  XNOR2_X1 U792 ( .A(n748), .B(KEYINPUT125), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(n363), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n747), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U796 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U798 ( .A1(G953), .A2(n750), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U800 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n755) );
  XNOR2_X1 U801 ( .A(G125), .B(n753), .ZN(n754) );
  XNOR2_X1 U802 ( .A(n755), .B(n754), .ZN(G27) );
  XNOR2_X1 U803 ( .A(n756), .B(G137), .ZN(G39) );
endmodule

