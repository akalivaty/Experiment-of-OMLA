//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  XOR2_X1   g006(.A(G127gat), .B(G134gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n210), .B(new_n213), .C1(new_n214), .C2(KEYINPUT2), .ZN(new_n215));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n210), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT69), .B(G113gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n206), .B(new_n220), .C1(new_n221), .C2(new_n205), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n209), .A2(new_n215), .A3(new_n219), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n209), .A2(new_n222), .B1(new_n219), .B2(new_n215), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n203), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n215), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n219), .A2(new_n215), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n222), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n209), .A2(new_n222), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n219), .A2(new_n215), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT4), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n223), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n233), .A2(new_n202), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n223), .B(KEYINPUT4), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n241), .A2(KEYINPUT5), .A3(new_n202), .A4(new_n233), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G1gat), .B(G29gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT0), .ZN(new_n245));
  XNOR2_X1  g044(.A(G57gat), .B(G85gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249));
  INV_X1    g048(.A(new_n247), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n240), .A2(new_n242), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n251), .A2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G78gat), .B(G106gat), .Z(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT31), .B(G50gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G22gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G228gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT76), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n260), .A2(new_n261), .B1(G211gat), .B2(G218gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G197gat), .B(G204gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n267), .A3(new_n265), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(KEYINPUT82), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n264), .A2(new_n272), .A3(new_n267), .A4(new_n265), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n235), .B1(new_n276), .B2(new_n230), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT77), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n264), .A2(new_n267), .A3(new_n265), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n267), .B1(new_n264), .B2(new_n265), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n269), .A2(KEYINPUT77), .A3(new_n270), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n281), .A2(new_n282), .B1(new_n274), .B2(new_n231), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n259), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n231), .A2(new_n274), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT29), .B1(new_n269), .B2(new_n270), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n228), .B1(new_n288), .B2(KEYINPUT3), .ZN(new_n289));
  INV_X1    g088(.A(new_n259), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n258), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n257), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n279), .A2(new_n280), .A3(new_n272), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n274), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n230), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n228), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n290), .B1(new_n298), .B2(new_n287), .ZN(new_n299));
  INV_X1    g098(.A(new_n291), .ZN(new_n300));
  OAI21_X1  g099(.A(G22gat), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n258), .A3(new_n291), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT35), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n301), .A2(new_n293), .A3(new_n302), .A4(new_n257), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n254), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT68), .ZN(new_n310));
  INV_X1    g109(.A(G169gat), .ZN(new_n311));
  INV_X1    g110(.A(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(KEYINPUT26), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT68), .B1(new_n308), .B2(new_n309), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G183gat), .ZN(new_n320));
  INV_X1    g119(.A(G190gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(KEYINPUT28), .ZN(new_n323));
  AND2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(new_n322), .B2(KEYINPUT28), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n316), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n327), .B(new_n328), .C1(G169gat), .C2(G176gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT66), .B1(new_n309), .B2(KEYINPUT23), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  AND4_X1   g131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n321), .A3(KEYINPUT65), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(G183gat), .B2(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT64), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT64), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n324), .A2(KEYINPUT24), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n337), .A2(new_n341), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT25), .B1(new_n333), .B2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n329), .A3(new_n331), .A4(new_n332), .ZN(new_n347));
  OR2_X1    g146(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n317), .A2(new_n321), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n338), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  NOR2_X1   g150(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n351), .B1(new_n324), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n326), .B1(new_n346), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G226gat), .ZN(new_n357));
  INV_X1    g156(.A(G233gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT29), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n359), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n326), .B(new_n363), .C1(new_n346), .C2(new_n355), .ZN(new_n364));
  INV_X1    g163(.A(new_n285), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n362), .A2(KEYINPUT79), .A3(new_n364), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n365), .B1(new_n362), .B2(new_n364), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT80), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n370), .A2(new_n372), .A3(new_n380), .A4(new_n373), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n382));
  OR3_X1    g181(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n327), .B1(new_n313), .B2(new_n328), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n331), .A2(new_n332), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n345), .A2(new_n386), .A3(new_n329), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n355), .B1(new_n387), .B2(new_n351), .ZN(new_n388));
  INV_X1    g187(.A(new_n326), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n234), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n326), .B(new_n232), .C1(new_n346), .C2(new_n355), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT70), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT70), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  XNOR2_X1  g198(.A(G15gat), .B(G43gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n394), .B2(KEYINPUT32), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n402), .A2(KEYINPUT71), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(KEYINPUT71), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT33), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n394), .A2(KEYINPUT32), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n392), .B1(new_n390), .B2(new_n393), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT34), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n390), .A2(new_n393), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n414), .A3(new_n391), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT74), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n410), .A2(new_n420), .A3(new_n414), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n416), .A3(new_n422), .A4(new_n408), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT75), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT75), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  AOI221_X4 g227(.A(new_n307), .B1(new_n382), .B2(new_n383), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n404), .A2(KEYINPUT72), .A3(new_n408), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT72), .B1(new_n404), .B2(new_n408), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n412), .A2(new_n415), .B1(new_n419), .B2(new_n421), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n425), .A2(new_n306), .A3(new_n304), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT86), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n248), .A2(new_n249), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n248), .A2(new_n438), .A3(new_n249), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n251), .A3(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n383), .A2(new_n382), .B1(new_n440), .B2(new_n253), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n409), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n404), .A2(KEYINPUT72), .A3(new_n408), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n423), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n304), .A2(new_n306), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n425), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n435), .A2(new_n441), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n429), .B1(new_n449), .B2(KEYINPUT35), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n426), .A2(new_n451), .A3(new_n428), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(KEYINPUT36), .A3(new_n425), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n382), .A2(new_n383), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n253), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n304), .A2(KEYINPUT84), .A3(new_n306), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT84), .B1(new_n304), .B2(new_n306), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n233), .A2(new_n238), .A3(new_n236), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n203), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n202), .B1(new_n241), .B2(new_n233), .ZN(new_n465));
  INV_X1    g264(.A(new_n225), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n202), .A3(new_n223), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT39), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n247), .B(new_n464), .C1(new_n465), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n251), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n470), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n382), .A2(new_n383), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT37), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n370), .A2(new_n372), .A3(new_n478), .A4(new_n373), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n479), .A2(new_n378), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n374), .B2(KEYINPUT37), .ZN(new_n482));
  INV_X1    g281(.A(new_n366), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n483), .B2(new_n371), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n378), .A3(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n480), .A2(new_n482), .B1(new_n485), .B2(new_n481), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n381), .A2(new_n252), .A3(new_n253), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n477), .B(new_n447), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n454), .A2(new_n461), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n450), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(G1gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493));
  AOI21_X1  g292(.A(G8gat), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n494), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G43gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G50gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(G50gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR3_X1    g306(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT91), .B(G36gat), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n511), .A2(G29gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n504), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(KEYINPUT92), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n502), .A2(KEYINPUT93), .ZN(new_n515));
  INV_X1    g314(.A(G50gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT93), .A3(G43gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n500), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n503), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT15), .B1(new_n499), .B2(G50gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n501), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n511), .A2(G29gat), .B1(new_n508), .B2(new_n505), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n514), .A2(new_n519), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n525), .A2(KEYINPUT17), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(KEYINPUT17), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n498), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n525), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n498), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT95), .B1(new_n498), .B2(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n532), .B(KEYINPUT13), .Z(new_n538));
  INV_X1    g337(.A(new_n498), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT95), .A3(new_n525), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT18), .A4(new_n532), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT88), .ZN(new_n545));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT89), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n545), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n548), .A2(new_n550), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT12), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n551), .B2(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n542), .A2(KEYINPUT96), .A3(new_n543), .A4(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n535), .A2(new_n541), .A3(new_n557), .A4(new_n543), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n543), .ZN(new_n562));
  INV_X1    g361(.A(new_n557), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n558), .A2(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n565), .A2(KEYINPUT97), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n539), .B1(KEYINPUT21), .B2(new_n569), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT98), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n574), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G190gat), .B(G218gat), .Z(new_n583));
  NOR2_X1   g382(.A1(new_n526), .A2(new_n527), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT102), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT7), .ZN(new_n587));
  AND2_X1   g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT101), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n585), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n591), .A2(new_n587), .A3(new_n588), .A4(KEYINPUT102), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n593), .B(new_n594), .C1(new_n590), .C2(new_n588), .ZN(new_n595));
  XNOR2_X1  g394(.A(G99gat), .B(G106gat), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT103), .B(G85gat), .Z(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n597), .A2(new_n598), .B1(KEYINPUT8), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n596), .B1(new_n595), .B2(new_n600), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n584), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n525), .ZN(new_n606));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT99), .Z(new_n608));
  INV_X1    g407(.A(KEYINPUT41), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n583), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n605), .A2(new_n611), .A3(new_n583), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n609), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT100), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OAI22_X1  g417(.A1(new_n613), .A2(new_n614), .B1(KEYINPUT104), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n614), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n612), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(KEYINPUT104), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n619), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n582), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n567), .B(new_n568), .Z(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n602), .B2(new_n603), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  INV_X1    g427(.A(new_n593), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n594), .B1(new_n590), .B2(new_n588), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n600), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n596), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n569), .A2(new_n633), .A3(new_n601), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT107), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n627), .A2(new_n634), .ZN(new_n641));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT107), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n644), .B(new_n642), .C1(new_n635), .C2(new_n636), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT106), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n635), .A2(KEYINPUT105), .A3(new_n636), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT105), .B1(new_n635), .B2(new_n636), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n653), .A2(new_n654), .A3(new_n642), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n643), .A3(new_n650), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n625), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n490), .A2(new_n564), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n456), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(new_n455), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT16), .B(G8gat), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT109), .Z(new_n670));
  XOR2_X1   g469(.A(new_n666), .B(KEYINPUT108), .Z(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n671), .B2(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(G8gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(G15gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n426), .A2(new_n428), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n454), .B(KEYINPUT110), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n677), .B1(new_n680), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n661), .A2(new_n460), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  OAI21_X1  g483(.A(new_n624), .B1(new_n450), .B2(new_n489), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n691));
  INV_X1    g490(.A(new_n429), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n454), .A2(new_n461), .A3(new_n488), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n450), .A2(new_n489), .A3(KEYINPUT112), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n624), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n688), .A2(new_n689), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n564), .A2(new_n658), .A3(new_n581), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT113), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n696), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT112), .B1(new_n450), .B2(new_n489), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n699), .ZN(new_n706));
  INV_X1    g505(.A(new_n689), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT111), .B1(new_n685), .B2(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n701), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n456), .ZN(new_n713));
  INV_X1    g512(.A(new_n685), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n701), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n456), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT45), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n717), .ZN(G1328gat));
  OAI21_X1  g517(.A(new_n511), .B1(new_n712), .B2(new_n455), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n715), .A2(new_n455), .A3(new_n511), .ZN(new_n723));
  MUX2_X1   g522(.A(new_n722), .B(new_n720), .S(new_n723), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n724), .ZN(G1329gat));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n701), .ZN(new_n726));
  OAI21_X1  g525(.A(G43gat), .B1(new_n726), .B2(new_n454), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n714), .A2(new_n499), .A3(new_n676), .A4(new_n701), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(KEYINPUT47), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n728), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n703), .A2(new_n678), .A3(new_n711), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(G43gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n732), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g532(.A(KEYINPUT48), .B(G50gat), .C1(new_n726), .C2(new_n447), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n516), .A3(new_n460), .A4(new_n701), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(KEYINPUT48), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n703), .A2(new_n460), .A3(new_n711), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G50gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g540(.A1(new_n625), .A2(new_n564), .A3(new_n658), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n695), .A2(new_n696), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n662), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n665), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT49), .B(G64gat), .Z(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n746), .B2(new_n748), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n743), .A2(new_n750), .A3(new_n676), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n743), .A2(new_n678), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n750), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n743), .A2(new_n460), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  INV_X1    g556(.A(new_n564), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n581), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n624), .B(new_n759), .C1(new_n450), .C2(new_n489), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n658), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n662), .A3(new_n597), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n759), .A2(new_n658), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n700), .A2(new_n456), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n597), .ZN(G1336gat));
  NOR2_X1   g567(.A1(new_n700), .A2(new_n766), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n598), .B1(new_n769), .B2(new_n665), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(KEYINPUT51), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n760), .B(new_n772), .ZN(new_n773));
  AND4_X1   g572(.A1(new_n598), .A2(new_n773), .A3(new_n665), .A4(new_n658), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n665), .A2(new_n598), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n763), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n770), .B2(new_n778), .ZN(G1337gat));
  XNOR2_X1  g578(.A(KEYINPUT118), .B(G99gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n676), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n769), .A2(new_n678), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(new_n780), .ZN(G1338gat));
  NOR2_X1   g582(.A1(new_n447), .A2(G106gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n773), .A2(new_n658), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT119), .ZN(new_n786));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n769), .B2(new_n460), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT53), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n764), .B2(new_n784), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n700), .A2(new_n447), .A3(new_n766), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n787), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT54), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT55), .B1(new_n655), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n639), .B2(new_n645), .ZN(new_n798));
  INV_X1    g597(.A(new_n650), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT121), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(KEYINPUT121), .A3(new_n799), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n657), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT122), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n795), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n656), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n798), .A2(KEYINPUT121), .A3(new_n799), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT121), .B1(new_n798), .B2(new_n799), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n564), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n796), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n809), .B2(new_n810), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n657), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n806), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n558), .A2(new_n561), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n538), .B1(new_n540), .B2(new_n537), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n532), .B1(new_n528), .B2(new_n531), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n553), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n658), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n624), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n811), .A2(new_n812), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(new_n624), .A3(new_n822), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AND4_X1   g626(.A1(new_n806), .A2(new_n817), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n582), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n625), .A2(new_n659), .A3(new_n564), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT120), .Z(new_n831));
  AOI21_X1  g630(.A(new_n456), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n435), .A2(new_n448), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n665), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n221), .A3(new_n758), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n460), .B1(new_n829), .B2(new_n831), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(new_n662), .A3(new_n676), .A4(new_n455), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n564), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(G1340gat));
  AOI21_X1  g640(.A(G120gat), .B1(new_n836), .B2(new_n658), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n839), .A2(new_n205), .A3(new_n659), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n839), .B2(new_n582), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n582), .A2(G127gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n835), .B2(new_n846), .ZN(G1342gat));
  NOR3_X1   g646(.A1(new_n835), .A2(G134gat), .A3(new_n698), .ZN(new_n848));
  XOR2_X1   g647(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n849));
  OR2_X1    g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n839), .B2(new_n698), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  AOI211_X1 g652(.A(new_n456), .B(new_n665), .C1(new_n452), .C2(new_n453), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n829), .A2(new_n831), .ZN(new_n855));
  INV_X1    g654(.A(new_n447), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n460), .A2(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n813), .A2(new_n657), .A3(new_n815), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n624), .B1(new_n859), .B2(new_n823), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n582), .B1(new_n860), .B2(new_n828), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n858), .B1(new_n861), .B2(new_n831), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n758), .B(new_n854), .C1(new_n857), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G141gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n678), .A2(new_n447), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n455), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n564), .A2(G141gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n832), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT58), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n864), .A2(new_n869), .A3(new_n873), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1344gat));
  AND2_X1   g676(.A1(new_n832), .A2(new_n867), .ZN(new_n878));
  INV_X1    g677(.A(G148gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n879), .A3(new_n658), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n854), .B1(new_n857), .B2(new_n862), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n659), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G148gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n447), .B1(new_n829), .B2(new_n831), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n861), .A2(new_n830), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n887), .A3(new_n460), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n888), .A2(new_n658), .A3(new_n854), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n883), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n880), .B1(new_n885), .B2(new_n892), .ZN(G1345gat));
  OAI21_X1  g692(.A(G155gat), .B1(new_n881), .B2(new_n582), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n211), .A3(new_n581), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n881), .B2(new_n698), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n212), .A3(new_n624), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  NAND4_X1  g698(.A1(new_n838), .A2(new_n456), .A3(new_n676), .A4(new_n665), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n311), .A3(new_n564), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n855), .B2(new_n456), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT125), .B(new_n662), .C1(new_n829), .C2(new_n831), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n833), .A2(new_n455), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n758), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n907), .B2(new_n311), .ZN(G1348gat));
  OAI21_X1  g707(.A(G176gat), .B1(new_n900), .B2(new_n659), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n658), .A2(new_n312), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1349gat));
  OAI21_X1  g711(.A(G183gat), .B1(new_n900), .B2(new_n582), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n581), .A2(new_n318), .A3(new_n320), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n906), .B(new_n914), .C1(new_n903), .C2(new_n904), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n900), .B2(new_n698), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT61), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n698), .A2(G190gat), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n906), .B(new_n920), .C1(new_n903), .C2(new_n904), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(G1351gat));
  NOR3_X1   g722(.A1(new_n678), .A2(new_n662), .A3(new_n455), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n890), .B(new_n924), .C1(new_n886), .C2(new_n887), .ZN(new_n925));
  INV_X1    g724(.A(G197gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n925), .A2(new_n926), .A3(new_n564), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n865), .A2(new_n665), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n905), .A2(new_n758), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n926), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n659), .A2(G204gat), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n929), .B(new_n932), .C1(new_n903), .C2(new_n904), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n934));
  OAI21_X1  g733(.A(G204gat), .B1(new_n925), .B2(new_n659), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G1353gat));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(KEYINPUT127), .ZN(new_n939));
  INV_X1    g738(.A(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(KEYINPUT127), .B2(new_n938), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n939), .B(new_n941), .C1(new_n925), .C2(new_n582), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n888), .A2(new_n581), .A3(new_n890), .A4(new_n924), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n939), .B1(new_n944), .B2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n905), .A2(new_n929), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n581), .A2(new_n940), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n943), .A2(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n925), .B2(new_n698), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n698), .A2(G218gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n946), .B2(new_n950), .ZN(G1355gat));
endmodule


