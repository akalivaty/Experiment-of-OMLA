//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0003(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n204), .B1(new_n205), .B2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G13), .ZN(new_n207));
  NAND4_X1  g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G50), .A2(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT67), .Z(new_n233));
  AOI211_X1 g0033(.A(new_n211), .B(new_n227), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT69), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n257), .A2(new_n258), .B1(new_n219), .B2(new_n252), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n251), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(G274), .C1(G41), .C2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND3_X1  g0066(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G226), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n260), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT76), .B(G200), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT74), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n275), .A2(new_n261), .A3(G13), .A4(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n228), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n279), .A3(new_n228), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n261), .A2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G50), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT73), .B1(new_n288), .B2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT73), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(new_n229), .A3(G33), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(KEYINPUT8), .A2(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT8), .A2(G58), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g0099(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n297), .A2(new_n299), .B1(new_n300), .B2(new_n229), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n284), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n287), .B(new_n302), .C1(G50), .C2(new_n277), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n271), .A2(new_n272), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n271), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G190), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n307), .C1(new_n304), .C2(new_n303), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n303), .C1(G169), .C2(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n268), .A2(G238), .A3(new_n269), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G226), .A2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n223), .B2(G1698), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n252), .B1(G33), .B2(G97), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n266), .A2(new_n263), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n315), .B(new_n262), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n223), .A2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G226), .B2(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n322), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n251), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n315), .A4(new_n262), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n314), .B1(new_n333), .B2(G169), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n310), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n314), .A3(G169), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT77), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n277), .B2(G68), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n340), .B(KEYINPUT12), .C1(new_n277), .C2(G68), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n214), .B1(new_n261), .B2(G20), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n343), .A2(new_n344), .B1(new_n285), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G50), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n299), .A2(new_n347), .B1(new_n229), .B2(G68), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n289), .A2(new_n291), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(G77), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n280), .A2(new_n279), .A3(new_n228), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n281), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT11), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT11), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n292), .A2(new_n219), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n354), .B(new_n284), .C1(new_n355), .C2(new_n348), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n346), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n339), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G190), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n258), .A2(new_n253), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n252), .B(new_n362), .C1(G226), .C2(new_n253), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n251), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n367), .A2(KEYINPUT82), .A3(new_n262), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT82), .B1(new_n367), .B2(new_n262), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n361), .B(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n319), .B1(new_n363), .B2(new_n364), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n262), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT80), .B1(new_n326), .B2(G33), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n288), .A3(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n379), .A3(new_n327), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n252), .B2(G20), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n214), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n222), .A2(new_n214), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n298), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n376), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n252), .A2(new_n382), .A3(G20), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n328), .B2(new_n229), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n389), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n390), .A2(new_n284), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n293), .A2(new_n286), .A3(new_n294), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n352), .A2(new_n277), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n278), .A2(new_n295), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT81), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT81), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n375), .A2(new_n396), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n383), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n389), .B1(new_n409), .B2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n352), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n390), .B1(new_n401), .B2(new_n403), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n310), .B(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n372), .B2(new_n373), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT18), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n396), .A2(new_n404), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n413), .A2(new_n415), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n375), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n407), .A2(new_n417), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n285), .A2(G77), .A3(new_n286), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT75), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n295), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT15), .B(G87), .Z(new_n428));
  AOI22_X1  g0228(.A1(new_n298), .A2(new_n427), .B1(new_n428), .B2(new_n349), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n229), .B2(new_n219), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n284), .B1(new_n219), .B2(new_n278), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n257), .A2(new_n215), .B1(new_n432), .B2(new_n252), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n328), .A2(new_n223), .A3(G1698), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n251), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n268), .A2(new_n269), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n262), .C1(new_n220), .C2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n426), .B(new_n431), .C1(new_n361), .C2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n272), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OR3_X1    g0240(.A1(new_n360), .A2(new_n423), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT78), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n321), .A2(G190), .A3(new_n332), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n357), .A3(new_n346), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n371), .B1(new_n321), .B2(new_n332), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n358), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n333), .A2(G200), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT78), .A4(new_n443), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n426), .A2(new_n431), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n437), .A2(new_n414), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n437), .A2(G179), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n313), .A2(new_n441), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT88), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n268), .A2(G274), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT85), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G41), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n464), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n251), .B1(new_n252), .B2(G303), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n253), .A2(G257), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G264), .A2(G1698), .ZN(new_n475));
  AND4_X1   g0275(.A1(new_n325), .A2(new_n327), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n472), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G303), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n319), .B1(new_n328), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n252), .A2(new_n475), .A3(new_n474), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n471), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n470), .A2(new_n268), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G270), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n371), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n278), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n261), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n352), .A2(G116), .A3(new_n277), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n229), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT83), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n492), .B1(new_n497), .B2(G33), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n280), .A2(new_n228), .B1(G20), .B2(new_n486), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT20), .B1(new_n498), .B2(new_n499), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n487), .B(new_n489), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n460), .B1(new_n485), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n477), .A2(new_n481), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n461), .A2(new_n470), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n484), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G200), .ZN(new_n507));
  INV_X1    g0307(.A(new_n502), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(KEYINPUT88), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n482), .A2(G190), .A3(new_n484), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n502), .A3(G169), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(new_n502), .A3(G169), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n504), .A2(G179), .A3(new_n505), .A4(new_n484), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n515), .A2(new_n512), .B1(new_n517), .B2(new_n502), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n381), .A2(new_n383), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(G107), .B1(G77), .B2(new_n298), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT83), .B(G97), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n523));
  XOR2_X1   g0323(.A(G97), .B(G107), .Z(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(KEYINPUT6), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G20), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n352), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n277), .A2(new_n282), .A3(new_n283), .A4(new_n488), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n352), .A2(KEYINPUT84), .A3(new_n277), .A4(new_n488), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(G97), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n278), .A2(new_n493), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n490), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n325), .A2(new_n327), .A3(G244), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n252), .A2(G250), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n253), .B1(new_n542), .B2(KEYINPUT4), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n251), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n470), .A2(G257), .A3(new_n268), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n544), .A2(new_n361), .A3(new_n505), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(new_n252), .B2(G250), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n539), .B(new_n540), .C1(new_n253), .C2(new_n548), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n471), .B(new_n545), .C1(new_n549), .C2(new_n251), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(G200), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n535), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n253), .A2(G257), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n252), .B(new_n553), .C1(G250), .C2(G1698), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G294), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n319), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n471), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n483), .A2(G264), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n361), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n251), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n561), .A2(new_n558), .A3(new_n505), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(G200), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n277), .A2(G107), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n564), .B(KEYINPUT25), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n530), .A2(G107), .A3(new_n531), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n325), .A2(new_n327), .A3(new_n229), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n252), .A2(new_n569), .A3(new_n229), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n288), .A2(new_n486), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n229), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n229), .A2(G107), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT23), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n571), .A2(KEYINPUT24), .A3(new_n573), .A4(new_n575), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n284), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n563), .A2(new_n565), .A3(new_n566), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n544), .A2(new_n505), .A3(new_n546), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n414), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n544), .A2(new_n310), .A3(new_n505), .A4(new_n546), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n527), .C2(new_n534), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n552), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n580), .A2(new_n565), .A3(new_n566), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n310), .A2(new_n561), .A3(new_n558), .A4(new_n505), .ZN(new_n588));
  AOI21_X1  g0388(.A(G169), .B1(new_n557), .B2(new_n558), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n277), .A2(new_n428), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n292), .B2(new_n497), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n229), .B1(new_n322), .B2(new_n593), .ZN(new_n595));
  INV_X1    g0395(.A(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n432), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n522), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n252), .A2(new_n229), .A3(G68), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n592), .B1(new_n600), .B2(new_n284), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n530), .A2(G87), .A3(new_n531), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n268), .A2(G274), .A3(new_n468), .ZN(new_n604));
  INV_X1    g0404(.A(new_n468), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n268), .A2(G250), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G238), .A2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n220), .B2(G1698), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n572), .B1(new_n608), .B2(new_n252), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n604), .B(new_n606), .C1(new_n609), .C2(new_n319), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(new_n361), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n272), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n603), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n530), .A2(new_n428), .A3(new_n531), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n601), .A2(new_n615), .B1(new_n414), .B2(new_n610), .ZN(new_n616));
  INV_X1    g0416(.A(new_n610), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n310), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n591), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n519), .A2(new_n586), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n459), .A2(new_n621), .ZN(G372));
  AND2_X1   g0422(.A1(new_n552), .A2(new_n585), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n601), .A2(new_n613), .A3(new_n602), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT89), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n611), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n601), .A2(KEYINPUT89), .A3(new_n602), .A4(new_n613), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n618), .B2(new_n616), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n591), .A2(new_n518), .A3(new_n514), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n623), .A2(new_n581), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n585), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n619), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n550), .A2(G169), .ZN(new_n635));
  INV_X1    g0435(.A(new_n584), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n527), .A2(new_n534), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n614), .A3(new_n619), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n630), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n459), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n312), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n457), .B1(new_n446), .B2(new_n449), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n407), .B(new_n422), .C1(new_n644), .C2(new_n360), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n417), .A2(new_n421), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n643), .B1(new_n647), .B2(new_n309), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n648), .ZN(G369));
  AND3_X1   g0449(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n261), .A2(new_n229), .A3(G13), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT90), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(new_n655), .A3(G213), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n508), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n518), .A2(new_n514), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  INV_X1    g0463(.A(new_n657), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n591), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n587), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n581), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n591), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n661), .A2(new_n664), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n209), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n522), .A2(G116), .A3(new_n597), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n232), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT92), .ZN(new_n679));
  XNOR2_X1  g0479(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n641), .A2(new_n657), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT29), .ZN(new_n683));
  INV_X1    g0483(.A(new_n628), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT26), .B1(new_n684), .B2(new_n585), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n630), .A3(new_n686), .A4(new_n619), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n657), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n617), .A2(new_n544), .A3(new_n546), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n557), .A2(new_n558), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n516), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT30), .B1(new_n693), .B2(KEYINPUT93), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n617), .A2(new_n544), .A3(new_n546), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n517), .A3(new_n562), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n582), .A2(new_n506), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n310), .A3(new_n610), .A4(new_n692), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n664), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n620), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n552), .A2(new_n581), .A3(new_n585), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n650), .A2(new_n706), .A3(new_n707), .A4(new_n657), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n690), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n681), .B1(new_n713), .B2(G1), .ZN(G364));
  NOR2_X1   g0514(.A1(new_n207), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n261), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n674), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n663), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G330), .B2(new_n662), .ZN(new_n720));
  INV_X1    g0520(.A(new_n718), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n228), .B1(G20), .B2(new_n414), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n310), .A2(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n229), .A2(G190), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G179), .A2(G200), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n229), .B1(new_n728), .B2(G190), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(G311), .A2(new_n727), .B1(new_n730), .B2(G294), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n229), .A2(new_n310), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n361), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(G317), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(KEYINPUT33), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(KEYINPUT33), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n229), .A2(new_n361), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n272), .A2(new_n310), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n725), .A2(new_n728), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n739), .A2(G303), .B1(G329), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n732), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n361), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n252), .B1(new_n744), .B2(G326), .ZN(new_n745));
  AND4_X1   g0545(.A1(new_n731), .A2(new_n736), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n272), .A2(new_n310), .A3(new_n725), .ZN(new_n748));
  INV_X1    g0548(.A(G322), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n737), .A2(new_n724), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n746), .B1(new_n747), .B2(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n252), .B1(new_n750), .B2(new_n222), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n748), .A2(new_n432), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(G50), .C2(new_n744), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n727), .A2(G77), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n733), .A2(new_n214), .B1(new_n729), .B2(new_n493), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(G87), .B2(new_n739), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n754), .A2(new_n755), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n723), .B1(new_n751), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n722), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n233), .A2(new_n467), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n673), .A2(new_n252), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n246), .C2(new_n467), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n209), .A2(G355), .A3(new_n252), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(G116), .C2(new_n209), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n721), .B(new_n762), .C1(new_n766), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n765), .B(KEYINPUT94), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n662), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n720), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  NAND2_X1  g0577(.A1(new_n454), .A2(new_n664), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n438), .B2(new_n439), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n457), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n457), .A2(new_n664), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n682), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT98), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n457), .B2(new_n779), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n641), .A2(new_n657), .A3(new_n786), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n784), .B1(new_n785), .B2(new_n787), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(new_n712), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n721), .ZN(new_n792));
  INV_X1    g0592(.A(new_n733), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G150), .ZN(new_n794));
  INV_X1    g0594(.A(new_n750), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G143), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  INV_X1    g0598(.A(new_n744), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n799), .C1(new_n756), .C2(new_n726), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n252), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n800), .ZN(new_n803));
  INV_X1    g0603(.A(new_n801), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(new_n222), .B2(new_n729), .ZN(new_n805));
  INV_X1    g0605(.A(new_n748), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n802), .B(new_n805), .C1(G68), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n347), .B2(new_n738), .C1(new_n808), .C2(new_n740), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n748), .A2(new_n596), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT95), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n733), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n811), .B1(new_n816), .B2(new_n747), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n328), .B1(new_n738), .B2(new_n432), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT96), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n740), .A2(new_n820), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n726), .A2(new_n486), .B1(new_n729), .B2(new_n493), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n817), .A2(new_n819), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n750), .C1(new_n478), .C2(new_n799), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n723), .B1(new_n809), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n722), .A2(new_n763), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n721), .B(new_n826), .C1(new_n219), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n764), .B2(new_n786), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n792), .A2(new_n829), .ZN(G384));
  AOI211_X1 g0630(.A(KEYINPUT14), .B(new_n414), .C1(new_n321), .C2(new_n332), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n334), .A2(new_n831), .A3(new_n336), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n452), .A2(new_n453), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n447), .A2(new_n657), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n446), .B2(new_n449), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n832), .A2(new_n837), .A3(new_n447), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT99), .B1(new_n339), .B2(new_n358), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n783), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT40), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n703), .B2(new_n704), .ZN(new_n844));
  AOI211_X1 g0644(.A(KEYINPUT103), .B(KEYINPUT31), .C1(new_n702), .C2(new_n664), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT104), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n709), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n702), .A2(KEYINPUT104), .A3(KEYINPUT31), .A4(new_n664), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n708), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n841), .B(new_n842), .C1(new_n846), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n214), .B1(new_n383), .B2(new_n408), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n376), .B1(new_n854), .B2(new_n389), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n395), .A2(new_n855), .A3(new_n284), .ZN(new_n856));
  INV_X1    g0656(.A(new_n400), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n856), .A2(KEYINPUT100), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT100), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n423), .A2(new_n656), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n857), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n656), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n416), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n856), .A2(KEYINPUT100), .A3(new_n857), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n862), .B1(new_n869), .B2(new_n405), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n656), .B1(new_n413), .B2(new_n415), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n405), .B(new_n862), .C1(new_n412), .C2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n853), .B1(new_n861), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n858), .A2(new_n859), .A3(new_n871), .ZN(new_n876));
  INV_X1    g0676(.A(new_n405), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n872), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n423), .A2(new_n656), .A3(new_n860), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n423), .A2(new_n418), .A3(new_n656), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n405), .B1(new_n412), .B2(new_n871), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n872), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n853), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n881), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n841), .C1(new_n846), .C2(new_n850), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n852), .A2(new_n882), .B1(KEYINPUT40), .B2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n621), .A2(new_n657), .B1(new_n709), .B2(new_n847), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n849), .C1(new_n844), .C2(new_n845), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n459), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n891), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G330), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n690), .A2(new_n459), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n648), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n837), .B1(new_n832), .B2(new_n447), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n339), .A2(KEYINPUT99), .A3(new_n358), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n833), .A2(new_n834), .B1(new_n904), .B2(new_n836), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n787), .B2(new_n782), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n882), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n904), .A2(new_n664), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n646), .A2(new_n656), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n901), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n261), .B2(new_n715), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n486), .B1(new_n525), .B2(KEYINPUT35), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n231), .C1(KEYINPUT35), .C2(new_n525), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n222), .B2(new_n214), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n232), .B1(G50), .B2(new_n214), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n207), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n922), .A3(new_n925), .ZN(G367));
  OAI21_X1  g0726(.A(new_n623), .B1(new_n535), .B2(new_n657), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n632), .A2(new_n664), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n668), .A3(new_n670), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n930), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n585), .B1(new_n927), .B2(new_n591), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n930), .A2(KEYINPUT42), .B1(new_n657), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT105), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n628), .B1(new_n603), .B2(new_n657), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n619), .A2(new_n603), .A3(new_n657), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n935), .A2(new_n943), .A3(new_n939), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n929), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n945), .A2(new_n669), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT106), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n945), .B1(new_n669), .B2(new_n946), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n674), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n668), .A2(new_n670), .ZN(new_n952));
  INV_X1    g0752(.A(new_n665), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n946), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT44), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n954), .B2(new_n946), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n671), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n957), .A2(new_n669), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n961), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n663), .B(new_n668), .C1(new_n956), .C2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT107), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n668), .B(new_n670), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n663), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n713), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n962), .A2(new_n964), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT107), .B1(new_n972), .B2(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n951), .B1(new_n974), .B2(new_n713), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n948), .B(new_n949), .C1(new_n975), .C2(new_n717), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n726), .A2(new_n347), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n252), .B1(new_n214), .B2(new_n729), .C1(new_n816), .C2(new_n756), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G137), .B2(new_n741), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n219), .B2(new_n748), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(G143), .C2(new_n744), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n222), .B2(new_n738), .C1(new_n297), .C2(new_n750), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n815), .A2(G294), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT108), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n739), .B(G116), .C1(new_n984), .C2(KEYINPUT46), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n738), .B2(new_n486), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n799), .A2(new_n820), .B1(new_n729), .B2(new_n432), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n750), .A2(new_n478), .B1(new_n740), .B2(new_n734), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n988), .A2(new_n252), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n747), .B2(new_n726), .C1(new_n497), .C2(new_n748), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n982), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n722), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n936), .A2(new_n773), .A3(new_n937), .ZN(new_n996));
  INV_X1    g0796(.A(new_n428), .ZN(new_n997));
  INV_X1    g0797(.A(new_n768), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n766), .B1(new_n209), .B2(new_n997), .C1(new_n242), .C2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n718), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n976), .A2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n676), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n295), .A2(G50), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n467), .C1(new_n214), .C2(new_n219), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1002), .B1(new_n1005), .B2(new_n328), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n238), .A2(new_n467), .A3(new_n252), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n209), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n766), .C1(new_n432), .C2(new_n209), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n718), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n733), .A2(new_n295), .B1(new_n726), .B2(new_n214), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT110), .Z(new_n1012));
  OAI22_X1  g0812(.A1(new_n738), .A2(new_n219), .B1(new_n297), .B2(new_n740), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT109), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n252), .B1(new_n750), .B2(new_n347), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n730), .A2(new_n428), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n493), .B2(new_n748), .C1(new_n756), .C2(new_n799), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n815), .A2(G311), .B1(G317), .B2(new_n795), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n478), .B2(new_n726), .C1(new_n749), .C2(new_n799), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT48), .Z(new_n1023));
  NOR2_X1   g0823(.A1(new_n729), .A2(new_n747), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n738), .A2(new_n824), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n806), .A2(G116), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n741), .A2(G326), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n328), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1010), .B1(new_n1032), .B2(new_n722), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n668), .B2(new_n774), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1035), .A2(new_n1036), .B1(new_n717), .B2(new_n968), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n713), .A2(new_n968), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n674), .A3(new_n969), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(G393));
  NAND2_X1  g0840(.A1(new_n965), .A2(new_n717), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n815), .A2(G303), .B1(G116), .B2(new_n730), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT113), .Z(new_n1043));
  AOI211_X1 g0843(.A(new_n753), .B(new_n1043), .C1(G322), .C2(new_n741), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n727), .A2(G294), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n739), .A2(G283), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n744), .A2(G317), .B1(new_n795), .B2(G311), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n252), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n427), .A2(new_n727), .B1(new_n730), .B2(G77), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n816), .B2(new_n347), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT112), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n328), .B(new_n1053), .C1(G143), .C2(new_n741), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n811), .C1(new_n214), .C2(new_n738), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n744), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT51), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1050), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n722), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n946), .A2(new_n765), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n766), .B1(new_n209), .B2(new_n497), .C1(new_n998), .C2(new_n249), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1059), .A2(new_n718), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1041), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n971), .A2(new_n973), .B1(new_n972), .B2(new_n969), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n674), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(G390));
  AND3_X1   g0866(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT79), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT79), .B1(new_n446), .B2(new_n449), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n339), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n834), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n840), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G330), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n783), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n893), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n710), .A3(G330), .A4(new_n786), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n687), .A2(new_n657), .A3(new_n780), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n782), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT115), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1073), .B1(new_n846), .B2(new_n850), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n905), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT115), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1076), .A2(new_n782), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1075), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n787), .A2(new_n782), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n893), .A2(G330), .A3(new_n841), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1071), .B1(new_n712), .B2(new_n786), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n459), .A2(new_n893), .A3(G330), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n897), .A2(new_n1091), .A3(new_n648), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1085), .A2(new_n1071), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n912), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n911), .A2(new_n913), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT114), .B1(new_n906), .B2(new_n912), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1097), .B(new_n889), .C1(new_n1082), .C2(new_n905), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1086), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1075), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1094), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1092), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1087), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1107), .A2(new_n674), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n717), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n750), .A2(new_n486), .B1(new_n740), .B2(new_n824), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n738), .A2(new_n596), .B1(new_n219), .B2(new_n729), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n252), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n816), .B2(new_n432), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1115), .B(new_n1118), .C1(G68), .C2(new_n806), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n747), .B2(new_n799), .C1(new_n497), .C2(new_n726), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n739), .A2(G150), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n328), .B(new_n1122), .C1(G159), .C2(new_n730), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n741), .A2(G125), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n815), .A2(G137), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n727), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n808), .B2(new_n750), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G128), .B2(new_n744), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n748), .A2(new_n347), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1120), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1099), .A2(new_n763), .B1(new_n722), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n827), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n718), .B1(new_n427), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT116), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1112), .A2(new_n1114), .A3(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1092), .B1(new_n1113), .B2(new_n1108), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n303), .A2(new_n656), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT55), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n309), .B2(new_n312), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n309), .A2(new_n1145), .A3(new_n312), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1148), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1144), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1150), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1143), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1150), .B2(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(new_n1148), .A3(new_n1144), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n1142), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n890), .A2(KEYINPUT40), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n893), .A2(new_n842), .A3(new_n882), .A4(new_n841), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1160), .A2(G330), .A3(new_n916), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n916), .B1(new_n1160), .B2(G330), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n917), .B1(new_n891), .B2(new_n1072), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1160), .A2(G330), .A3(new_n916), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1157), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1140), .B1(new_n1141), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1111), .A2(new_n1093), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1161), .A2(new_n1162), .A3(new_n1157), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1166), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n1173), .A3(KEYINPUT57), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1169), .A2(new_n1174), .A3(new_n674), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n717), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n718), .B1(G50), .B2(new_n1135), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n806), .A2(G58), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n219), .B2(new_n738), .C1(new_n486), .C2(new_n799), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n997), .A2(new_n726), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n252), .B1(new_n741), .B2(G283), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n465), .C1(new_n432), .C2(new_n750), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n733), .A2(new_n493), .B1(new_n729), .B2(new_n214), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT118), .Z(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n465), .B1(new_n326), .B2(new_n288), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1185), .A2(new_n1186), .B1(new_n347), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT119), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n726), .A2(new_n798), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1127), .B2(new_n739), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n793), .A2(G132), .B1(new_n730), .B2(G150), .ZN(new_n1192));
  INV_X1    g0992(.A(G128), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1192), .C1(new_n1193), .C2(new_n750), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G125), .B2(new_n744), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n288), .B(new_n465), .C1(new_n748), .C2(new_n756), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G124), .B2(new_n741), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1189), .B(new_n1200), .C1(new_n1186), .C2(new_n1185), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1177), .B1(new_n1201), .B2(new_n722), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1166), .B2(new_n764), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1176), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1175), .A2(new_n1204), .ZN(G375));
  OAI221_X1 g1005(.A(new_n1017), .B1(new_n219), .B2(new_n748), .C1(new_n816), .C2(new_n486), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n740), .A2(new_n478), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n799), .A2(new_n824), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G283), .A2(new_n795), .B1(new_n727), .B2(G107), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n328), .C1(new_n493), .C2(new_n738), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n815), .A2(new_n1127), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n730), .A2(G50), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1212), .A2(new_n252), .A3(new_n1178), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n740), .A2(new_n1193), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n799), .A2(new_n808), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G137), .A2(new_n795), .B1(new_n727), .B2(G150), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n756), .B2(new_n738), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n722), .B1(new_n1211), .B2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n718), .C1(G68), .C2(new_n1135), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n905), .B2(new_n763), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n716), .B(KEYINPUT122), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1090), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1084), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n950), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1226), .B2(new_n1108), .ZN(G381));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1175), .A3(new_n1204), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(G384), .A3(G381), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n976), .A2(new_n1065), .A3(new_n1000), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1037), .A2(new_n776), .A3(new_n1039), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .ZN(G407));
  INV_X1    g1034(.A(G343), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G213), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT123), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(new_n1229), .C2(new_n1238), .ZN(G409));
  NAND2_X1  g1039(.A1(G375), .A2(G378), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1225), .A2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1084), .A2(KEYINPUT60), .A3(new_n1089), .A4(new_n1092), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(new_n1094), .A3(new_n674), .A4(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1244), .A2(G384), .A3(new_n1224), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1244), .B2(new_n1224), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1173), .A2(new_n1223), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1248), .A2(new_n1203), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1170), .A2(new_n1173), .A3(new_n950), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1170), .A2(new_n1173), .A3(KEYINPUT124), .A4(new_n950), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1228), .A2(new_n1249), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1240), .A2(new_n1238), .A3(new_n1247), .A4(new_n1254), .ZN(new_n1255));
  XOR2_X1   g1055(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1240), .A2(new_n1238), .A3(new_n1254), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1245), .A2(new_n1246), .A3(KEYINPUT125), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT125), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1237), .A2(G2897), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(KEYINPUT125), .B(new_n1261), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1259), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1237), .B1(G375), .B2(G378), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1247), .A4(new_n1254), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1257), .A2(new_n1266), .A3(new_n1267), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1232), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1065), .B1(new_n976), .B2(new_n1000), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1231), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n976), .A2(new_n1065), .A3(new_n1000), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1272), .A2(new_n1232), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT126), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1274), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1278), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1271), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1282), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1247), .A4(new_n1254), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1255), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1286), .B(new_n1287), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1285), .A2(new_n1291), .ZN(G405));
  NAND2_X1  g1092(.A1(new_n1240), .A2(new_n1229), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1293), .A2(new_n1247), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1247), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1283), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1284), .A2(new_n1295), .A3(new_n1294), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G402));
endmodule


