

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XNOR2_X1 U322 ( .A(n390), .B(n291), .ZN(n393) );
  XOR2_X1 U323 ( .A(n417), .B(n416), .Z(n290) );
  AND2_X1 U324 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U325 ( .A(G127GAT), .B(KEYINPUT85), .Z(n292) );
  INV_X1 U326 ( .A(KEYINPUT33), .ZN(n420) );
  XNOR2_X1 U327 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U328 ( .A(n423), .B(n422), .ZN(n427) );
  XNOR2_X1 U329 ( .A(n393), .B(n392), .ZN(n398) );
  XNOR2_X1 U330 ( .A(n403), .B(KEYINPUT100), .ZN(n564) );
  XOR2_X1 U331 ( .A(n571), .B(KEYINPUT41), .Z(n558) );
  XNOR2_X1 U332 ( .A(n400), .B(n399), .ZN(n525) );
  INV_X1 U333 ( .A(G29GAT), .ZN(n450) );
  XNOR2_X1 U334 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n474) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U336 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n453), .B(n452), .ZN(G1328GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT6), .B(KEYINPUT96), .Z(n294) );
  XNOR2_X1 U339 ( .A(G1GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n302) );
  XOR2_X1 U341 ( .A(KEYINPUT97), .B(KEYINPUT4), .Z(n300) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n292), .B(n295), .ZN(n391) );
  XOR2_X1 U344 ( .A(KEYINPUT2), .B(KEYINPUT95), .Z(n297) );
  XNOR2_X1 U345 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U347 ( .A(G141GAT), .B(n298), .Z(n366) );
  XNOR2_X1 U348 ( .A(n391), .B(n366), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n314) );
  NAND2_X1 U351 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XOR2_X1 U352 ( .A(KEYINPUT78), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(G120GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U355 ( .A(G134GAT), .B(G162GAT), .Z(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U358 ( .A(G57GAT), .B(KEYINPUT1), .Z(n310) );
  XNOR2_X1 U359 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n542) );
  XOR2_X1 U363 ( .A(KEYINPUT75), .B(KEYINPUT66), .Z(n316) );
  XNOR2_X1 U364 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n334) );
  XOR2_X1 U366 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n318) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U369 ( .A(G106GAT), .B(G99GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(G190GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U372 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U373 ( .A(G43GAT), .B(G134GAT), .Z(n387) );
  XOR2_X1 U374 ( .A(G85GAT), .B(G92GAT), .Z(n417) );
  XOR2_X1 U375 ( .A(G50GAT), .B(G162GAT), .Z(n354) );
  XNOR2_X1 U376 ( .A(n417), .B(n354), .ZN(n324) );
  AND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n387), .B(n325), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n328), .B(KEYINPUT77), .Z(n332) );
  XOR2_X1 U382 ( .A(G29GAT), .B(KEYINPUT8), .Z(n330) );
  XNOR2_X1 U383 ( .A(KEYINPUT7), .B(KEYINPUT71), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n436) );
  XNOR2_X1 U385 ( .A(n436), .B(KEYINPUT78), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U387 ( .A(n334), .B(n333), .Z(n477) );
  INV_X1 U388 ( .A(n477), .ZN(n550) );
  XNOR2_X1 U389 ( .A(KEYINPUT36), .B(n550), .ZN(n577) );
  XOR2_X1 U390 ( .A(G78GAT), .B(G211GAT), .Z(n336) );
  XNOR2_X1 U391 ( .A(G71GAT), .B(G155GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .Z(n429) );
  XOR2_X1 U394 ( .A(n337), .B(n429), .Z(n339) );
  XNOR2_X1 U395 ( .A(G183GAT), .B(G127GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U397 ( .A(G15GAT), .B(G22GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n340), .B(G1GAT), .ZN(n433) );
  XOR2_X1 U399 ( .A(n433), .B(KEYINPUT12), .Z(n342) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n344), .B(n343), .Z(n352) );
  XOR2_X1 U403 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n346) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(G64GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U406 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X1 U407 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n575) );
  INV_X1 U411 ( .A(n542), .ZN(n409) );
  XNOR2_X1 U412 ( .A(G106GAT), .B(G78GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n353), .B(G148GAT), .ZN(n416) );
  XOR2_X1 U414 ( .A(KEYINPUT22), .B(n416), .Z(n356) );
  XNOR2_X1 U415 ( .A(G22GAT), .B(n354), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U417 ( .A(G211GAT), .B(KEYINPUT21), .Z(n358) );
  XNOR2_X1 U418 ( .A(G197GAT), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n370) );
  XOR2_X1 U420 ( .A(n370), .B(KEYINPUT94), .Z(n360) );
  NAND2_X1 U421 ( .A1(G228GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U423 ( .A(n362), .B(n361), .Z(n368) );
  XOR2_X1 U424 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n364) );
  XNOR2_X1 U425 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n471) );
  XNOR2_X1 U429 ( .A(n471), .B(KEYINPUT68), .ZN(n369) );
  XOR2_X1 U430 ( .A(n369), .B(KEYINPUT28), .Z(n521) );
  AND2_X1 U431 ( .A1(n409), .A2(n521), .ZN(n386) );
  XOR2_X1 U432 ( .A(G204GAT), .B(G64GAT), .Z(n428) );
  XOR2_X1 U433 ( .A(n428), .B(n370), .Z(n372) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U436 ( .A(n373), .B(KEYINPUT99), .Z(n375) );
  XOR2_X1 U437 ( .A(G36GAT), .B(G8GAT), .Z(n432) );
  XNOR2_X1 U438 ( .A(n432), .B(G92GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n384) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(G176GAT), .ZN(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n377) );
  XNOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U444 ( .A(n378), .B(KEYINPUT19), .Z(n380) );
  XNOR2_X1 U445 ( .A(G190GAT), .B(G183GAT), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n400) );
  INV_X1 U448 ( .A(n400), .ZN(n383) );
  XOR2_X1 U449 ( .A(n384), .B(n383), .Z(n515) );
  INV_X1 U450 ( .A(n515), .ZN(n467) );
  XOR2_X1 U451 ( .A(n467), .B(KEYINPUT27), .Z(n404) );
  INV_X1 U452 ( .A(n404), .ZN(n385) );
  NAND2_X1 U453 ( .A1(n386), .A2(n385), .ZN(n524) );
  XNOR2_X1 U454 ( .A(n387), .B(KEYINPUT90), .ZN(n389) );
  XNOR2_X1 U455 ( .A(G99GAT), .B(G71GAT), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n388), .B(G120GAT), .ZN(n419) );
  XNOR2_X1 U457 ( .A(n389), .B(n419), .ZN(n390) );
  XOR2_X1 U458 ( .A(n391), .B(KEYINPUT86), .Z(n392) );
  XOR2_X1 U459 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n395) );
  XNOR2_X1 U460 ( .A(KEYINPUT65), .B(KEYINPUT89), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U462 ( .A(G15GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U464 ( .A(KEYINPUT92), .B(n525), .Z(n401) );
  NOR2_X1 U465 ( .A1(n524), .A2(n401), .ZN(n412) );
  NAND2_X1 U466 ( .A1(n525), .A2(n471), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT26), .ZN(n403) );
  NOR2_X1 U468 ( .A1(n564), .A2(n404), .ZN(n540) );
  NOR2_X1 U469 ( .A1(n525), .A2(n515), .ZN(n405) );
  NOR2_X1 U470 ( .A1(n471), .A2(n405), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n406), .B(KEYINPUT25), .ZN(n407) );
  XNOR2_X1 U472 ( .A(KEYINPUT101), .B(n407), .ZN(n408) );
  NOR2_X1 U473 ( .A1(n540), .A2(n408), .ZN(n410) );
  NOR2_X1 U474 ( .A1(n410), .A2(n409), .ZN(n411) );
  NOR2_X1 U475 ( .A1(n412), .A2(n411), .ZN(n476) );
  NOR2_X1 U476 ( .A1(n575), .A2(n476), .ZN(n413) );
  NAND2_X1 U477 ( .A1(n577), .A2(n413), .ZN(n414) );
  XNOR2_X1 U478 ( .A(KEYINPUT106), .B(n414), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n415), .B(KEYINPUT37), .ZN(n510) );
  NAND2_X1 U480 ( .A1(G230GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n290), .B(n418), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n419), .B(KEYINPUT74), .ZN(n421) );
  XOR2_X1 U483 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n425) );
  XNOR2_X1 U484 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n571) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U490 ( .A(G50GAT), .B(G43GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U492 ( .A(n436), .B(KEYINPUT69), .Z(n438) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n448) );
  XOR2_X1 U496 ( .A(G141GAT), .B(G197GAT), .Z(n442) );
  XNOR2_X1 U497 ( .A(G169GAT), .B(G113GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U499 ( .A(KEYINPUT72), .B(KEYINPUT30), .Z(n444) );
  XNOR2_X1 U500 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n566) );
  INV_X1 U504 ( .A(n566), .ZN(n499) );
  NOR2_X1 U505 ( .A1(n571), .A2(n499), .ZN(n481) );
  NAND2_X1 U506 ( .A1(n510), .A2(n481), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n449), .B(KEYINPUT38), .ZN(n497) );
  NOR2_X1 U508 ( .A1(n542), .A2(n497), .ZN(n453) );
  XNOR2_X1 U509 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n469) );
  XNOR2_X1 U511 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n466) );
  NAND2_X1 U512 ( .A1(n566), .A2(n558), .ZN(n454) );
  XNOR2_X1 U513 ( .A(KEYINPUT46), .B(n454), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n455), .A2(n477), .ZN(n456) );
  NOR2_X1 U515 ( .A1(n575), .A2(n456), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT47), .ZN(n464) );
  INV_X1 U517 ( .A(KEYINPUT67), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n575), .A2(n577), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT45), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n461), .A2(n571), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n462), .A2(n499), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n539) );
  NAND2_X1 U525 ( .A1(n467), .A2(n539), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n542), .A2(n470), .ZN(n565) );
  NOR2_X1 U528 ( .A1(n471), .A2(n565), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT55), .ZN(n473) );
  NOR2_X2 U530 ( .A1(n525), .A2(n473), .ZN(n561) );
  NAND2_X1 U531 ( .A1(n550), .A2(n561), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n575), .A2(n477), .ZN(n478) );
  XNOR2_X1 U533 ( .A(n478), .B(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U534 ( .A(n479), .B(KEYINPUT84), .ZN(n480) );
  NOR2_X1 U535 ( .A1(n476), .A2(n480), .ZN(n500) );
  NAND2_X1 U536 ( .A1(n481), .A2(n500), .ZN(n489) );
  NOR2_X1 U537 ( .A1(n542), .A2(n489), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT34), .B(n482), .Z(n483) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n515), .A2(n489), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT102), .B(n484), .Z(n485) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n485), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n525), .A2(n489), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NOR2_X1 U547 ( .A1(n521), .A2(n489), .ZN(n490) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(n490), .Z(n491) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  NOR2_X1 U550 ( .A1(n497), .A2(n515), .ZN(n493) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1329GAT) );
  NOR2_X1 U553 ( .A1(n497), .A2(n525), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U556 ( .A(G43GAT), .B(n496), .Z(G1330GAT) );
  NOR2_X1 U557 ( .A1(n497), .A2(n521), .ZN(n498) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  AND2_X1 U559 ( .A1(n499), .A2(n558), .ZN(n511) );
  NAND2_X1 U560 ( .A1(n511), .A2(n500), .ZN(n507) );
  NOR2_X1 U561 ( .A1(n542), .A2(n507), .ZN(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U565 ( .A1(n515), .A2(n507), .ZN(n504) );
  XOR2_X1 U566 ( .A(KEYINPUT110), .B(n504), .Z(n505) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(n505), .ZN(G1333GAT) );
  NOR2_X1 U568 ( .A1(n525), .A2(n507), .ZN(n506) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n521), .A2(n507), .ZN(n509) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n520) );
  NOR2_X1 U574 ( .A1(n542), .A2(n520), .ZN(n513) );
  XNOR2_X1 U575 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n515), .A2(n520), .ZN(n517) );
  XNOR2_X1 U579 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n525), .A2(n520), .ZN(n519) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n539), .A2(n526), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT115), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n535), .A2(n566), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT116), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U594 ( .A1(n535), .A2(n558), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n533) );
  NAND2_X1 U597 ( .A1(n535), .A2(n575), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U601 ( .A1(n535), .A2(n550), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n551), .A2(n566), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n545) );
  NAND2_X1 U609 ( .A1(n551), .A2(n558), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U613 ( .A1(n551), .A2(n575), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT120), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n549), .ZN(G1346GAT) );
  XOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT121), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n566), .A2(n561), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n557), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n575), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n578) );
  NAND2_X1 U631 ( .A1(n578), .A2(n566), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

