//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n205), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n208), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  OR3_X1    g0021(.A1(new_n208), .A2(KEYINPUT64), .A3(G13), .ZN(new_n222));
  OAI21_X1  g0022(.A(KEYINPUT64), .B1(new_n208), .B2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n221), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n210), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n257), .B1(new_n216), .B2(new_n255), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(G1), .B(G13), .C1(new_n252), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(G274), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n266), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(G226), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  OAI21_X1  g0078(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n252), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n279), .B1(new_n280), .B2(new_n282), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n227), .B1(new_n208), .B2(new_n252), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n266), .A2(KEYINPUT66), .A3(G13), .A4(G20), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n286), .A2(new_n287), .B1(new_n244), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(new_n287), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n228), .A2(G1), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(G50), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n277), .B1(new_n278), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n301), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(KEYINPUT9), .B1(G200), .B2(new_n275), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n275), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n301), .C1(G179), .C2(new_n275), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n252), .A2(new_n212), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT68), .B(G33), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n253), .B1(new_n312), .B2(new_n251), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G223), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G226), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT69), .B1(new_n317), .B2(new_n262), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n323), .B2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g0124(.A(new_n316), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(new_n252), .B2(new_n212), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n263), .ZN(new_n328));
  INV_X1    g0128(.A(G232), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n272), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n271), .A2(new_n330), .A3(G190), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n318), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n317), .A2(new_n262), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n269), .A2(new_n270), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n335), .A2(new_n265), .B1(new_n329), .B2(new_n272), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n210), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n281), .A2(G159), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n228), .B(new_n253), .C1(new_n312), .C2(new_n251), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n344), .B2(KEYINPUT7), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n324), .B2(new_n228), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT16), .B(new_n343), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n320), .A2(new_n322), .A3(new_n251), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n253), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n349), .A2(new_n351), .B1(new_n353), .B2(new_n346), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n343), .B1(new_n354), .B2(new_n210), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n348), .A2(new_n357), .A3(new_n287), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n296), .A2(new_n283), .A3(new_n298), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n292), .B2(new_n283), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n338), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n338), .A2(KEYINPUT17), .A3(new_n358), .A4(new_n360), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n271), .A2(new_n330), .A3(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n318), .A2(new_n328), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n307), .B1(new_n334), .B2(new_n336), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n358), .A2(new_n360), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT18), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n285), .A2(new_n216), .B1(new_n228), .B2(G68), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n282), .A2(new_n244), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n287), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT11), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n292), .A2(new_n210), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT12), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT67), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n296), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT67), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n387), .A2(G68), .A3(new_n299), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n271), .B1(G238), .B2(new_n273), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n255), .A2(G226), .A3(new_n256), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n258), .C2(new_n329), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n263), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G179), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n391), .A2(new_n398), .A3(new_n395), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n398), .B1(new_n391), .B2(new_n395), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n403), .B2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT14), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n397), .A2(new_n399), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(G169), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n390), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(G200), .B1(new_n401), .B2(new_n402), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n397), .A2(G190), .A3(new_n399), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n389), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n387), .A2(G77), .A3(new_n299), .ZN(new_n413));
  INV_X1    g0213(.A(new_n283), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n285), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n287), .B1(new_n216), .B2(new_n292), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n420), .B1(new_n205), .B2(new_n255), .C1(new_n258), .C2(new_n211), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n263), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n271), .B1(G244), .B2(new_n273), .ZN(new_n423));
  INV_X1    g0223(.A(G179), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n307), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(G200), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n422), .A2(new_n423), .A3(G190), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n413), .A4(new_n418), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n310), .A2(new_n376), .A3(new_n412), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G45), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G1), .ZN(new_n435));
  AND2_X1   g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  NOR2_X1   g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(G270), .A3(new_n262), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT5), .B(G41), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n440), .A2(new_n262), .A3(G274), .A4(new_n435), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT77), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n251), .B1(new_n320), .B2(new_n322), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(new_n256), .C1(new_n447), .C2(new_n319), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n253), .A2(new_n254), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G303), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n313), .A2(new_n452), .A3(G264), .A4(G1698), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G264), .A2(G1698), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT78), .B1(new_n324), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n446), .B1(new_n456), .B2(new_n262), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G200), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n266), .B2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n385), .A2(new_n386), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT79), .B1(new_n294), .B2(G116), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n290), .A2(new_n464), .A3(new_n459), .A4(new_n291), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n228), .C1(G33), .C2(new_n204), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n459), .A2(G20), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n287), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT20), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n287), .A3(KEYINPUT20), .A4(new_n468), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n463), .A2(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n462), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n458), .B(new_n475), .C1(new_n276), .C2(new_n457), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n457), .A2(new_n424), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n462), .B2(new_n474), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n307), .B1(new_n461), .B2(new_n473), .ZN(new_n480));
  AOI211_X1 g0280(.A(KEYINPUT80), .B(new_n479), .C1(new_n457), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n455), .A2(new_n453), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n448), .A2(new_n450), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n262), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n443), .A2(new_n445), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT21), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n476), .B(new_n478), .C1(new_n481), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n487), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n479), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT21), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(KEYINPUT81), .A3(new_n478), .A4(new_n476), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G244), .B(G1698), .C1(new_n447), .C2(new_n319), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n313), .A2(KEYINPUT73), .A3(G244), .A4(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n323), .A2(G116), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n313), .A2(G238), .A3(new_n256), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n263), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n435), .A2(new_n213), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n262), .ZN(new_n507));
  INV_X1    g0307(.A(new_n435), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n265), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n505), .A2(G190), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT75), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n505), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n504), .B2(new_n263), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(G190), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n228), .B(G68), .C1(new_n447), .C2(new_n319), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n284), .A2(G97), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n228), .B1(new_n393), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n212), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(new_n287), .B1(new_n292), .B2(new_n416), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n296), .B1(new_n266), .B2(G33), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G87), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n512), .A2(new_n514), .A3(new_n517), .A4(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT76), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n513), .A2(new_n307), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(new_n287), .ZN(new_n533));
  INV_X1    g0333(.A(new_n416), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n266), .A2(G33), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n297), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n292), .A2(new_n416), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT74), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n515), .A2(new_n424), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n532), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n530), .A2(new_n531), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n531), .B1(new_n530), .B2(new_n544), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n441), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n438), .A2(new_n262), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n218), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n313), .A2(G250), .A3(new_n256), .ZN(new_n552));
  OAI211_X1 g0352(.A(G257), .B(G1698), .C1(new_n447), .C2(new_n319), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n323), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n549), .B(new_n551), .C1(new_n555), .C2(new_n263), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n212), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n228), .B(new_n558), .C1(new_n447), .C2(new_n319), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n228), .A2(G87), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n449), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n323), .A2(new_n228), .A3(G116), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n205), .A2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n559), .A2(new_n561), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT24), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n565), .A2(new_n562), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n559), .A4(new_n561), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n295), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n294), .A2(G107), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT25), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n527), .A2(G107), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI22_X1  g0375(.A1(G169), .A2(new_n556), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n551), .B1(new_n555), .B2(new_n263), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n441), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(G179), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT82), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n571), .A2(new_n575), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n307), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n556), .A2(new_n424), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n571), .A2(new_n575), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(G200), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n276), .C2(new_n578), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n580), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT72), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT71), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n438), .A2(G257), .A3(new_n262), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n441), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n441), .A3(new_n591), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n217), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n255), .A2(new_n256), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n466), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n313), .A2(G244), .A3(new_n256), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n596), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n594), .B(new_n595), .C1(new_n602), .C2(new_n262), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n307), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n294), .A2(G97), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n527), .B2(G97), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT6), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n609), .B2(new_n522), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n350), .B1(new_n312), .B2(new_n251), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT7), .B1(new_n253), .B2(new_n352), .ZN(new_n615));
  OAI21_X1  g0415(.A(G107), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI211_X1 g0416(.A(KEYINPUT70), .B(new_n295), .C1(new_n613), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT70), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n281), .A2(G77), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT6), .B1(new_n206), .B2(new_n608), .ZN(new_n620));
  INV_X1    g0420(.A(new_n611), .ZN(new_n621));
  OAI21_X1  g0421(.A(G20), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n619), .B(new_n622), .C1(new_n354), .C2(new_n205), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n623), .B2(new_n287), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n606), .B1(new_n617), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n595), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n593), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n424), .C1(new_n262), .C2(new_n602), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n604), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n287), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT70), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n623), .A2(new_n618), .A3(new_n287), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n601), .A2(new_n596), .ZN(new_n634));
  INV_X1    g0434(.A(new_n600), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n262), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n594), .A2(new_n595), .ZN(new_n637));
  OAI21_X1  g0437(.A(G200), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n627), .B(G190), .C1(new_n262), .C2(new_n602), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n633), .A2(new_n638), .A3(new_n639), .A4(new_n606), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n590), .B1(new_n629), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n629), .A2(new_n640), .A3(new_n590), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n589), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n433), .A2(new_n497), .A3(new_n548), .A4(new_n643), .ZN(G372));
  AND3_X1   g0444(.A1(new_n515), .A2(new_n516), .A3(G190), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n529), .B1(new_n515), .B2(new_n333), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n516), .B1(new_n515), .B2(G190), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n532), .A2(new_n542), .A3(new_n543), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT76), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n604), .A2(new_n625), .A3(new_n628), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n545), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n511), .B(new_n529), .C1(new_n333), .C2(new_n515), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n544), .A2(new_n651), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n544), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n484), .A2(new_n485), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G179), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n475), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n493), .B2(new_n494), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT83), .B1(new_n576), .B2(new_n579), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT83), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n581), .A2(new_n582), .A3(new_n663), .A4(new_n584), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n588), .A2(new_n629), .A3(new_n640), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n544), .A2(new_n655), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n657), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n653), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n433), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  INV_X1    g0473(.A(new_n309), .ZN(new_n674));
  XNOR2_X1  g0474(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT18), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT18), .B1(new_n369), .B2(new_n370), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n373), .A2(new_n374), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n365), .A2(new_n411), .ZN(new_n682));
  INV_X1    g0482(.A(new_n428), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n406), .A2(new_n405), .A3(G169), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n400), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n686), .B2(new_n390), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n681), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n674), .B1(new_n688), .B2(new_n306), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n673), .A2(new_n689), .ZN(G369));
  NAND3_X1  g0490(.A1(new_n266), .A2(new_n228), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n497), .B1(new_n475), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n462), .B2(new_n474), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n661), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n589), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n586), .B2(new_n697), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n581), .A2(new_n584), .A3(new_n582), .A4(new_n696), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(G330), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n661), .A2(new_n696), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n701), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n696), .B(KEYINPUT87), .Z(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n665), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n224), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n523), .A2(G116), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n713), .A2(new_n266), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n231), .B2(new_n713), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  NAND3_X1  g0518(.A1(new_n661), .A2(new_n580), .A3(new_n585), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n669), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n650), .A2(new_n654), .A3(new_n545), .A4(new_n651), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n544), .A2(new_n651), .A3(new_n655), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n649), .B1(new_n722), .B2(KEYINPUT26), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT88), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(KEYINPUT88), .A3(new_n723), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n696), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n708), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n671), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n497), .A2(new_n548), .A3(new_n643), .A4(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n636), .A2(new_n637), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n515), .A3(new_n577), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT30), .B1(new_n659), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n577), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n603), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n477), .A2(new_n739), .A3(new_n740), .A4(new_n515), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n513), .A2(new_n578), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n603), .A2(new_n424), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(new_n658), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n747), .B2(new_n696), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n737), .B2(new_n741), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n749), .A2(new_n750), .A3(new_n730), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n734), .A2(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n729), .A2(new_n733), .B1(G330), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n718), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n712), .A2(new_n313), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G45), .B2(new_n230), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n249), .A2(new_n434), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n224), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n224), .A2(new_n255), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT90), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n759), .B1(G355), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(G1), .B(G13), .C1(new_n228), .C2(G169), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT91), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT92), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n762), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n228), .A2(G13), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n266), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n713), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT89), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n333), .A2(G190), .ZN(new_n779));
  OAI21_X1  g0579(.A(G20), .B1(new_n779), .B2(G179), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT93), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT94), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT94), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n204), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n228), .A2(G179), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n228), .A2(new_n424), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n276), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n787), .A2(new_n276), .A3(G200), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n244), .B1(new_n797), .B2(new_n205), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n794), .A2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n210), .B1(new_n801), .B2(new_n212), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n793), .A2(new_n788), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n779), .A2(new_n228), .A3(new_n424), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n255), .B1(new_n216), .B2(new_n803), .C1(new_n805), .C2(new_n339), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n792), .A2(new_n798), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n781), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G294), .ZN(new_n809));
  INV_X1    g0609(.A(new_n803), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G311), .A2(new_n810), .B1(new_n790), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G322), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n449), .C1(new_n812), .C2(new_n805), .ZN(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n796), .A2(new_n814), .B1(new_n801), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n800), .A2(new_n817), .B1(new_n797), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n813), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n786), .A2(new_n807), .B1(new_n809), .B2(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n778), .B1(new_n764), .B2(new_n821), .C1(new_n700), .C2(new_n768), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n700), .A2(G330), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n777), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n700), .A2(G330), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n428), .A2(KEYINPUT97), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n419), .A2(new_n696), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT97), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n419), .A2(new_n829), .A3(new_n425), .A4(new_n427), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n827), .A2(new_n431), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n683), .A2(new_n696), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n708), .B(new_n834), .C1(new_n653), .C2(new_n670), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n731), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n753), .A2(G330), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n776), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n764), .A2(new_n766), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT95), .Z(new_n843));
  OAI21_X1  g0643(.A(new_n776), .B1(new_n843), .B2(G77), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n255), .B1(new_n804), .B2(G294), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n459), .B2(new_n803), .C1(new_n846), .C2(new_n789), .ZN(new_n847));
  INV_X1    g0647(.A(new_n801), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n799), .A2(G283), .B1(new_n848), .B2(G107), .ZN(new_n849));
  INV_X1    g0649(.A(new_n797), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G87), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n815), .C2(new_n796), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n785), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n810), .A2(G159), .B1(new_n804), .B2(G143), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n796), .B2(new_n857), .C1(new_n280), .C2(new_n800), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n808), .A2(G58), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n244), .A2(new_n801), .B1(new_n797), .B2(new_n210), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n324), .B(new_n863), .C1(G132), .C2(new_n790), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n854), .A2(new_n855), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n764), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n844), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n833), .B2(new_n766), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n841), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  OAI211_X1 g0671(.A(G116), .B(new_n229), .C1(new_n612), .C2(KEYINPUT35), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n872), .A2(KEYINPUT98), .B1(KEYINPUT35), .B2(new_n612), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(KEYINPUT98), .B2(new_n872), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT36), .Z(new_n875));
  OR3_X1    g0675(.A1(new_n230), .A2(new_n216), .A3(new_n340), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n266), .B(G13), .C1(new_n876), .C2(new_n245), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n343), .B1(new_n345), .B2(new_n347), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n356), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n348), .A2(new_n287), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n360), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n694), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n365), .B2(new_n375), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n370), .A2(new_n884), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n371), .A2(new_n887), .A3(new_n361), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n883), .B1(new_n369), .B2(new_n884), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .A3(new_n361), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n879), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n885), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n677), .A2(new_n678), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n363), .A2(new_n364), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n890), .A4(new_n892), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n390), .A2(new_n696), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n408), .A2(new_n411), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n411), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n390), .B(new_n696), .C1(new_n686), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n827), .A2(new_n830), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n697), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT99), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n900), .B(new_n905), .C1(new_n835), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n681), .A2(new_n884), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(KEYINPUT100), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n887), .B1(new_n681), .B2(new_n365), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n887), .A2(new_n361), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n916), .B2(KEYINPUT85), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n888), .ZN(new_n918));
  INV_X1    g0718(.A(new_n916), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(KEYINPUT85), .A3(KEYINPUT37), .A4(new_n371), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n879), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n899), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n914), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n686), .A2(new_n390), .A3(new_n697), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n913), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT100), .B1(new_n910), .B2(new_n912), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n729), .A2(new_n433), .A3(new_n733), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n689), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(G330), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n905), .A2(new_n833), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n749), .A2(new_n750), .A3(new_n697), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n748), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n937), .B1(new_n734), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT101), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n923), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT40), .ZN(new_n943));
  NAND2_X1  g0743(.A1(KEYINPUT101), .A2(KEYINPUT40), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n940), .B(new_n944), .C1(KEYINPUT40), .C2(new_n900), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n734), .A2(new_n939), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n433), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n936), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n935), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n266), .B2(new_n772), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n935), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n878), .B1(new_n953), .B2(new_n954), .ZN(G367));
  INV_X1    g0755(.A(new_n770), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n756), .A2(new_n239), .B1(new_n712), .B2(new_n534), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n777), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n324), .B1(new_n796), .B2(new_n846), .ZN(new_n959));
  INV_X1    g0759(.A(G294), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n800), .A2(new_n960), .B1(new_n797), .B2(new_n204), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(G107), .C2(new_n808), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n790), .A2(G317), .B1(new_n804), .B2(G303), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n818), .B2(new_n803), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n848), .A2(G116), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n962), .B(new_n967), .C1(new_n965), .C2(new_n966), .ZN(new_n968));
  INV_X1    g0768(.A(new_n784), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(G68), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n449), .B1(G150), .B2(new_n804), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n244), .B2(new_n803), .C1(new_n857), .C2(new_n789), .ZN(new_n972));
  INV_X1    g0772(.A(G159), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n800), .A2(new_n973), .B1(new_n801), .B2(new_n339), .ZN(new_n974));
  INV_X1    g0774(.A(G143), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n796), .A2(new_n975), .B1(new_n797), .B2(new_n216), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n972), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n970), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n968), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT47), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n867), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(KEYINPUT47), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n958), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n529), .A2(new_n697), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n649), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n985), .B(KEYINPUT102), .C1(new_n668), .C2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(KEYINPUT102), .B2(new_n985), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n983), .B1(new_n987), .B2(new_n767), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n625), .A2(new_n708), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n629), .A2(new_n640), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n629), .B2(new_n730), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT103), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n709), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT45), .ZN(new_n995));
  NOR2_X1   g0795(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n996));
  INV_X1    g0796(.A(new_n993), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n710), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n709), .B(new_n993), .C1(KEYINPUT105), .C2(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(new_n705), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n995), .A2(new_n705), .A3(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n823), .A2(KEYINPUT106), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n707), .B1(new_n704), .B2(new_n706), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n754), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n754), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n713), .B(KEYINPUT41), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT107), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1010), .A2(KEYINPUT107), .A3(new_n1011), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1014), .A2(new_n773), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n993), .A2(new_n707), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT42), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n580), .A2(new_n585), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n997), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n708), .B1(new_n1020), .B2(new_n629), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT43), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1018), .A2(new_n1021), .B1(new_n1022), .B2(new_n987), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n987), .A2(new_n1022), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n705), .A2(new_n993), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(KEYINPUT104), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(KEYINPUT104), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n989), .B1(new_n1016), .B2(new_n1032), .ZN(G387));
  NAND3_X1  g0833(.A1(new_n702), .A2(new_n703), .A3(new_n767), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n810), .A2(G303), .B1(new_n804), .B2(G317), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n796), .B2(new_n812), .C1(new_n846), .C2(new_n800), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n808), .A2(G283), .B1(G294), .B2(new_n848), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n324), .B1(new_n814), .B2(new_n789), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G116), .B2(new_n850), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n784), .A2(new_n416), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n795), .A2(G159), .B1(new_n848), .B2(G77), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n283), .B2(new_n800), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G68), .A2(new_n810), .B1(new_n790), .B2(G150), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n244), .B2(new_n805), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n313), .B1(new_n204), .B2(new_n797), .ZN(new_n1053));
  OR4_X1    g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n764), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n761), .A2(new_n715), .B1(new_n205), .B2(new_n712), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n715), .C1(G68), .C2(G77), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT108), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(KEYINPUT108), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(KEYINPUT109), .A3(new_n756), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n434), .B2(new_n236), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT109), .B1(new_n1062), .B2(new_n756), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1056), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n777), .B(new_n1055), .C1(new_n956), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1008), .A2(new_n774), .B1(new_n1034), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1009), .A2(new_n713), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1008), .A2(new_n754), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  AOI22_X1  g0871(.A1(new_n795), .A2(G150), .B1(G159), .B2(new_n804), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT51), .Z(new_n1073));
  OAI221_X1 g0873(.A(new_n851), .B1(new_n210), .B2(new_n801), .C1(new_n800), .C2(new_n244), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n803), .A2(new_n283), .B1(new_n789), .B2(new_n975), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1074), .A2(new_n324), .A3(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1073), .B(new_n1076), .C1(new_n784), .C2(new_n216), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n795), .A2(G317), .B1(G311), .B2(new_n804), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n808), .A2(G116), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n449), .B1(new_n803), .B2(new_n960), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G322), .B2(new_n790), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n800), .A2(new_n815), .B1(new_n797), .B2(new_n205), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G283), .B2(new_n848), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n764), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n756), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n956), .B1(new_n204), .B2(new_n224), .C1(new_n243), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n777), .B1(new_n1088), .B2(KEYINPUT110), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(KEYINPUT110), .B2(new_n1088), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1086), .B(new_n1090), .C1(new_n993), .C2(new_n767), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1005), .B2(new_n773), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n713), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(G390));
  OAI21_X1  g0899(.A(new_n905), .B1(new_n835), .B2(new_n909), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n925), .B1(new_n1100), .B2(new_n926), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n906), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n431), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n696), .B(new_n1103), .C1(new_n726), .C2(new_n727), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n907), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n905), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n926), .B(KEYINPUT111), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n923), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1101), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n833), .A2(G330), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n948), .A2(new_n905), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT112), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT112), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n948), .A2(new_n1115), .A3(new_n905), .A4(new_n1112), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT113), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1103), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1105), .B1(new_n728), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n905), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1109), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1101), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1111), .B(new_n1122), .C1(new_n734), .C2(new_n752), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT113), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n724), .A2(new_n725), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n720), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n727), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n697), .A3(new_n1120), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n907), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1108), .B1(new_n1133), .B2(new_n905), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1128), .B(new_n1117), .C1(new_n1134), .C2(new_n1101), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1119), .A2(new_n774), .A3(new_n1127), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(new_n1128), .B1(new_n1110), .B2(new_n1126), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n774), .A4(new_n1119), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n800), .A2(new_n857), .B1(new_n803), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n969), .B2(G159), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n848), .A2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n449), .B1(new_n790), .B2(G125), .ZN(new_n1149));
  INV_X1    g0949(.A(G132), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n805), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n796), .A2(new_n1152), .B1(new_n797), .B2(new_n244), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1146), .A2(new_n1148), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n790), .A2(G294), .B1(new_n804), .B2(G116), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n449), .C1(new_n204), .C2(new_n803), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n848), .A2(G87), .B1(new_n850), .B2(G68), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n205), .B2(new_n800), .C1(new_n818), .C2(new_n796), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(new_n969), .C2(G77), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n867), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n776), .C1(new_n414), .C2(new_n843), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n925), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n765), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n753), .A2(new_n1112), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1122), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1114), .A2(new_n1116), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n836), .A2(new_n908), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n905), .B1(new_n948), .B2(new_n1112), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(new_n1125), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1168), .A2(new_n1169), .B1(new_n1121), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT114), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n949), .B2(new_n936), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n948), .A2(new_n433), .A3(KEYINPUT114), .A4(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n933), .A2(new_n1176), .A3(new_n689), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1135), .A2(new_n1127), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1128), .B1(new_n1181), .B2(new_n1117), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1119), .A2(new_n1127), .A3(new_n1135), .A4(new_n1178), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n713), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1142), .A2(new_n1165), .A3(new_n1185), .ZN(G378));
  INV_X1    g0986(.A(new_n1177), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n946), .A2(G330), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n929), .A2(new_n1189), .A3(new_n931), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n301), .A2(new_n884), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n310), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  AOI21_X1  g0994(.A(new_n936), .B1(new_n943), .B2(new_n945), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n913), .A2(new_n928), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n930), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1190), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1194), .B1(new_n1190), .B2(new_n1197), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n713), .B1(new_n1188), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1194), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1197), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1196), .A2(new_n1195), .A3(new_n930), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1190), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1201), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n774), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n776), .B1(G50), .B2(new_n842), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n324), .A2(new_n261), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n244), .C1(G33), .C2(G41), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n970), .B1(new_n459), .B2(new_n796), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT119), .Z(new_n1216));
  OAI22_X1  g1016(.A1(new_n801), .A2(new_n216), .B1(new_n789), .B2(new_n818), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1217), .B(new_n1213), .C1(G58), .C2(new_n850), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT118), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n810), .A2(new_n534), .B1(new_n804), .B2(G107), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n204), .B2(new_n800), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1216), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1214), .B1(new_n1222), .B2(KEYINPUT58), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT120), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT120), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n805), .A2(new_n1152), .B1(new_n803), .B2(new_n857), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G132), .B2(new_n799), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1143), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n795), .A2(G125), .B1(new_n848), .B2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(new_n784), .C2(new_n280), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n973), .B2(new_n797), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1230), .B2(KEYINPUT59), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1222), .A2(KEYINPUT58), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1224), .A2(new_n1225), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1212), .B1(new_n1236), .B2(new_n867), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1202), .B2(new_n766), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1211), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1210), .A2(new_n1240), .ZN(G375));
  OR2_X1    g1041(.A1(new_n1172), .A2(new_n773), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT121), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n776), .B1(new_n843), .B2(G68), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n799), .A2(G116), .B1(new_n850), .B2(G77), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n795), .A2(G294), .B1(new_n848), .B2(G97), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n255), .B1(new_n790), .B2(G303), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n810), .A2(G107), .B1(new_n804), .B2(G283), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n784), .A2(new_n244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n795), .A2(G132), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n803), .A2(new_n280), .B1(new_n789), .B2(new_n1152), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G137), .B2(new_n804), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n324), .B1(G58), .B2(new_n850), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n799), .A2(new_n1228), .B1(new_n848), .B2(G159), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1048), .A2(new_n1249), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1244), .B1(new_n1258), .B2(new_n867), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n905), .B2(new_n766), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1242), .A2(KEYINPUT121), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1243), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1179), .A2(new_n1011), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(G381));
  NOR4_X1   g1065(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1267));
  OR4_X1    g1067(.A1(G387), .A2(new_n1267), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  INV_X1    g1070(.A(G213), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(G343), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n695), .A2(KEYINPUT123), .A3(G213), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT124), .Z(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G375), .C2(new_n1276), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1240), .C1(new_n1201), .C2(new_n1209), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1119), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1095), .B1(new_n1280), .B2(new_n1179), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1164), .B1(new_n1281), .B2(new_n1184), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1207), .A2(new_n1208), .A3(new_n1011), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1142), .B(new_n1282), .C1(new_n1283), .C2(new_n1239), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1279), .A2(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1263), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT60), .B1(new_n1263), .B2(KEYINPUT125), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n713), .B(new_n1179), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1262), .A2(G384), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1262), .B2(new_n1288), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AND4_X1   g1092(.A1(KEYINPUT126), .A2(new_n1285), .A3(new_n1274), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1274), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT126), .B1(new_n1295), .B2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1278), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1291), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1298), .A2(new_n1289), .B1(G2897), .B2(new_n1275), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1294), .A2(G2897), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1292), .B2(new_n1300), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1301), .A2(new_n1295), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G390), .B(new_n989), .C1(new_n1016), .C2(new_n1032), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n774), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1032), .B1(new_n1304), .B2(new_n1015), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1098), .B1(new_n1305), .B2(new_n988), .ZN(new_n1306));
  XOR2_X1   g1106(.A(G393), .B(G396), .Z(new_n1307));
  AND3_X1   g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1308), .A2(new_n1309), .A3(KEYINPUT61), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1275), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(KEYINPUT63), .A3(new_n1292), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1297), .A2(new_n1302), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1301), .B2(new_n1311), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1311), .A2(KEYINPUT62), .A3(new_n1292), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1315), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1313), .B1(new_n1319), .B2(new_n1320), .ZN(G405));
  INV_X1    g1121(.A(new_n1292), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G378), .B1(new_n1210), .B2(new_n1240), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1322), .B1(new_n1324), .B2(new_n1279), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1279), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1323), .A2(new_n1326), .A3(new_n1292), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1320), .ZN(G402));
endmodule


