

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762;

  NAND2_X1 U378 ( .A1(n637), .A2(n704), .ZN(n372) );
  XNOR2_X1 U379 ( .A(n592), .B(n398), .ZN(n637) );
  NOR2_X1 U380 ( .A1(n661), .A2(n573), .ZN(n574) );
  XNOR2_X1 U381 ( .A(n405), .B(n404), .ZN(n559) );
  NOR2_X1 U382 ( .A1(G902), .A2(n646), .ZN(n511) );
  XOR2_X1 U383 ( .A(G122), .B(G104), .Z(n499) );
  XNOR2_X2 U384 ( .A(n355), .B(n444), .ZN(n638) );
  NAND2_X2 U385 ( .A1(n443), .A2(n426), .ZN(n355) );
  AND2_X2 U386 ( .A1(n636), .A2(n390), .ZN(n357) );
  NOR2_X2 U387 ( .A1(G902), .A2(n721), .ZN(n484) );
  AND2_X2 U388 ( .A1(n408), .A2(n407), .ZN(n550) );
  AND2_X2 U389 ( .A1(n389), .A2(n388), .ZN(n387) );
  XOR2_X1 U390 ( .A(G137), .B(G140), .Z(n522) );
  XNOR2_X1 U391 ( .A(n579), .B(KEYINPUT39), .ZN(n591) );
  NAND2_X4 U392 ( .A1(n387), .A2(n384), .ZN(n631) );
  INV_X2 U393 ( .A(n604), .ZN(n675) );
  XNOR2_X2 U394 ( .A(n383), .B(n515), .ZN(n742) );
  INV_X1 U395 ( .A(n679), .ZN(n356) );
  INV_X1 U396 ( .A(n583), .ZN(n519) );
  XNOR2_X1 U397 ( .A(n428), .B(KEYINPUT87), .ZN(n625) );
  AND2_X1 U398 ( .A1(n578), .A2(n371), .ZN(n566) );
  INV_X1 U399 ( .A(KEYINPUT84), .ZN(n398) );
  NAND2_X1 U400 ( .A1(n624), .A2(n625), .ZN(n370) );
  XNOR2_X1 U401 ( .A(n400), .B(KEYINPUT46), .ZN(n588) );
  NAND2_X1 U402 ( .A1(n402), .A2(n401), .ZN(n400) );
  XNOR2_X1 U403 ( .A(n599), .B(n454), .ZN(n606) );
  NOR2_X1 U404 ( .A1(n693), .A2(n694), .ZN(n585) );
  XNOR2_X1 U405 ( .A(n533), .B(n532), .ZN(n679) );
  NOR2_X1 U406 ( .A1(G902), .A2(n729), .ZN(n533) );
  XNOR2_X1 U407 ( .A(n494), .B(n483), .ZN(n721) );
  XNOR2_X1 U408 ( .A(n445), .B(n528), .ZN(n729) );
  XNOR2_X1 U409 ( .A(n494), .B(n495), .ZN(n648) );
  XNOR2_X1 U410 ( .A(n410), .B(n409), .ZN(n527) );
  XNOR2_X1 U411 ( .A(n478), .B(n395), .ZN(n482) );
  XNOR2_X1 U412 ( .A(n522), .B(n396), .ZN(n395) );
  XOR2_X1 U413 ( .A(G116), .B(G107), .Z(n514) );
  INV_X2 U414 ( .A(KEYINPUT68), .ZN(n365) );
  NAND2_X1 U415 ( .A1(n369), .A2(n357), .ZN(n368) );
  XNOR2_X1 U416 ( .A(n370), .B(n424), .ZN(n369) );
  INV_X1 U417 ( .A(KEYINPUT73), .ZN(n380) );
  INV_X1 U418 ( .A(KEYINPUT22), .ZN(n382) );
  INV_X1 U419 ( .A(n603), .ZN(n375) );
  INV_X1 U420 ( .A(KEYINPUT6), .ZN(n392) );
  INV_X1 U421 ( .A(KEYINPUT8), .ZN(n409) );
  NAND2_X1 U422 ( .A1(n537), .A2(G234), .ZN(n410) );
  NAND2_X1 U423 ( .A1(n371), .A2(n691), .ZN(n558) );
  NAND2_X1 U424 ( .A1(n418), .A2(n416), .ZN(n415) );
  NOR2_X1 U425 ( .A1(n417), .A2(n731), .ZN(n416) );
  NAND2_X1 U426 ( .A1(n728), .A2(n363), .ZN(n418) );
  NOR2_X1 U427 ( .A1(n360), .A2(G472), .ZN(n417) );
  NOR2_X1 U428 ( .A1(n663), .A2(n590), .ZN(n695) );
  INV_X1 U429 ( .A(KEYINPUT10), .ZN(n452) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT11), .ZN(n500) );
  INV_X1 U431 ( .A(G902), .ZN(n386) );
  NAND2_X1 U432 ( .A1(n496), .A2(G902), .ZN(n388) );
  XNOR2_X1 U433 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n607) );
  AND2_X1 U434 ( .A1(n554), .A2(n663), .ZN(n407) );
  XNOR2_X1 U435 ( .A(n617), .B(n391), .ZN(n619) );
  INV_X1 U436 ( .A(KEYINPUT79), .ZN(n391) );
  NAND2_X1 U437 ( .A1(n374), .A2(n373), .ZN(n622) );
  NAND2_X1 U438 ( .A1(n375), .A2(n359), .ZN(n374) );
  NAND2_X1 U439 ( .A1(n378), .A2(n377), .ZN(n376) );
  OR2_X1 U440 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U441 ( .A(n414), .B(KEYINPUT30), .ZN(n565) );
  XNOR2_X1 U442 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U443 ( .A(KEYINPUT94), .ZN(n471) );
  INV_X1 U444 ( .A(G478), .ZN(n404) );
  OR2_X1 U445 ( .A1(n726), .A2(G902), .ZN(n405) );
  XNOR2_X1 U446 ( .A(n510), .B(G475), .ZN(n453) );
  XNOR2_X1 U447 ( .A(n525), .B(n447), .ZN(n446) );
  NAND2_X1 U448 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U449 ( .A1(G953), .A2(G237), .ZN(n504) );
  XNOR2_X1 U450 ( .A(n497), .B(KEYINPUT69), .ZN(n383) );
  INV_X1 U451 ( .A(KEYINPUT44), .ZN(n424) );
  NOR2_X1 U452 ( .A1(n425), .A2(n358), .ZN(n390) );
  INV_X1 U453 ( .A(n651), .ZN(n425) );
  INV_X1 U454 ( .A(KEYINPUT86), .ZN(n444) );
  INV_X1 U455 ( .A(KEYINPUT76), .ZN(n396) );
  XOR2_X1 U456 ( .A(KEYINPUT75), .B(G107), .Z(n480) );
  XNOR2_X1 U457 ( .A(G110), .B(G104), .ZN(n479) );
  XOR2_X1 U458 ( .A(KEYINPUT4), .B(G101), .Z(n476) );
  NAND2_X1 U459 ( .A1(n382), .A2(n380), .ZN(n378) );
  NAND2_X1 U460 ( .A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(n377) );
  NAND2_X1 U461 ( .A1(n382), .A2(KEYINPUT73), .ZN(n381) );
  NAND2_X1 U462 ( .A1(n380), .A2(KEYINPUT22), .ZN(n379) );
  BUF_X1 U463 ( .A(n707), .Z(n745) );
  XNOR2_X1 U464 ( .A(n422), .B(n421), .ZN(n493) );
  XNOR2_X1 U465 ( .A(G113), .B(KEYINPUT72), .ZN(n421) );
  XNOR2_X1 U466 ( .A(n423), .B(KEYINPUT3), .ZN(n422) );
  XNOR2_X1 U467 ( .A(KEYINPUT93), .B(G119), .ZN(n423) );
  XNOR2_X1 U468 ( .A(n526), .B(KEYINPUT23), .ZN(n447) );
  INV_X1 U469 ( .A(KEYINPUT64), .ZN(n411) );
  XNOR2_X1 U470 ( .A(G113), .B(G143), .ZN(n498) );
  NOR2_X1 U471 ( .A1(n707), .A2(n640), .ZN(n639) );
  XNOR2_X1 U472 ( .A(n666), .B(KEYINPUT106), .ZN(n590) );
  NAND2_X1 U473 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U474 ( .A1(G472), .A2(n386), .ZN(n385) );
  XNOR2_X1 U475 ( .A(n512), .B(n513), .ZN(n406) );
  NAND2_X1 U476 ( .A1(n728), .A2(G475), .ZN(n436) );
  XNOR2_X1 U477 ( .A(n550), .B(KEYINPUT113), .ZN(n551) );
  NOR2_X1 U478 ( .A1(n356), .A2(n620), .ZN(n621) );
  NAND2_X1 U479 ( .A1(n430), .A2(n429), .ZN(n658) );
  NOR2_X1 U480 ( .A1(n616), .A2(n356), .ZN(n429) );
  INV_X1 U481 ( .A(n615), .ZN(n430) );
  NOR2_X1 U482 ( .A1(n419), .A2(n415), .ZN(n650) );
  NOR2_X1 U483 ( .A1(n728), .A2(n360), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n413), .B(n412), .ZN(n730) );
  NAND2_X1 U485 ( .A1(n728), .A2(G217), .ZN(n413) );
  INV_X1 U486 ( .A(KEYINPUT56), .ZN(n448) );
  AND2_X1 U487 ( .A1(n717), .A2(n399), .ZN(n719) );
  AND2_X1 U488 ( .A1(n716), .A2(n737), .ZN(n399) );
  INV_X1 U489 ( .A(n426), .ZN(n673) );
  NOR2_X1 U490 ( .A1(n695), .A2(n635), .ZN(n358) );
  XNOR2_X1 U491 ( .A(n558), .B(KEYINPUT19), .ZN(n598) );
  NAND2_X1 U492 ( .A1(n381), .A2(n379), .ZN(n359) );
  XOR2_X1 U493 ( .A(n648), .B(KEYINPUT62), .Z(n360) );
  XNOR2_X1 U494 ( .A(KEYINPUT92), .B(n457), .ZN(n731) );
  INV_X1 U495 ( .A(n731), .ZN(n420) );
  XOR2_X1 U496 ( .A(n647), .B(KEYINPUT59), .Z(n361) );
  XOR2_X1 U497 ( .A(n720), .B(n455), .Z(n362) );
  AND2_X1 U498 ( .A1(n360), .A2(G472), .ZN(n363) );
  XOR2_X1 U499 ( .A(KEYINPUT60), .B(KEYINPUT66), .Z(n364) );
  INV_X1 U500 ( .A(G953), .ZN(n737) );
  AND2_X4 U501 ( .A1(n645), .A2(n372), .ZN(n728) );
  XNOR2_X1 U502 ( .A(n436), .B(n361), .ZN(n435) );
  XNOR2_X2 U503 ( .A(n365), .B(G131), .ZN(n497) );
  NAND2_X1 U504 ( .A1(n728), .A2(G210), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n366), .B(KEYINPUT74), .ZN(n632) );
  NAND2_X1 U506 ( .A1(n675), .A2(n676), .ZN(n366) );
  NAND2_X1 U507 ( .A1(n616), .A2(n691), .ZN(n414) );
  XNOR2_X2 U508 ( .A(n631), .B(KEYINPUT107), .ZN(n616) );
  NOR2_X1 U509 ( .A1(n367), .A2(n575), .ZN(n576) );
  XNOR2_X1 U510 ( .A(n574), .B(KEYINPUT81), .ZN(n367) );
  XNOR2_X1 U511 ( .A(n406), .B(n518), .ZN(n726) );
  NAND2_X1 U512 ( .A1(n435), .A2(n420), .ZN(n434) );
  OR2_X2 U513 ( .A1(n632), .A2(n617), .ZN(n608) );
  INV_X1 U514 ( .A(n758), .ZN(n401) );
  XNOR2_X2 U515 ( .A(n628), .B(n486), .ZN(n604) );
  XNOR2_X2 U516 ( .A(n484), .B(n485), .ZN(n628) );
  XNOR2_X2 U517 ( .A(n368), .B(KEYINPUT45), .ZN(n704) );
  XNOR2_X1 U518 ( .A(n371), .B(n577), .ZN(n690) );
  OR2_X1 U519 ( .A1(n549), .A2(n371), .ZN(n426) );
  XNOR2_X2 U520 ( .A(n474), .B(n473), .ZN(n371) );
  NAND2_X1 U521 ( .A1(n706), .A2(n372), .ZN(n710) );
  NAND2_X1 U522 ( .A1(n603), .A2(n376), .ZN(n373) );
  XNOR2_X2 U523 ( .A(n475), .B(G134), .ZN(n515) );
  XNOR2_X2 U524 ( .A(G143), .B(G128), .ZN(n475) );
  OR2_X1 U525 ( .A1(n648), .A2(n385), .ZN(n384) );
  NAND2_X1 U526 ( .A1(n648), .A2(n496), .ZN(n389) );
  XNOR2_X1 U527 ( .A(n631), .B(n392), .ZN(n617) );
  BUF_X1 U528 ( .A(n661), .Z(n394) );
  XNOR2_X1 U529 ( .A(n475), .B(n397), .ZN(n458) );
  INV_X1 U530 ( .A(n427), .ZN(n397) );
  NAND2_X1 U531 ( .A1(n759), .A2(n658), .ZN(n428) );
  XNOR2_X1 U532 ( .A(n431), .B(KEYINPUT32), .ZN(n759) );
  XNOR2_X2 U533 ( .A(n742), .B(n477), .ZN(n494) );
  XNOR2_X1 U534 ( .A(n576), .B(KEYINPUT70), .ZN(n442) );
  INV_X1 U535 ( .A(n761), .ZN(n402) );
  XNOR2_X1 U536 ( .A(n434), .B(n364), .ZN(G60) );
  XNOR2_X1 U537 ( .A(n744), .B(n446), .ZN(n445) );
  INV_X1 U538 ( .A(n570), .ZN(n569) );
  NAND2_X1 U539 ( .A1(n403), .A2(n598), .ZN(n570) );
  INV_X1 U540 ( .A(n586), .ZN(n403) );
  NOR2_X4 U541 ( .A1(n582), .A2(n519), .ZN(n663) );
  INV_X1 U542 ( .A(n617), .ZN(n408) );
  XNOR2_X2 U543 ( .A(n411), .B(G953), .ZN(n537) );
  XNOR2_X1 U544 ( .A(n729), .B(KEYINPUT122), .ZN(n412) );
  INV_X1 U545 ( .A(n631), .ZN(n674) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n427), .B(n452), .ZN(n520) );
  XNOR2_X2 U548 ( .A(G146), .B(G125), .ZN(n427) );
  NAND2_X1 U549 ( .A1(n622), .A2(n623), .ZN(n431) );
  AND2_X1 U550 ( .A1(n432), .A2(n420), .ZN(G54) );
  XNOR2_X1 U551 ( .A(n433), .B(n724), .ZN(n432) );
  NAND2_X1 U552 ( .A1(n728), .A2(G469), .ZN(n433) );
  NAND2_X1 U553 ( .A1(n437), .A2(n589), .ZN(n441) );
  NAND2_X1 U554 ( .A1(n442), .A2(n438), .ZN(n437) );
  INV_X1 U555 ( .A(n588), .ZN(n438) );
  NOR2_X1 U556 ( .A1(n588), .A2(n589), .ZN(n440) );
  NAND2_X1 U557 ( .A1(n441), .A2(n439), .ZN(n443) );
  NAND2_X1 U558 ( .A1(n442), .A2(n440), .ZN(n439) );
  XNOR2_X1 U559 ( .A(n449), .B(n448), .ZN(G51) );
  NAND2_X1 U560 ( .A1(n450), .A2(n420), .ZN(n449) );
  XNOR2_X1 U561 ( .A(n451), .B(n362), .ZN(n450) );
  NOR2_X2 U562 ( .A1(n559), .A2(n583), .ZN(n666) );
  XNOR2_X2 U563 ( .A(n511), .B(n453), .ZN(n583) );
  NOR2_X2 U564 ( .A1(n567), .A2(n611), .ZN(n661) );
  XOR2_X1 U565 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n454) );
  XNOR2_X1 U566 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n455) );
  AND2_X1 U567 ( .A1(n672), .A2(KEYINPUT2), .ZN(n456) );
  XNOR2_X1 U568 ( .A(n581), .B(n580), .ZN(n761) );
  INV_X1 U569 ( .A(KEYINPUT48), .ZN(n589) );
  XNOR2_X1 U570 ( .A(n489), .B(KEYINPUT100), .ZN(n490) );
  INV_X1 U571 ( .A(n563), .ZN(n544) );
  XNOR2_X1 U572 ( .A(n491), .B(n490), .ZN(n492) );
  AND2_X1 U573 ( .A1(n679), .A2(n544), .ZN(n554) );
  INV_X1 U574 ( .A(G472), .ZN(n496) );
  INV_X1 U575 ( .A(n646), .ZN(n647) );
  INV_X1 U576 ( .A(n537), .ZN(n748) );
  XNOR2_X1 U577 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n580) );
  NOR2_X1 U578 ( .A1(n537), .A2(G952), .ZN(n457) );
  NAND2_X1 U579 ( .A1(G224), .A2(n537), .ZN(n459) );
  XNOR2_X1 U580 ( .A(n459), .B(n458), .ZN(n462) );
  INV_X1 U581 ( .A(n462), .ZN(n460) );
  NAND2_X1 U582 ( .A1(n460), .A2(KEYINPUT18), .ZN(n464) );
  INV_X1 U583 ( .A(KEYINPUT18), .ZN(n461) );
  NAND2_X1 U584 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U585 ( .A1(n464), .A2(n463), .ZN(n466) );
  XNOR2_X1 U586 ( .A(n476), .B(KEYINPUT17), .ZN(n465) );
  XNOR2_X1 U587 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U588 ( .A(KEYINPUT16), .B(n514), .Z(n468) );
  XNOR2_X1 U589 ( .A(G110), .B(n499), .ZN(n467) );
  XNOR2_X1 U590 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U591 ( .A(n493), .B(n469), .ZN(n732) );
  XNOR2_X1 U592 ( .A(n470), .B(n732), .ZN(n720) );
  XNOR2_X1 U593 ( .A(G902), .B(KEYINPUT15), .ZN(n640) );
  NAND2_X1 U594 ( .A1(n720), .A2(n640), .ZN(n474) );
  OR2_X1 U595 ( .A1(G237), .A2(G902), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G210), .A2(n545), .ZN(n472) );
  XNOR2_X1 U597 ( .A(KEYINPUT71), .B(G469), .ZN(n485) );
  XOR2_X1 U598 ( .A(G146), .B(n476), .Z(n477) );
  NAND2_X1 U599 ( .A1(G227), .A2(n537), .ZN(n478) );
  XOR2_X1 U600 ( .A(n480), .B(n479), .Z(n481) );
  INV_X1 U601 ( .A(KEYINPUT1), .ZN(n486) );
  NAND2_X1 U602 ( .A1(n504), .A2(G210), .ZN(n488) );
  XOR2_X1 U603 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n487) );
  XNOR2_X1 U604 ( .A(n488), .B(n487), .ZN(n491) );
  XOR2_X1 U605 ( .A(G116), .B(G137), .Z(n489) );
  XNOR2_X1 U606 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n497), .B(n498), .ZN(n509) );
  XNOR2_X1 U608 ( .A(n499), .B(KEYINPUT103), .ZN(n503) );
  XOR2_X1 U609 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n501) );
  XNOR2_X1 U610 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n503), .B(n502), .ZN(n507) );
  NAND2_X1 U612 ( .A1(G214), .A2(n504), .ZN(n505) );
  XNOR2_X1 U613 ( .A(n520), .B(n505), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U615 ( .A(n509), .B(n508), .ZN(n646) );
  XNOR2_X1 U616 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n510) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n513) );
  NAND2_X1 U618 ( .A1(G217), .A2(n527), .ZN(n512) );
  XOR2_X1 U619 ( .A(KEYINPUT7), .B(n514), .Z(n517) );
  XNOR2_X1 U620 ( .A(n515), .B(G122), .ZN(n516) );
  XNOR2_X1 U621 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U622 ( .A(n559), .ZN(n582) );
  INV_X1 U623 ( .A(n520), .ZN(n521) );
  XOR2_X1 U624 ( .A(n522), .B(n521), .Z(n744) );
  XOR2_X1 U625 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n524) );
  XNOR2_X1 U626 ( .A(G128), .B(KEYINPUT96), .ZN(n523) );
  XNOR2_X1 U627 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U628 ( .A(G119), .B(G110), .ZN(n526) );
  NAND2_X1 U629 ( .A1(G221), .A2(n527), .ZN(n528) );
  XOR2_X1 U630 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n531) );
  NAND2_X1 U631 ( .A1(n640), .A2(G234), .ZN(n529) );
  XNOR2_X1 U632 ( .A(n529), .B(KEYINPUT20), .ZN(n541) );
  NAND2_X1 U633 ( .A1(G217), .A2(n541), .ZN(n530) );
  XNOR2_X1 U634 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U635 ( .A1(G234), .A2(G237), .ZN(n534) );
  XNOR2_X1 U636 ( .A(n534), .B(KEYINPUT14), .ZN(n536) );
  NAND2_X1 U637 ( .A1(G952), .A2(n536), .ZN(n703) );
  NOR2_X1 U638 ( .A1(n703), .A2(G953), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n535), .B(KEYINPUT95), .ZN(n595) );
  NAND2_X1 U640 ( .A1(G902), .A2(n536), .ZN(n593) );
  NOR2_X1 U641 ( .A1(G900), .A2(n593), .ZN(n538) );
  NAND2_X1 U642 ( .A1(n538), .A2(n748), .ZN(n539) );
  NAND2_X1 U643 ( .A1(n595), .A2(n539), .ZN(n540) );
  XNOR2_X1 U644 ( .A(n540), .B(KEYINPUT80), .ZN(n543) );
  NAND2_X1 U645 ( .A1(G221), .A2(n541), .ZN(n542) );
  XNOR2_X1 U646 ( .A(KEYINPUT21), .B(n542), .ZN(n678) );
  INV_X1 U647 ( .A(n678), .ZN(n600) );
  NAND2_X1 U648 ( .A1(n543), .A2(n600), .ZN(n563) );
  NAND2_X1 U649 ( .A1(G214), .A2(n545), .ZN(n691) );
  NAND2_X1 U650 ( .A1(n550), .A2(n691), .ZN(n546) );
  NOR2_X1 U651 ( .A1(n675), .A2(n546), .ZN(n547) );
  XOR2_X1 U652 ( .A(KEYINPUT43), .B(n547), .Z(n548) );
  XOR2_X1 U653 ( .A(KEYINPUT108), .B(n548), .Z(n549) );
  NOR2_X1 U654 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U655 ( .A(KEYINPUT36), .B(n552), .ZN(n553) );
  XOR2_X1 U656 ( .A(KEYINPUT90), .B(n604), .Z(n618) );
  NAND2_X1 U657 ( .A1(n553), .A2(n618), .ZN(n671) );
  AND2_X1 U658 ( .A1(n616), .A2(n554), .ZN(n556) );
  XNOR2_X1 U659 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n555) );
  XNOR2_X1 U660 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U661 ( .A1(n557), .A2(n628), .ZN(n586) );
  NOR2_X1 U662 ( .A1(KEYINPUT47), .A2(n695), .ZN(n560) );
  NAND2_X1 U663 ( .A1(n569), .A2(n560), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n671), .A2(n561), .ZN(n575) );
  NAND2_X1 U665 ( .A1(n356), .A2(n628), .ZN(n562) );
  NOR2_X2 U666 ( .A1(n565), .A2(n564), .ZN(n578) );
  XNOR2_X1 U667 ( .A(n566), .B(KEYINPUT109), .ZN(n567) );
  NAND2_X1 U668 ( .A1(n582), .A2(n583), .ZN(n611) );
  NAND2_X1 U669 ( .A1(n695), .A2(KEYINPUT47), .ZN(n568) );
  XNOR2_X1 U670 ( .A(n568), .B(KEYINPUT82), .ZN(n572) );
  NAND2_X1 U671 ( .A1(n570), .A2(KEYINPUT47), .ZN(n571) );
  NAND2_X1 U672 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U673 ( .A(KEYINPUT38), .ZN(n577) );
  NAND2_X1 U674 ( .A1(n690), .A2(n578), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n591), .A2(n663), .ZN(n581) );
  NOR2_X1 U676 ( .A1(n583), .A2(n582), .ZN(n601) );
  INV_X1 U677 ( .A(n601), .ZN(n693) );
  NAND2_X1 U678 ( .A1(n691), .A2(n690), .ZN(n694) );
  XNOR2_X1 U679 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n584) );
  XNOR2_X1 U680 ( .A(n585), .B(n584), .ZN(n714) );
  NOR2_X1 U681 ( .A1(n586), .A2(n714), .ZN(n587) );
  XNOR2_X1 U682 ( .A(n587), .B(KEYINPUT42), .ZN(n758) );
  NAND2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n672) );
  NAND2_X1 U684 ( .A1(n638), .A2(n456), .ZN(n592) );
  INV_X1 U685 ( .A(n593), .ZN(n594) );
  NOR2_X1 U686 ( .A1(G898), .A2(n737), .ZN(n733) );
  NAND2_X1 U687 ( .A1(n594), .A2(n733), .ZN(n596) );
  NAND2_X1 U688 ( .A1(n596), .A2(n595), .ZN(n597) );
  AND2_X1 U689 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U690 ( .A1(n606), .A2(n602), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n604), .A2(n622), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n408), .A2(n615), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n356), .A2(n605), .ZN(n651) );
  INV_X1 U694 ( .A(n606), .ZN(n630) );
  NOR2_X1 U695 ( .A1(n678), .A2(n679), .ZN(n676) );
  XNOR2_X2 U696 ( .A(n608), .B(n607), .ZN(n713) );
  NOR2_X1 U697 ( .A1(n630), .A2(n713), .ZN(n610) );
  XNOR2_X1 U698 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n609) );
  XNOR2_X1 U699 ( .A(n610), .B(n609), .ZN(n612) );
  NOR2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U701 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n613) );
  XNOR2_X1 U702 ( .A(n614), .B(n613), .ZN(n756) );
  NOR2_X1 U703 ( .A1(n756), .A2(KEYINPUT67), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT78), .ZN(n623) );
  AND2_X1 U706 ( .A1(n756), .A2(KEYINPUT67), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n636) );
  AND2_X1 U708 ( .A1(n631), .A2(n676), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n653) );
  XOR2_X1 U711 ( .A(KEYINPUT101), .B(KEYINPUT31), .Z(n634) );
  NOR2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n686) );
  NAND2_X1 U713 ( .A1(n686), .A2(n606), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n634), .B(n633), .ZN(n667) );
  NOR2_X1 U715 ( .A1(n653), .A2(n667), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n638), .A2(n672), .ZN(n707) );
  NAND2_X1 U717 ( .A1(n639), .A2(n704), .ZN(n644) );
  INV_X1 U718 ( .A(n640), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT65), .B(n642), .Z(n643) );
  XNOR2_X1 U721 ( .A(KEYINPUT63), .B(KEYINPUT91), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(G57) );
  XNOR2_X1 U723 ( .A(G101), .B(n651), .ZN(G3) );
  NAND2_X1 U724 ( .A1(n653), .A2(n663), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(G104), .ZN(G6) );
  XNOR2_X1 U726 ( .A(G107), .B(KEYINPUT114), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n655) );
  NAND2_X1 U728 ( .A1(n653), .A2(n666), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(G9) );
  XNOR2_X1 U731 ( .A(n658), .B(G110), .ZN(G12) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n660) );
  NAND2_X1 U733 ( .A1(n569), .A2(n666), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(G30) );
  XOR2_X1 U735 ( .A(n394), .B(G143), .Z(G45) );
  NAND2_X1 U736 ( .A1(n569), .A2(n663), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n662), .B(G146), .ZN(G48) );
  XOR2_X1 U738 ( .A(G113), .B(KEYINPUT115), .Z(n665) );
  NAND2_X1 U739 ( .A1(n667), .A2(n663), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n668), .B(KEYINPUT116), .ZN(n669) );
  XNOR2_X1 U743 ( .A(G116), .B(n669), .ZN(G18) );
  XOR2_X1 U744 ( .A(G125), .B(KEYINPUT37), .Z(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(G27) );
  XNOR2_X1 U746 ( .A(G134), .B(n672), .ZN(G36) );
  XOR2_X1 U747 ( .A(G140), .B(n673), .Z(G42) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U749 ( .A(KEYINPUT50), .B(n677), .Z(n683) );
  NAND2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT49), .ZN(n681) );
  XNOR2_X1 U752 ( .A(KEYINPUT117), .B(n681), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n674), .A2(n684), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U756 ( .A(n687), .B(KEYINPUT118), .Z(n688) );
  XNOR2_X1 U757 ( .A(KEYINPUT51), .B(n688), .ZN(n689) );
  NOR2_X1 U758 ( .A1(n714), .A2(n689), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U763 ( .A1(n698), .A2(n713), .ZN(n699) );
  NOR2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U765 ( .A(n701), .B(KEYINPUT52), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n704), .A2(KEYINPUT2), .ZN(n705) );
  XNOR2_X1 U768 ( .A(n705), .B(KEYINPUT83), .ZN(n706) );
  INV_X1 U769 ( .A(n745), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n708), .A2(KEYINPUT2), .ZN(n709) );
  NOR2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U774 ( .A(n715), .B(KEYINPUT119), .ZN(n716) );
  XNOR2_X1 U775 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n718) );
  XNOR2_X1 U776 ( .A(n719), .B(n718), .ZN(G75) );
  XOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n723) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT121), .ZN(n722) );
  XNOR2_X1 U779 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U780 ( .A1(G478), .A2(n728), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U782 ( .A1(n731), .A2(n727), .ZN(G63) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(G66) );
  XNOR2_X1 U784 ( .A(n732), .B(G101), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n741) );
  NAND2_X1 U786 ( .A1(G953), .A2(G224), .ZN(n735) );
  XNOR2_X1 U787 ( .A(KEYINPUT61), .B(n735), .ZN(n736) );
  NAND2_X1 U788 ( .A1(n736), .A2(G898), .ZN(n739) );
  NAND2_X1 U789 ( .A1(n704), .A2(n737), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(G69) );
  XOR2_X1 U792 ( .A(n742), .B(KEYINPUT4), .Z(n743) );
  XOR2_X1 U793 ( .A(n744), .B(n743), .Z(n750) );
  INV_X1 U794 ( .A(n750), .ZN(n746) );
  XOR2_X1 U795 ( .A(n746), .B(n745), .Z(n747) );
  NOR2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U797 ( .A(KEYINPUT123), .B(n749), .ZN(n755) );
  XOR2_X1 U798 ( .A(G227), .B(n750), .Z(n751) );
  NAND2_X1 U799 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U800 ( .A1(G953), .A2(n752), .ZN(n753) );
  XNOR2_X1 U801 ( .A(KEYINPUT124), .B(n753), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U803 ( .A(n756), .B(G122), .Z(G24) );
  XOR2_X1 U804 ( .A(G137), .B(KEYINPUT126), .Z(n757) );
  XNOR2_X1 U805 ( .A(n758), .B(n757), .ZN(G39) );
  XOR2_X1 U806 ( .A(G119), .B(n759), .Z(n760) );
  XNOR2_X1 U807 ( .A(KEYINPUT125), .B(n760), .ZN(G21) );
  XNOR2_X1 U808 ( .A(G131), .B(KEYINPUT127), .ZN(n762) );
  XNOR2_X1 U809 ( .A(n762), .B(n761), .ZN(G33) );
endmodule

