//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n201), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n209), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n214), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G68), .A2(G77), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n203), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT65), .ZN(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n216), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n227), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n256), .B1(new_n208), .B2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n254), .B1(new_n258), .B2(new_n216), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G58), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n209), .A2(G33), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n216), .A2(new_n263), .A3(new_n201), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n259), .B1(new_n271), .B2(new_n256), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n285), .C2(new_n276), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n282), .A2(G274), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G222), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G223), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n294), .B1(new_n202), .B2(new_n292), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n288), .B1(new_n297), .B2(new_n275), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n298), .A2(G190), .B1(KEYINPUT70), .B2(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n274), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n303), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n274), .A2(new_n305), .A3(new_n300), .A4(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n255), .A2(new_n227), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n267), .B2(new_n270), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(G169), .B2(new_n298), .C1(new_n310), .C2(new_n259), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G107), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n292), .A2(new_n293), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n315), .B1(new_n295), .B2(new_n218), .C1(new_n233), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n275), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n279), .A2(G244), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n319), .A2(new_n287), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G200), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G20), .A2(G77), .ZN(new_n323));
  INV_X1    g0123(.A(new_n269), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n323), .B1(new_n260), .B2(new_n324), .C1(new_n266), .C2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n326), .A2(new_n256), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n253), .A2(new_n202), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n258), .B2(new_n202), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n322), .B(new_n330), .C1(new_n331), .C2(new_n321), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n321), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n318), .A2(new_n307), .A3(new_n320), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n304), .A2(new_n306), .A3(new_n311), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n257), .A2(G68), .ZN(new_n339));
  XOR2_X1   g0139(.A(new_n339), .B(KEYINPUT71), .Z(new_n340));
  OAI22_X1  g0140(.A1(new_n324), .A2(new_n216), .B1(new_n209), .B2(G68), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n266), .A2(new_n202), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n256), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT11), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT72), .B1(new_n252), .B2(G68), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n347), .B(KEYINPUT12), .Z(new_n348));
  AND4_X1   g0148(.A1(new_n340), .A2(new_n345), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n292), .A2(G232), .A3(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n351), .C1(new_n316), .C2(new_n217), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n275), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n279), .A2(G238), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(new_n287), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n353), .B2(new_n355), .ZN(new_n358));
  OAI21_X1  g0158(.A(G169), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n355), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(G179), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT73), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n349), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G200), .B1(new_n357), .B2(new_n358), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(G190), .A3(new_n364), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n349), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n338), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(G58), .B(G68), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n291), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n314), .A2(KEYINPUT74), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n290), .A2(new_n209), .A3(new_n291), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n385), .A2(KEYINPUT75), .A3(G68), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT75), .B1(new_n385), .B2(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n377), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n201), .B1(new_n384), .B2(new_n378), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n376), .B1(new_n389), .B2(new_n375), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n390), .A3(new_n256), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n265), .A2(new_n257), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n252), .B2(new_n265), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(KEYINPUT76), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n286), .A2(G232), .A3(new_n283), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n287), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n217), .A2(G1698), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n401), .B1(G223), .B2(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n286), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n333), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n400), .A2(new_n404), .A3(G179), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT77), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n407), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT77), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n405), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n397), .A2(new_n398), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT18), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n397), .A2(new_n415), .A3(new_n398), .A4(new_n412), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n400), .A2(new_n404), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n331), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G200), .B2(new_n417), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n391), .A2(new_n394), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT17), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n414), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n372), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n209), .B(G87), .C1(new_n312), .C2(new_n313), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT22), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT23), .ZN(new_n429));
  INV_X1    g0229(.A(G107), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(G20), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT83), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n428), .A2(new_n431), .A3(new_n432), .A4(KEYINPUT83), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT24), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n427), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n427), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n256), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n208), .A2(G33), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n309), .A2(new_n252), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT25), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n252), .A2(new_n444), .A3(G107), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n252), .B2(G107), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n443), .A2(G107), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G257), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n450));
  OAI211_X1 g0250(.A(G250), .B(new_n293), .C1(new_n312), .C2(new_n313), .ZN(new_n451));
  INV_X1    g0251(.A(G294), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n450), .B(new_n451), .C1(new_n285), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n275), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n277), .A2(G1), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n286), .A3(G274), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n275), .B1(new_n456), .B2(new_n455), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G264), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G179), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n453), .A2(new_n275), .B1(new_n458), .B2(G264), .ZN(new_n462));
  AOI21_X1  g0262(.A(G169), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT85), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n466), .A3(new_n299), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n331), .A3(new_n457), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n460), .B2(new_n299), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n449), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT84), .B1(new_n449), .B2(new_n464), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n465), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT80), .ZN(new_n475));
  INV_X1    g0275(.A(G274), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n208), .A2(new_n476), .A3(G45), .ZN(new_n477));
  INV_X1    g0277(.A(G250), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n277), .B2(G1), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n286), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G238), .B(new_n293), .C1(new_n312), .C2(new_n313), .ZN(new_n481));
  OAI211_X1 g0281(.A(G244), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n484), .B2(new_n275), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n333), .ZN(new_n486));
  AOI211_X1 g0286(.A(new_n307), .B(new_n480), .C1(new_n484), .C2(new_n275), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(G179), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(KEYINPUT80), .C1(new_n333), .C2(new_n485), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n292), .A2(new_n209), .A3(G68), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n209), .B1(new_n351), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(G87), .B2(new_n206), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n266), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n256), .B1(new_n253), .B2(new_n325), .ZN(new_n498));
  INV_X1    g0298(.A(new_n325), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n443), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n488), .A2(new_n490), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n485), .A2(G190), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(new_n256), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n325), .A2(new_n253), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n443), .A2(G87), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n485), .A2(new_n299), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT81), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n292), .A2(G244), .A3(new_n293), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT79), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(KEYINPUT4), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n516), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n292), .A2(new_n518), .A3(G244), .A4(new_n293), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n275), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n455), .A2(new_n456), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G257), .A3(new_n286), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n457), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n523), .A2(G179), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n522), .B2(new_n275), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n333), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  AND2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(new_n205), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n430), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n535), .A2(new_n209), .B1(new_n202), .B2(new_n324), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n430), .B1(new_n384), .B2(new_n378), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n256), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n252), .A2(G97), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n443), .B2(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n523), .A2(new_n527), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n384), .A2(new_n378), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G107), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n533), .A2(new_n534), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n309), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n540), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT78), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n538), .A2(new_n552), .A3(new_n540), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n529), .A2(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n544), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n512), .A2(new_n513), .A3(new_n542), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n542), .A2(new_n555), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT81), .B1(new_n557), .B2(new_n511), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n443), .A2(G116), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n253), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n255), .A2(new_n227), .B1(G20), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n521), .B(new_n209), .C1(G33), .C2(new_n495), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT20), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n563), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n559), .B(new_n561), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n524), .A2(G270), .A3(new_n286), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n568), .A2(new_n457), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n292), .A2(G264), .A3(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n292), .A2(G257), .A3(new_n293), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n314), .A2(G303), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n275), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(new_n574), .A3(G179), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n567), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n566), .B1(new_n575), .B2(G200), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n331), .B2(new_n575), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n575), .A2(new_n566), .A3(G169), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n579), .B(new_n581), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n474), .A2(new_n556), .A3(new_n558), .A4(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n425), .A2(new_n589), .ZN(G372));
  OAI21_X1  g0390(.A(KEYINPUT86), .B1(new_n486), .B2(new_n487), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT86), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n489), .B(new_n592), .C1(new_n333), .C2(new_n485), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n509), .B1(new_n594), .B2(new_n501), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n441), .B(new_n448), .C1(new_n469), .C2(new_n470), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n542), .A3(new_n596), .A4(new_n555), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n449), .A2(new_n464), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n579), .B1(new_n585), .B2(new_n586), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT26), .B1(new_n511), .B2(new_n542), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n543), .A2(G169), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n604), .A2(new_n528), .B1(new_n551), .B2(new_n553), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n595), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n501), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n591), .B2(new_n593), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n602), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n424), .B1(new_n601), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n395), .A2(new_n412), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(new_n415), .ZN(new_n613));
  INV_X1    g0413(.A(new_n336), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n370), .B1(new_n367), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n421), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n304), .A2(new_n306), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(new_n311), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n620), .ZN(G369));
  NAND3_X1  g0421(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G213), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT87), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(G343), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(G343), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n567), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n599), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n587), .B2(new_n632), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G330), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n631), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n449), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n474), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n598), .B2(new_n631), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n449), .A2(new_n464), .A3(new_n631), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n599), .A2(new_n631), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n474), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(G399));
  INV_X1    g0446(.A(new_n212), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G41), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G1), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n226), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT28), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n602), .A2(new_n606), .A3(new_n609), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n598), .B(new_n579), .C1(new_n586), .C2(new_n585), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n542), .A2(new_n555), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n596), .A4(new_n595), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n637), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT88), .B1(new_n659), .B2(KEYINPUT29), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n631), .B1(new_n601), .B2(new_n610), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n465), .A2(new_n473), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n597), .B1(new_n666), .B2(new_n600), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n604), .A2(new_n528), .B1(new_n538), .B2(new_n540), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(new_n603), .A3(new_n510), .A4(new_n502), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n551), .A2(new_n553), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n530), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n671), .A2(new_n509), .A3(new_n608), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n609), .B(new_n669), .C1(new_n672), .C2(new_n603), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT29), .B(new_n631), .C1(new_n667), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT89), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n595), .A2(new_n605), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n608), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n599), .A2(new_n465), .A3(new_n473), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n677), .B(new_n669), .C1(new_n678), .C2(new_n597), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT89), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT29), .A4(new_n631), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n462), .A2(new_n569), .A3(new_n574), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n529), .A3(new_n487), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n529), .A4(new_n487), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n485), .A2(G179), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n543), .A2(new_n460), .A3(new_n575), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n637), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n693), .B(new_n694), .C1(new_n589), .C2(new_n637), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n665), .A2(new_n682), .B1(G330), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n654), .B1(new_n696), .B2(G1), .ZN(G364));
  AND2_X1   g0497(.A1(new_n209), .A2(G13), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n208), .B1(new_n698), .B2(G45), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n648), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n636), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(G330), .B2(new_n634), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n212), .A2(new_n292), .ZN(new_n704));
  INV_X1    g0504(.A(G355), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(G116), .B2(new_n212), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n250), .A2(G45), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n647), .A2(new_n292), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n226), .B2(new_n277), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n706), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n227), .B1(G20), .B2(new_n333), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n701), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n209), .A2(new_n331), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n307), .A2(G200), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n209), .A2(G190), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(new_n720), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n722), .A2(new_n263), .B1(new_n725), .B2(new_n202), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT32), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G159), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n730), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT32), .A3(G159), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n726), .A2(new_n727), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n299), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT91), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT91), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G87), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n735), .B(new_n742), .C1(new_n727), .C2(new_n726), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n723), .A2(new_n736), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n209), .A2(new_n307), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n292), .B1(new_n744), .B2(new_n430), .C1(new_n746), .C2(new_n216), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n331), .A3(G200), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n209), .B1(new_n729), .B2(G190), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n201), .B1(new_n749), .B2(new_n495), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n743), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n753));
  INV_X1    g0553(.A(G322), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT33), .B(G317), .Z(new_n755));
  OAI22_X1  g0555(.A1(new_n722), .A2(new_n754), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT93), .Z(new_n757));
  AOI22_X1  g0557(.A1(G329), .A2(new_n733), .B1(new_n724), .B2(G311), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n314), .C1(new_n759), .C2(new_n744), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n746), .A2(new_n761), .B1(new_n749), .B2(new_n452), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G303), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n757), .B(new_n763), .C1(new_n764), .C2(new_n740), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n753), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n718), .B1(new_n767), .B2(new_n715), .ZN(new_n768));
  INV_X1    g0568(.A(new_n714), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n634), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n703), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  INV_X1    g0572(.A(new_n744), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G87), .A2(new_n773), .B1(new_n733), .B2(G311), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n774), .B(new_n314), .C1(new_n452), .C2(new_n722), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n746), .A2(new_n764), .B1(new_n749), .B2(new_n495), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n748), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G283), .B1(new_n724), .B2(G116), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n777), .B(new_n780), .C1(new_n430), .C2(new_n740), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G143), .A2(new_n721), .B1(new_n724), .B2(G159), .ZN(new_n782));
  INV_X1    g0582(.A(G137), .ZN(new_n783));
  INV_X1    g0583(.A(G150), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n782), .B1(new_n783), .B2(new_n746), .C1(new_n784), .C2(new_n748), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT34), .Z(new_n786));
  OAI21_X1  g0586(.A(new_n292), .B1(new_n744), .B2(new_n201), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G132), .B2(new_n733), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n788), .B1(new_n263), .B2(new_n749), .C1(new_n216), .C2(new_n740), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n781), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n791));
  INV_X1    g0591(.A(new_n715), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n790), .B2(KEYINPUT95), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n701), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n715), .A2(new_n712), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n202), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n637), .B1(new_n327), .B2(new_n329), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n614), .B1(new_n332), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n614), .A2(new_n631), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n798), .B1(new_n712), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n803), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n659), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n661), .A2(new_n803), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n695), .A2(G330), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n701), .B1(new_n811), .B2(KEYINPUT96), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(KEYINPUT96), .B2(new_n811), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT97), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n809), .A2(new_n810), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT98), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n813), .B2(new_n814), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n805), .B1(new_n815), .B2(new_n818), .ZN(G384));
  NAND2_X1  g0619(.A1(new_n385), .A2(G68), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT75), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n385), .A2(KEYINPUT75), .A3(G68), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n309), .B1(new_n824), .B2(new_n377), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n374), .B1(new_n386), .B2(new_n387), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n376), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n393), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n420), .B1(new_n828), .B2(new_n625), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n408), .A2(new_n411), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT37), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n829), .C2(new_n831), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n397), .A2(new_n398), .A3(new_n626), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n413), .A2(new_n836), .A3(new_n837), .A4(new_n420), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n828), .A2(new_n625), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n422), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n839), .A2(new_n841), .A3(KEYINPUT38), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT38), .B1(new_n839), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n807), .A2(new_n801), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n361), .A2(new_n366), .ZN(new_n846));
  INV_X1    g0646(.A(new_n349), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n637), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n370), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n847), .B(new_n637), .C1(new_n846), .C2(new_n371), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n844), .A2(new_n853), .B1(new_n613), .B2(new_n626), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n842), .A2(new_n843), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n413), .A2(new_n837), .A3(new_n420), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n830), .B1(new_n391), .B2(new_n394), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n391), .A2(new_n394), .A3(new_n419), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT102), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n612), .A2(new_n862), .A3(new_n420), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n836), .A3(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n858), .A2(new_n836), .B1(new_n864), .B2(KEYINPUT37), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n836), .B1(new_n613), .B2(new_n421), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n857), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n839), .A2(new_n841), .A3(KEYINPUT38), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT39), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n856), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n848), .A2(new_n637), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n854), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n665), .A2(new_n682), .A3(new_n424), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n620), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n872), .B(new_n874), .Z(new_n875));
  XNOR2_X1  g0675(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n691), .B2(new_n692), .ZN(new_n878));
  AOI211_X1 g0678(.A(KEYINPUT104), .B(KEYINPUT31), .C1(new_n690), .C2(new_n637), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n880), .B(new_n694), .C1(new_n589), .C2(new_n637), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n803), .B1(new_n850), .B2(new_n851), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n876), .B1(new_n844), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n881), .A2(new_n882), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n838), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n613), .A2(new_n421), .ZN(new_n888));
  INV_X1    g0688(.A(new_n836), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n885), .B(KEYINPUT40), .C1(new_n842), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n424), .A2(new_n881), .ZN(new_n894));
  OAI21_X1  g0694(.A(G330), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n875), .A2(new_n896), .B1(new_n208), .B2(new_n698), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n875), .B2(new_n896), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(G116), .A3(new_n228), .A4(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT36), .Z(new_n902));
  AOI211_X1 g0702(.A(new_n202), .B(new_n652), .C1(G58), .C2(G68), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n904), .A2(KEYINPUT99), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n216), .A2(G68), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT100), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n904), .B2(KEYINPUT99), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n208), .B(G13), .C1(new_n905), .C2(new_n908), .ZN(new_n909));
  OR3_X1    g0709(.A1(new_n898), .A2(new_n902), .A3(new_n909), .ZN(G367));
  INV_X1    g0710(.A(new_n670), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n657), .B1(new_n911), .B2(new_n631), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n605), .A2(new_n637), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n474), .A3(new_n644), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT42), .Z(new_n916));
  AOI21_X1  g0716(.A(new_n666), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n631), .B1(new_n917), .B2(new_n668), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n637), .A2(new_n507), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n595), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n609), .B2(new_n920), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT43), .B1(new_n922), .B2(KEYINPUT105), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT105), .B2(new_n922), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n919), .B2(new_n925), .ZN(new_n927));
  INV_X1    g0727(.A(new_n641), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n914), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n927), .B(new_n929), .Z(new_n930));
  XOR2_X1   g0730(.A(new_n648), .B(KEYINPUT41), .Z(new_n931));
  INV_X1    g0731(.A(KEYINPUT44), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n914), .B1(KEYINPUT106), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n645), .A2(new_n642), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n933), .B(new_n934), .C1(KEYINPUT106), .C2(new_n932), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n645), .A2(new_n914), .A3(new_n642), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT45), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n641), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n928), .B1(new_n939), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n645), .B1(new_n640), .B2(new_n644), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n636), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n696), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT107), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT107), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(new_n951), .A3(new_n943), .A4(new_n944), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n931), .B1(new_n953), .B2(new_n696), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n930), .B1(new_n954), .B2(new_n700), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n716), .B1(new_n212), .B2(new_n325), .C1(new_n709), .C2(new_n239), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n956), .A2(new_n701), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n773), .A2(G77), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n725), .B2(new_n216), .C1(new_n784), .C2(new_n722), .ZN(new_n959));
  INV_X1    g0759(.A(new_n746), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n778), .A2(G159), .B1(new_n960), .B2(G143), .ZN(new_n961));
  INV_X1    g0761(.A(new_n749), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(G68), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n314), .B1(new_n733), .B2(G137), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n959), .B(new_n965), .C1(G58), .C2(new_n741), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT108), .ZN(new_n967));
  INV_X1    g0767(.A(G311), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n748), .A2(new_n452), .B1(new_n746), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n314), .B1(new_n722), .B2(new_n764), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(G107), .C2(new_n962), .ZN(new_n971));
  INV_X1    g0771(.A(G317), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n744), .A2(new_n495), .B1(new_n730), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G283), .B2(new_n724), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n740), .B2(new_n560), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n741), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n971), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n967), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  OAI221_X1 g0780(.A(new_n957), .B1(new_n769), .B2(new_n922), .C1(new_n980), .C2(new_n792), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n955), .A2(new_n981), .ZN(G387));
  XNOR2_X1  g0782(.A(new_n648), .B(KEYINPUT114), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n950), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n696), .B2(new_n947), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n640), .A2(new_n769), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G317), .A2(new_n721), .B1(new_n724), .B2(G303), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n968), .B2(new_n748), .C1(new_n754), .C2(new_n746), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n740), .A2(new_n452), .B1(new_n759), .B2(new_n749), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT112), .Z(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(KEYINPUT49), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(KEYINPUT49), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n314), .B1(new_n730), .B2(new_n761), .C1(new_n560), .C2(new_n744), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G150), .A2(new_n733), .B1(new_n724), .B2(G68), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n216), .B2(new_n722), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n740), .A2(new_n202), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n265), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1001), .C1(new_n1002), .C2(new_n778), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n749), .A2(new_n325), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n292), .B1(new_n744), .B2(new_n495), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(G159), .C2(new_n960), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n792), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n704), .A2(new_n650), .B1(G107), .B2(new_n212), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n260), .A2(G50), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT50), .Z(new_n1011));
  NAND3_X1  g0811(.A1(new_n650), .A2(new_n277), .A3(new_n246), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n708), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT109), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1013), .A2(new_n1014), .B1(G45), .B2(new_n236), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n701), .B1(new_n1017), .B2(new_n717), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT110), .Z(new_n1019));
  OR2_X1    g0819(.A1(new_n1008), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT113), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n987), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1008), .A2(new_n1021), .A3(new_n1019), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1022), .A2(new_n1023), .B1(new_n700), .B2(new_n947), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n986), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT115), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n986), .A2(KEYINPUT115), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(G393));
  NAND3_X1  g0829(.A1(new_n943), .A2(KEYINPUT116), .A3(new_n944), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT116), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n942), .A2(new_n1031), .A3(new_n641), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n700), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n244), .A2(new_n708), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n716), .B1(new_n495), .B2(new_n212), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n701), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n960), .A2(G150), .B1(new_n721), .B2(G159), .ZN(new_n1038));
  XOR2_X1   g0838(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n741), .A2(G68), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n314), .B1(new_n773), .B2(G87), .ZN(new_n1042));
  INV_X1    g0842(.A(G143), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n725), .A2(new_n260), .B1(new_n730), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n749), .A2(new_n202), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G50), .B2(new_n778), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n741), .A2(G283), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n292), .B1(new_n773), .B2(G107), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G322), .A2(new_n733), .B1(new_n724), .B2(G294), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n778), .A2(G303), .B1(new_n962), .B2(G116), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n960), .A2(G317), .B1(new_n721), .B2(G311), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1040), .A2(new_n1048), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1037), .B1(new_n715), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n914), .B2(new_n769), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1033), .A2(new_n950), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1060), .A2(new_n984), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1061), .B2(new_n953), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(new_n796), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n701), .B1(new_n1002), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n722), .A2(new_n560), .B1(new_n730), .B2(new_n452), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G97), .B2(new_n724), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n292), .B(new_n1046), .C1(G68), .C2(new_n773), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n778), .A2(G107), .B1(new_n960), .B2(G283), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1067), .A2(new_n742), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n741), .A2(G150), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT53), .ZN(new_n1072));
  INV_X1    g0872(.A(G125), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n744), .A2(new_n216), .B1(new_n730), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n314), .B(new_n1074), .C1(G132), .C2(new_n721), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT54), .B(G143), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n778), .A2(G137), .B1(new_n724), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT121), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n960), .A2(G128), .B1(new_n962), .B2(G159), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1075), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1070), .B1(new_n1072), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1065), .B1(new_n1084), .B2(new_n715), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n870), .B2(new_n713), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n881), .A2(new_n882), .A3(G330), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n871), .B1(new_n845), .B2(new_n852), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n855), .B1(new_n842), .B2(new_n891), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n839), .A2(new_n841), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n857), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1089), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n871), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n631), .B1(new_n667), .B2(new_n673), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n800), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n802), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n852), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n842), .A2(new_n891), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1088), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n853), .A2(new_n1095), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n856), .B2(new_n869), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1095), .B1(new_n842), .B2(new_n891), .C1(new_n1099), .C2(new_n1098), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n695), .A2(G330), .A3(new_n852), .A4(new_n806), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1086), .B1(new_n1109), .B2(new_n699), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n424), .A2(G330), .A3(new_n881), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n873), .A2(new_n620), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n695), .A2(G330), .A3(new_n806), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1114), .A2(new_n1099), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n845), .B1(new_n1115), .B2(new_n1088), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n881), .A2(G330), .A3(new_n806), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1098), .B(new_n1107), .C1(new_n1117), .C2(new_n852), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1109), .B2(KEYINPUT120), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(KEYINPUT120), .B2(new_n1109), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1103), .A2(new_n1108), .A3(new_n1119), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1103), .A2(new_n1108), .A3(new_n1119), .A4(KEYINPUT118), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n984), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT119), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(KEYINPUT119), .B(new_n984), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1111), .B1(new_n1128), .B2(new_n1129), .ZN(G378));
  NAND2_X1  g0930(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1113), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT122), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n618), .A2(new_n311), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n272), .A2(new_n625), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1138), .B(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n884), .A3(G330), .A4(new_n892), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n883), .B1(new_n1092), .B2(new_n868), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n876), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n892), .B(G330), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1141), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n872), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n872), .A3(new_n1142), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1135), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1133), .A2(new_n1134), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1113), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1147), .A2(new_n872), .A3(new_n1142), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n1148), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1135), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1148), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT122), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1152), .A2(new_n1156), .A3(new_n1158), .A4(new_n983), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n721), .A2(G128), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n725), .B2(new_n783), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G150), .B2(new_n962), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n778), .A2(G132), .B1(new_n960), .B2(G125), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n740), .C2(new_n1076), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n773), .A2(G159), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n733), .C2(G124), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n778), .A2(G97), .B1(new_n960), .B2(G116), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n292), .A2(G41), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n744), .A2(new_n263), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n1175), .A3(new_n963), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n724), .A2(new_n499), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n759), .B2(new_n730), .C1(new_n722), .C2(new_n430), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1176), .A2(new_n1001), .A3(new_n1178), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1173), .B(new_n216), .C1(G33), .C2(G41), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n715), .B1(new_n1170), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n701), .C1(G50), .C2(new_n1064), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1146), .B2(new_n712), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1155), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n700), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1159), .A2(new_n1188), .ZN(G375));
  INV_X1    g0989(.A(new_n1119), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n931), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1116), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n699), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1099), .A2(new_n712), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n701), .B1(G68), .B2(new_n1064), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n722), .A2(new_n783), .B1(new_n725), .B2(new_n784), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G128), .B2(new_n733), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n314), .B(new_n1174), .C1(new_n778), .C2(new_n1077), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n960), .A2(G132), .B1(new_n962), .B2(G50), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n741), .A2(G159), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n958), .A2(new_n314), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT124), .Z(new_n1204));
  NOR2_X1   g1004(.A1(new_n730), .A2(new_n764), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1205), .B(new_n1004), .C1(G283), .C2(new_n721), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n495), .C2(new_n740), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n778), .A2(G116), .B1(new_n724), .B2(G107), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n452), .B2(new_n746), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT123), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1202), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1196), .B1(new_n1211), .B2(new_n715), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1194), .B1(new_n1195), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1193), .A2(new_n1213), .ZN(G381));
  NOR2_X1   g1014(.A1(G375), .A2(G378), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n955), .A2(new_n981), .A3(new_n1062), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1027), .A2(new_n771), .A3(new_n1028), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1218), .A2(G384), .A3(G381), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1215), .A2(new_n1217), .A3(new_n1219), .ZN(G407));
  NAND3_X1  g1020(.A1(new_n628), .A2(new_n629), .A3(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1215), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(G213), .A3(new_n1223), .ZN(G409));
  NAND2_X1  g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1062), .B1(new_n955), .B2(new_n981), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1218), .B(new_n1225), .C1(new_n1217), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1226), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1218), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1216), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1159), .A2(G378), .A3(new_n1188), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1129), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1121), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1133), .A2(new_n1191), .A3(new_n1187), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1188), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1237), .A3(new_n1111), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1232), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1192), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT60), .B1(new_n1192), .B2(new_n1241), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n983), .B(new_n1190), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1213), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n805), .C1(new_n815), .C2(new_n818), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(G384), .A3(new_n1213), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1239), .A2(new_n1240), .A3(new_n1221), .A4(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1222), .B1(new_n1232), .B2(new_n1238), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(G2897), .A3(new_n1222), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1222), .A2(G2897), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(new_n1249), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1252), .B(new_n1253), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1222), .B(new_n1250), .C1(new_n1232), .C2(new_n1238), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(new_n1240), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1231), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1227), .A2(new_n1230), .A3(new_n1253), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1260), .B2(KEYINPUT63), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1254), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1250), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1258), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1254), .A2(new_n1258), .A3(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1264), .B(new_n1267), .C1(new_n1269), .C2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1262), .A2(new_n1272), .ZN(G405));
  INV_X1    g1073(.A(new_n1232), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G378), .B1(new_n1159), .B2(new_n1188), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1251), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1232), .A3(new_n1250), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1278), .A3(new_n1231), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT127), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1276), .A2(new_n1278), .A3(new_n1283), .A4(new_n1231), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1284), .ZN(G402));
endmodule


