//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  INV_X1    g005(.A(G110), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n190), .A2(new_n191), .A3(new_n192), .A4(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(new_n195), .A2(KEYINPUT73), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n188), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(KEYINPUT73), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT72), .A2(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT72), .A3(G125), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT16), .B1(new_n207), .B2(G125), .ZN(new_n210));
  OAI21_X1  g024(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G125), .B(G140), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n196), .A2(KEYINPUT74), .A3(new_n199), .A4(new_n200), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n203), .A2(new_n211), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OR3_X1    g030(.A1(new_n209), .A2(G146), .A3(new_n210), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n190), .A2(new_n194), .A3(new_n191), .ZN(new_n219));
  OAI221_X1 g033(.A(new_n218), .B1(new_n192), .B2(new_n219), .C1(new_n197), .C2(new_n198), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n220), .A3(new_n225), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT25), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G234), .B2(new_n228), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n227), .A2(new_n234), .A3(new_n228), .A4(new_n229), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n227), .A2(new_n229), .ZN(new_n237));
  INV_X1    g051(.A(new_n233), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n228), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT68), .B(G116), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT69), .B1(new_n241), .B2(new_n193), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n193), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n244), .B(G119), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n249), .B2(new_n250), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n213), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT64), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n256), .B1(new_n261), .B2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n260), .A3(new_n213), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n257), .A2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(G134), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT65), .A3(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT11), .B1(new_n273), .B2(G134), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n275), .A2(G137), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT11), .ZN(new_n281));
  AND4_X1   g095(.A1(new_n271), .A2(new_n277), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n273), .A2(KEYINPUT11), .A3(G134), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n278), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n271), .B1(new_n284), .B2(new_n277), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n265), .B(new_n270), .C1(new_n282), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n266), .A2(new_n267), .B1(new_n287), .B2(G128), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G128), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT64), .B(G143), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n255), .B(new_n291), .C1(new_n292), .C2(new_n213), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n261), .A2(G146), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n255), .A4(new_n291), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n288), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n271), .A3(new_n277), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n273), .A2(G134), .ZN(new_n300));
  OAI21_X1  g114(.A(G131), .B1(new_n280), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n286), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT30), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n286), .B(new_n305), .C1(new_n298), .C2(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n254), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n249), .A2(new_n250), .ZN(new_n308));
  INV_X1    g122(.A(new_n251), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G237), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G210), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(G101), .Z(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n307), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n322));
  INV_X1    g136(.A(new_n288), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n296), .B1(new_n262), .B2(new_n291), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n213), .B1(new_n258), .B2(new_n260), .ZN(new_n325));
  NOR4_X1   g139(.A1(new_n325), .A2(KEYINPUT66), .A3(new_n256), .A4(new_n290), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n302), .ZN(new_n328));
  INV_X1    g142(.A(new_n285), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n299), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n331), .A2(new_n269), .B1(new_n262), .B2(new_n264), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n327), .A2(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n254), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n303), .A2(new_n312), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n313), .A2(KEYINPUT28), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n318), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n319), .A2(new_n339), .A3(new_n320), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n327), .A2(new_n328), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n305), .B1(new_n341), .B2(new_n286), .ZN(new_n342));
  INV_X1    g156(.A(new_n306), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n312), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n318), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n334), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT70), .B1(new_n346), .B2(KEYINPUT31), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n321), .B(new_n338), .C1(new_n340), .C2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT71), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT32), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G472), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n336), .A2(new_n337), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n356), .B2(new_n345), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n344), .A2(new_n334), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n318), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(KEYINPUT29), .A3(new_n345), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n348), .A2(new_n349), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n240), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n218), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n314), .A2(G214), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT83), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n314), .A2(new_n370), .A3(G214), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n261), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n223), .A3(G143), .A4(G214), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n314), .A2(KEYINPUT84), .A3(G143), .A4(G214), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n271), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n378), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G131), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n378), .A3(new_n271), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n367), .B(new_n380), .C1(new_n384), .C2(KEYINPUT17), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n206), .A2(new_n208), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n214), .B1(new_n386), .B2(new_n213), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT18), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n271), .ZN(new_n389));
  OAI221_X1 g203(.A(new_n387), .B1(new_n389), .B2(new_n381), .C1(new_n382), .C2(new_n388), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT85), .B(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n387), .B1(new_n381), .B2(new_n389), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(KEYINPUT18), .B2(new_n379), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT19), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n212), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n386), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n211), .B1(new_n400), .B2(G146), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n382), .B2(new_n383), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n393), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G475), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n228), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT86), .B1(new_n395), .B2(new_n403), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(KEYINPUT20), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n411));
  AOI21_X1  g225(.A(G475), .B1(new_n395), .B2(new_n403), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n228), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n385), .A2(new_n390), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n393), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT87), .A3(new_n395), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n417), .A3(new_n393), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n228), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n408), .A2(new_n413), .B1(new_n419), .B2(G475), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n187), .B1(new_n258), .B2(new_n260), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT89), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n257), .A2(G128), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n429), .B(new_n422), .C1(new_n292), .C2(new_n187), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G116), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n241), .B2(new_n432), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n434), .A2(G107), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(G107), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n431), .A2(G134), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n275), .B(new_n427), .C1(new_n292), .C2(new_n187), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT14), .B(G122), .C1(new_n246), .C2(new_n247), .ZN(new_n440));
  OAI211_X1 g254(.A(G107), .B(new_n440), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n441));
  OAI21_X1  g255(.A(G134), .B1(new_n424), .B2(new_n426), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n435), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT9), .B(G234), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n447), .A2(new_n232), .A3(G953), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n444), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n437), .B2(new_n438), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n448), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n421), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G221), .B1(new_n447), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n228), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n294), .A2(new_n297), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT76), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n187), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n262), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n255), .B1(new_n292), .B2(new_n213), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n289), .B1(new_n292), .B2(new_n213), .ZN(new_n470));
  OAI211_X1 g284(.A(KEYINPUT76), .B(new_n469), .C1(new_n470), .C2(new_n187), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G104), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT3), .B1(new_n473), .B2(G107), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n475));
  INV_X1    g289(.A(G107), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(G104), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(G107), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(G101), .ZN(new_n480));
  INV_X1    g294(.A(new_n478), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n473), .A2(G107), .ZN(new_n482));
  OAI21_X1  g296(.A(G101), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n472), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n298), .A2(new_n484), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n464), .B1(new_n488), .B2(new_n330), .ZN(new_n489));
  INV_X1    g303(.A(new_n330), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT12), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n490), .B(new_n492), .C1(new_n486), .C2(new_n487), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT79), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G140), .ZN(new_n495));
  INV_X1    g309(.A(G227), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n495), .B(new_n497), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT10), .B1(new_n472), .B2(new_n485), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n479), .A2(new_n501), .A3(G101), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT75), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT75), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n479), .A2(new_n504), .A3(new_n501), .A4(G101), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n501), .B1(new_n479), .B2(G101), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n480), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n506), .A2(new_n332), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n298), .A2(new_n510), .A3(new_n484), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n500), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n499), .B1(new_n512), .B2(new_n490), .ZN(new_n513));
  INV_X1    g327(.A(new_n492), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n468), .A2(new_n471), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n484), .B1(new_n515), .B2(new_n465), .ZN(new_n516));
  INV_X1    g330(.A(new_n487), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n330), .B(new_n514), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT79), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n490), .B1(new_n486), .B2(new_n487), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n464), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n494), .A2(new_n513), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT80), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n494), .A2(new_n521), .A3(new_n524), .A4(new_n513), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT78), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n512), .B2(new_n490), .ZN(new_n528));
  INV_X1    g342(.A(new_n509), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n327), .A2(KEYINPUT10), .A3(new_n485), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n529), .B(new_n530), .C1(new_n516), .C2(KEYINPUT10), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT78), .A3(new_n330), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n512), .A2(new_n490), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n498), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n463), .B1(new_n537), .B2(new_n462), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n533), .A2(new_n513), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(new_n489), .B2(new_n493), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n499), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n541), .A3(G469), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n461), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n270), .A2(new_n265), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G125), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n327), .B2(G125), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n223), .A2(G224), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n546), .B(new_n548), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n503), .A2(new_n505), .B1(new_n480), .B2(new_n507), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n252), .B2(new_n253), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT5), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n193), .A3(G116), .ZN(new_n553));
  OAI211_X1 g367(.A(G113), .B(new_n553), .C1(new_n249), .C2(new_n552), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n242), .A2(new_n248), .A3(new_n309), .A4(new_n243), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n485), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(G110), .B(G122), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n555), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n485), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n557), .B(KEYINPUT8), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n549), .B(new_n559), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n551), .A2(new_n556), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n564), .A2(new_n557), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n558), .B(new_n566), .C1(new_n551), .C2(new_n556), .ZN(new_n567));
  INV_X1    g381(.A(new_n559), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n546), .B(new_n547), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n228), .B(new_n563), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n564), .A2(new_n557), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n566), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n564), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n557), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n559), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n570), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n574), .A3(new_n563), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(G234), .A2(G237), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(G952), .A3(new_n223), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT90), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT21), .B(G898), .Z(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(G902), .A3(G953), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G214), .B1(G237), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n366), .A2(new_n459), .A3(new_n543), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(new_n543), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n348), .A2(new_n228), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n364), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n598), .A2(new_n240), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT91), .B1(new_n582), .B2(new_n563), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n593), .B1(new_n603), .B2(new_n572), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT91), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n571), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n582), .A2(KEYINPUT91), .A3(new_n563), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n573), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT92), .B1(new_n452), .B2(new_n448), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n445), .A2(new_n449), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n452), .A2(new_n448), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n610), .B(KEYINPUT33), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n450), .B(new_n453), .C1(KEYINPUT92), .C2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(G478), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n455), .A2(new_n228), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n454), .A2(new_n455), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n420), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n609), .A2(new_n591), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n602), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n419), .A2(G475), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT20), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n406), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n406), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n458), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n604), .A3(new_n590), .A4(new_n608), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n602), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n221), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n228), .A3(new_n238), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n644), .A2(KEYINPUT96), .A3(new_n228), .A4(new_n238), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n236), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n601), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n543), .A2(new_n651), .A3(new_n459), .A4(new_n595), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT97), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n354), .A2(new_n365), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n585), .A2(new_n657), .A3(G902), .A4(G953), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT98), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n587), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n635), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n609), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n543), .A2(new_n656), .A3(new_n649), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n660), .B(KEYINPUT39), .Z(new_n665));
  NOR2_X1   g479(.A1(new_n598), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n649), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n584), .B(KEYINPUT99), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT38), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n420), .A2(new_n457), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n593), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT40), .B1(new_n598), .B2(new_n665), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n364), .A2(new_n363), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n345), .B1(new_n334), .B2(new_n335), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n228), .B1(new_n319), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(G472), .ZN(new_n678));
  INV_X1    g492(.A(new_n349), .ZN(new_n679));
  INV_X1    g493(.A(new_n338), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n339), .B1(new_n319), .B2(new_n320), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n346), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n679), .B1(new_n683), .B2(new_n321), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n352), .B1(new_n684), .B2(KEYINPUT32), .ZN(new_n685));
  INV_X1    g499(.A(new_n353), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n675), .B(new_n678), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n354), .A2(new_n689), .A3(new_n675), .A4(new_n678), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n668), .A2(new_n673), .A3(new_n674), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n261), .B(KEYINPUT101), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G45));
  AOI21_X1  g508(.A(new_n650), .B1(new_n354), .B2(new_n365), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n609), .A2(new_n622), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n543), .A3(new_n696), .A4(new_n660), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  NAND2_X1  g512(.A1(new_n526), .A2(new_n536), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n462), .A3(new_n228), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n535), .B1(new_n523), .B2(new_n525), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n702), .A3(new_n460), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n366), .A2(new_n623), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  OAI211_X1 g521(.A(new_n366), .B(new_n704), .C1(new_n638), .C2(new_n639), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR2_X1   g523(.A1(new_n703), .A2(new_n609), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n421), .A2(new_n458), .A3(new_n591), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n695), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  INV_X1    g527(.A(new_n240), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n356), .A2(KEYINPUT102), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n336), .B2(new_n337), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n318), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n346), .A2(KEYINPUT31), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n321), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n349), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n600), .A2(new_n714), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n710), .A2(new_n590), .A3(new_n671), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  AOI21_X1  g538(.A(G902), .B1(new_n683), .B2(new_n321), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n649), .B(new_n721), .C1(new_n725), .C2(new_n355), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT103), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n600), .A2(new_n728), .A3(new_n649), .A4(new_n721), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n660), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n622), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n710), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n701), .A2(G469), .A3(G902), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n542), .A2(KEYINPUT104), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n513), .A2(new_n533), .B1(new_n540), .B2(new_n499), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(G469), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n736), .A2(new_n463), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT105), .B1(new_n742), .B2(new_n461), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n576), .A2(new_n583), .A3(new_n592), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n576), .A2(new_n583), .A3(KEYINPUT106), .A4(new_n592), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n463), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n739), .B1(new_n738), .B2(G469), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n739), .A2(new_n539), .A3(G469), .A4(new_n541), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n700), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n460), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n743), .A2(new_n366), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n732), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n735), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI211_X1 g573(.A(KEYINPUT105), .B(new_n461), .C1(new_n538), .C2(new_n753), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n755), .B1(new_n754), .B2(new_n460), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n240), .B1(new_n365), .B2(new_n350), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n758), .A2(new_n735), .A3(new_n748), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR3_X1   g581(.A1(new_n760), .A2(new_n761), .A3(new_n748), .ZN(new_n768));
  INV_X1    g582(.A(new_n661), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(KEYINPUT107), .A3(new_n366), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n757), .B2(new_n661), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT108), .B(G134), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G36));
  OAI21_X1  g589(.A(G469), .B1(new_n738), .B2(KEYINPUT45), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT109), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n738), .A2(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT46), .B1(new_n779), .B2(new_n750), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n736), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n460), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n665), .ZN(new_n785));
  INV_X1    g599(.A(new_n620), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n420), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n601), .A3(new_n649), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n749), .A3(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n785), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n784), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n758), .A2(new_n748), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n354), .A2(new_n365), .A3(new_n240), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n609), .A2(new_n672), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n660), .B(KEYINPUT115), .Z(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n688), .B2(new_n690), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n742), .A2(new_n461), .A3(new_n649), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n733), .A2(new_n663), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n733), .A2(new_n663), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n814), .A2(new_n816), .A3(new_n697), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n733), .A2(new_n663), .A3(new_n817), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n733), .B2(new_n663), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n697), .A4(new_n814), .ZN(new_n825));
  INV_X1    g639(.A(new_n697), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n812), .A2(new_n813), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n820), .A2(new_n825), .B1(new_n808), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n708), .A2(new_n723), .A3(new_n712), .A4(new_n705), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n759), .B2(new_n765), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n457), .A2(new_n628), .A3(new_n660), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n746), .A2(new_n634), .A3(new_n747), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n695), .A2(new_n543), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n834), .A2(new_n835), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n695), .A2(new_n836), .A3(new_n543), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT113), .B1(new_n842), .B2(new_n839), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n621), .A2(new_n584), .A3(new_n594), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n621), .A2(new_n584), .A3(KEYINPUT111), .A4(new_n594), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n584), .A2(new_n458), .A3(new_n420), .A4(new_n594), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n601), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n543), .A3(new_n714), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n596), .A2(new_n852), .A3(new_n652), .ZN(new_n853));
  INV_X1    g667(.A(new_n730), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n758), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n853), .B1(new_n855), .B2(new_n768), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n832), .A2(new_n773), .A3(new_n844), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n807), .B1(new_n830), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n829), .A2(new_n808), .B1(new_n827), .B2(new_n814), .ZN(new_n859));
  XNOR2_X1  g673(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n806), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n857), .B2(new_n859), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n770), .A2(new_n772), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n768), .A2(new_n855), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n596), .A2(new_n652), .A3(new_n852), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n838), .B1(new_n837), .B2(new_n840), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n842), .A2(KEYINPUT113), .A3(new_n839), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n743), .A2(new_n764), .A3(new_n756), .A4(new_n763), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n762), .A2(new_n366), .A3(new_n732), .A4(new_n749), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n735), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT118), .B1(new_n874), .B2(new_n831), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n832), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n871), .A2(new_n875), .A3(KEYINPUT53), .A4(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n864), .B(new_n806), .C1(new_n878), .C2(new_n830), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n863), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n587), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n789), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n722), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n710), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n700), .A2(new_n702), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n460), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n749), .B(new_n885), .C1(new_n800), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n703), .A2(new_n748), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n730), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n670), .A2(new_n593), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n892), .A2(new_n703), .A3(new_n884), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n893), .A2(KEYINPUT50), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(KEYINPUT50), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n691), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n714), .A3(new_n882), .A4(new_n890), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n421), .A3(new_n786), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n889), .A2(KEYINPUT51), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT51), .B1(new_n889), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n223), .A2(G952), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n883), .A2(new_n763), .A3(new_n890), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT48), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI221_X1 g720(.A(new_n906), .B1(new_n905), .B2(new_n904), .C1(new_n898), .C2(new_n622), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n881), .A2(new_n886), .A3(new_n901), .A4(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(G952), .B2(G953), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n787), .A2(new_n461), .A3(new_n593), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n887), .B2(KEYINPUT49), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(KEYINPUT49), .B2(new_n887), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n897), .A2(new_n714), .A3(new_n670), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(G75));
  NAND2_X1  g729(.A1(new_n829), .A2(new_n808), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n824), .B1(new_n917), .B2(new_n814), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n773), .A2(new_n856), .A3(new_n844), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n876), .B2(new_n832), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n228), .B1(new_n924), .B2(new_n864), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n580), .B(new_n570), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(KEYINPUT119), .B2(KEYINPUT56), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n926), .A2(new_n930), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n223), .A2(G952), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(G51));
  AOI211_X1 g748(.A(new_n228), .B(new_n779), .C1(new_n924), .C2(new_n864), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n463), .B(KEYINPUT57), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n806), .B1(new_n924), .B2(new_n864), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n880), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n938), .B2(new_n699), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT120), .B1(new_n939), .B2(new_n933), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  INV_X1    g755(.A(new_n933), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n864), .B1(new_n878), .B2(new_n830), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n879), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n701), .B1(new_n945), .B2(new_n936), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n941), .B(new_n942), .C1(new_n946), .C2(new_n935), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n940), .A2(new_n947), .ZN(G54));
  NAND3_X1  g762(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  INV_X1    g763(.A(new_n404), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n933), .ZN(G60));
  AND2_X1   g767(.A1(new_n613), .A2(new_n615), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n617), .B(KEYINPUT59), .Z(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n863), .B2(new_n880), .ZN(new_n956));
  INV_X1    g770(.A(new_n954), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n957), .B(new_n955), .C1(new_n937), .C2(new_n880), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT121), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n945), .A2(new_n960), .A3(new_n957), .A4(new_n955), .ZN(new_n961));
  AOI221_X4 g775(.A(new_n933), .B1(new_n954), .B2(new_n956), .C1(new_n959), .C2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND3_X1  g778(.A1(new_n943), .A2(new_n644), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n943), .A2(new_n964), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n942), .B(new_n965), .C1(new_n966), .C2(new_n237), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT61), .B1(new_n967), .B2(KEYINPUT122), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  NAND2_X1  g785(.A1(new_n588), .A2(G224), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(G953), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n831), .A2(new_n853), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n569), .B1(G898), .B2(new_n223), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  NAND3_X1  g791(.A1(new_n804), .A2(new_n773), .A3(new_n917), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n795), .A2(new_n796), .B1(new_n763), .B2(new_n809), .ZN(new_n979));
  INV_X1    g793(.A(new_n785), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n766), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n223), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n304), .A2(new_n306), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n400), .B(KEYINPUT123), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n982), .B(new_n985), .C1(G900), .C2(new_n223), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n917), .A2(new_n692), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n622), .B1(new_n457), .B2(new_n421), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n666), .A2(new_n366), .A3(new_n749), .A4(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n797), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n992), .A3(new_n804), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT124), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n989), .A2(new_n992), .A3(new_n995), .A4(new_n804), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n985), .A2(G953), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n986), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n496), .B2(new_n657), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n986), .B(new_n1002), .C1(new_n997), .C2(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G72));
  XNOR2_X1  g818(.A(new_n358), .B(KEYINPUT126), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n978), .A2(new_n981), .A3(new_n831), .A4(new_n853), .ZN(new_n1006));
  XNOR2_X1  g820(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n355), .A2(new_n228), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1007), .B(new_n1008), .Z(new_n1009));
  OAI211_X1 g823(.A(new_n318), .B(new_n1005), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n858), .A2(new_n862), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1009), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n359), .A2(new_n346), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1010), .A2(new_n1014), .A3(new_n942), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n994), .A2(new_n974), .A3(new_n996), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1005), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n345), .B2(new_n1017), .ZN(G57));
endmodule


