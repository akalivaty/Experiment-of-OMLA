//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n459), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(new_n462), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(KEYINPUT70), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  OR2_X1    g048(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n465), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n470), .A2(new_n471), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n475), .A2(new_n480), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n475), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(G124), .A2(new_n485), .B1(new_n486), .B2(G136), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n480), .C2(G112), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n459), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n475), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n466), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n480), .A2(new_n497), .A3(new_n498), .A4(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n506), .B2(KEYINPUT72), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(new_n516), .B1(new_n504), .B2(new_n505), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n503), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  AOI22_X1  g093(.A1(G88), .A2(new_n517), .B1(new_n518), .B2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n511), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND2_X1  g096(.A1(new_n517), .A2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n504), .A2(new_n505), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n528), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n522), .A2(new_n523), .A3(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n518), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n514), .A2(new_n516), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n524), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n532), .B1(new_n534), .B2(new_n535), .C1(new_n513), .C2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n504), .A2(new_n505), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(G81), .B2(new_n517), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT73), .B(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n518), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n518), .A2(G53), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n518), .A2(new_n555), .A3(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n540), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(G91), .B2(new_n517), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g138(.A1(G168), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n522), .A2(new_n523), .A3(new_n530), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  NAND2_X1  g143(.A1(new_n517), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n518), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n540), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n517), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n518), .A2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n517), .A2(G85), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n513), .C2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT75), .B(G66), .Z(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n540), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT10), .B1(new_n534), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n517), .A2(new_n591), .A3(G92), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n518), .A2(G54), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n588), .A2(new_n590), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n584), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n584), .B1(new_n595), .B2(G868), .ZN(G321));
  NOR2_X1   g172(.A1(G299), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G868), .B2(new_n567), .ZN(G297));
  AOI21_X1  g174(.A(new_n598), .B1(G868), .B2(new_n567), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n546), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n587), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n605), .A2(new_n601), .A3(new_n592), .A4(new_n590), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n607), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g184(.A1(G123), .A2(new_n485), .B1(new_n486), .B2(G135), .ZN(new_n610));
  OAI221_X1 g185(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n480), .C2(G111), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2096), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n615), .B(new_n616), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT77), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n614), .B(new_n621), .C1(new_n619), .C2(new_n618), .ZN(G156));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G1341), .B(G1348), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n632), .A2(new_n635), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT18), .Z(new_n644));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n641), .ZN(new_n647));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n641), .B(KEYINPUT17), .Z(new_n649));
  INV_X1    g224(.A(new_n642), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n640), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT81), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n658), .A2(new_n663), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n666));
  AOI211_X1 g241(.A(new_n662), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n665), .B2(new_n666), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G23), .ZN(new_n680));
  INV_X1    g255(.A(G288), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT33), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1976), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n679), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(G1971), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(G1971), .ZN(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n684), .A2(new_n687), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n694));
  AOI22_X1  g269(.A1(G119), .A2(new_n485), .B1(new_n486), .B2(G131), .ZN(new_n695));
  OAI221_X1 g270(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n480), .C2(G107), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G25), .B(new_n697), .S(G29), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT83), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1986), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n693), .A2(new_n694), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT31), .B(G11), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(G28), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT30), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n708), .B1(new_n710), .B2(new_n713), .C1(new_n612), .C2(new_n712), .ZN(new_n714));
  NOR2_X1   g289(.A1(G162), .A2(new_n712), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n712), .B2(G35), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT29), .B(G2090), .Z(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT24), .B(G34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(new_n712), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT87), .Z(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n483), .B2(new_n712), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n718), .B1(new_n716), .B2(new_n717), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n712), .A2(G26), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT28), .Z(new_n727));
  AOI22_X1  g302(.A1(G128), .A2(new_n485), .B1(new_n486), .B2(G140), .ZN(new_n728));
  OAI221_X1 g303(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n480), .C2(G116), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT84), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n727), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT85), .B(G2067), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n679), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n679), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1966), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n679), .A2(G5), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G171), .B2(new_n679), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n737), .B1(G1961), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G4), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n595), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1348), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n679), .A2(G20), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT23), .Z(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G299), .B2(G16), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AND4_X1   g324(.A1(new_n734), .A2(new_n740), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n712), .A2(G32), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n486), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n485), .A2(G129), .ZN(new_n757));
  AND4_X1   g332(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(new_n712), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G16), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n547), .B2(G16), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(G1341), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n712), .A2(G33), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  INV_X1    g344(.A(G127), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n475), .B2(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n771), .A2(new_n481), .B1(new_n486), .B2(G139), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n765), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT86), .B(G2072), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G1961), .B2(new_n739), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n763), .A2(G1341), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n774), .B2(new_n775), .ZN(new_n779));
  NOR2_X1   g354(.A1(G27), .A2(G29), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G164), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT90), .B(G2078), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n764), .A2(new_n777), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n725), .A2(new_n750), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n707), .A2(new_n785), .ZN(G150));
  INV_X1    g361(.A(G150), .ZN(G311));
  NOR2_X1   g362(.A1(new_n594), .A2(new_n601), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n518), .A2(G55), .ZN(new_n791));
  INV_X1    g366(.A(G93), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n791), .B1(new_n534), .B2(new_n792), .C1(new_n513), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n793), .A2(new_n513), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n534), .A2(new_n792), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n798), .A2(new_n545), .A3(new_n543), .A4(new_n791), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n790), .B(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n801), .A2(KEYINPUT39), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(KEYINPUT39), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n802), .A2(new_n803), .A3(G860), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n794), .A2(G860), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT37), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n806), .ZN(G145));
  XNOR2_X1  g382(.A(new_n483), .B(new_n612), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(new_n489), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n496), .A2(new_n499), .ZN(new_n810));
  INV_X1    g385(.A(new_n494), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n773), .A2(KEYINPUT93), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(new_n758), .Z(new_n814));
  INV_X1    g389(.A(new_n731), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n814), .A2(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(new_n815), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n819), .A2(G164), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n485), .A2(G130), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT94), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n486), .A2(G142), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n480), .A2(G118), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n697), .ZN(new_n829));
  INV_X1    g404(.A(new_n617), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(KEYINPUT95), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n809), .B1(new_n822), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n818), .B(new_n821), .C1(KEYINPUT95), .C2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n822), .A2(new_n831), .ZN(new_n836));
  INV_X1    g411(.A(new_n831), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n837), .A2(new_n821), .A3(new_n818), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n809), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT96), .B(KEYINPUT40), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(G395));
  OR2_X1    g418(.A1(G290), .A2(G288), .ZN(new_n844));
  NAND2_X1  g419(.A1(G290), .A2(G288), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n844), .A2(KEYINPUT100), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT100), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(G303), .A2(G305), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n575), .A2(G651), .B1(G48), .B2(new_n518), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n511), .A2(new_n849), .A3(new_n519), .A4(new_n577), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n846), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n681), .B(G290), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n851), .A2(new_n853), .A3(KEYINPUT100), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n800), .A2(new_n607), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n795), .A2(new_n799), .A3(new_n606), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(G299), .A2(new_n592), .A3(new_n590), .A4(new_n605), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n594), .A2(new_n861), .A3(new_n557), .A4(new_n561), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G299), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n861), .B1(new_n864), .B2(new_n594), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT98), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT97), .B1(new_n595), .B2(G299), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n860), .A3(new_n862), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n869), .A2(new_n870), .A3(new_n857), .A4(new_n858), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n863), .B2(new_n865), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n868), .A2(KEYINPUT41), .A3(new_n860), .A4(new_n862), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT99), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n869), .A2(new_n878), .A3(new_n874), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n859), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n872), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n873), .B1(new_n872), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n856), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n881), .A3(new_n855), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G868), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n794), .A2(new_n603), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(G295));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n891), .A3(new_n889), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n603), .B1(new_n884), .B2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(new_n889), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT101), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  NAND2_X1  g472(.A1(G301), .A2(new_n565), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n800), .B(new_n898), .C1(G286), .C2(G301), .ZN(new_n899));
  AOI21_X1  g474(.A(G301), .B1(new_n564), .B2(new_n566), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n795), .B(new_n799), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n877), .A2(new_n903), .A3(new_n879), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n869), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n855), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n852), .B2(new_n854), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n844), .A2(new_n845), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n844), .A2(KEYINPUT100), .A3(new_n845), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n848), .A4(new_n850), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n851), .A2(new_n853), .A3(KEYINPUT100), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT103), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n910), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n897), .B1(new_n909), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n875), .A2(new_n876), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n906), .B1(new_n923), .B2(new_n905), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n907), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n909), .A2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n910), .A2(new_n920), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n931), .A2(new_n840), .A3(new_n907), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n932), .B2(new_n908), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(new_n897), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n908), .B1(new_n921), .B2(new_n907), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n920), .A2(new_n924), .ZN(new_n936));
  AND4_X1   g511(.A1(new_n840), .A2(new_n936), .A3(new_n907), .A4(new_n908), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n929), .B(new_n897), .C1(new_n935), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n928), .B1(new_n934), .B2(new_n939), .ZN(G397));
  OR3_X1    g515(.A1(G164), .A2(KEYINPUT105), .A3(G1384), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT105), .B1(G164), .B2(G1384), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT106), .B(G40), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n470), .A2(new_n471), .A3(new_n482), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n758), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n731), .B(G2067), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n951), .A2(new_n952), .A3(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n951), .B2(new_n947), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n957), .B(new_n950), .C1(new_n953), .C2(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(new_n947), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n697), .B(new_n700), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n956), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(G290), .B(G1986), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n947), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n470), .A2(KEYINPUT123), .A3(new_n471), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT123), .B1(new_n470), .B2(new_n471), .ZN(new_n965));
  INV_X1    g540(.A(G2078), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n482), .A2(KEYINPUT53), .A3(G40), .A4(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n812), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n944), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n972));
  AND4_X1   g547(.A1(new_n470), .A2(new_n471), .A3(new_n482), .A4(new_n945), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n942), .B1(G164), .B2(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n975), .B2(G2078), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n812), .A2(new_n977), .A3(new_n969), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1961), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n971), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G171), .ZN(new_n984));
  INV_X1    g559(.A(new_n975), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(KEYINPUT53), .A3(new_n966), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(new_n976), .A3(G301), .A4(new_n982), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(KEYINPUT54), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT124), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT124), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n984), .A2(new_n990), .A3(KEYINPUT54), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT109), .B(G1971), .Z(new_n993));
  NAND2_X1  g568(.A1(new_n975), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n977), .B1(new_n812), .B2(new_n969), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT113), .B1(new_n995), .B2(new_n946), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n973), .A2(new_n979), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n978), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(G2090), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n975), .A2(KEYINPUT110), .A3(new_n993), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n1009), .C1(G2090), .C2(new_n980), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1005), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(G8), .A3(new_n1011), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n946), .A2(G1384), .A3(G164), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1976), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT111), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT52), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1016), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1015), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(G305), .A2(G1981), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G305), .A2(G1981), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1015), .A3(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1020), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1006), .A2(new_n1012), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1966), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n975), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n978), .A2(new_n979), .A3(new_n973), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n723), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n975), .A2(KEYINPUT114), .A3(new_n1032), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1035), .A2(G168), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1014), .B1(KEYINPUT121), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT51), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT114), .B1(new_n975), .B2(new_n1032), .ZN(new_n1046));
  OAI211_X1 g621(.A(G8), .B(new_n565), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1039), .B(new_n1041), .C1(KEYINPUT121), .C2(new_n1040), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n976), .A2(new_n982), .ZN(new_n1051));
  AOI21_X1  g626(.A(G301), .B1(new_n1051), .B2(new_n986), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n983), .A2(G171), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n992), .A2(new_n1031), .A3(new_n1049), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n561), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n561), .A2(new_n1056), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n557), .B(KEYINPUT116), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1059), .A2(new_n1060), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT56), .B(G2072), .Z(new_n1062));
  OR2_X1    g637(.A1(new_n975), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1956), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n998), .A2(new_n978), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n997), .B1(new_n973), .B2(new_n979), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT115), .B(new_n1066), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT115), .B1(new_n999), .B2(new_n1066), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1065), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT61), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1069), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1061), .B1(new_n1077), .B2(new_n1063), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT119), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1064), .B1(new_n1076), .B2(new_n1069), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1063), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1061), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1080), .B1(new_n1077), .B2(new_n1065), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT58), .B(G1341), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n975), .A2(G1996), .B1(new_n1013), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n547), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G2067), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1013), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(KEYINPUT60), .C1(new_n1036), .C2(G1348), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1096), .A2(KEYINPUT120), .A3(new_n594), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n594), .B1(new_n1096), .B2(KEYINPUT120), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1097), .A2(new_n1098), .B1(KEYINPUT120), .B2(new_n1096), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n980), .A2(new_n743), .B1(new_n1013), .B2(new_n1094), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1093), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1079), .A2(new_n1082), .A3(new_n1088), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1100), .A2(new_n594), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1106), .B2(new_n1081), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT118), .B(new_n1072), .C1(new_n1078), .C2(new_n1105), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1055), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1048), .A2(new_n1047), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT121), .B(new_n1040), .C1(new_n1039), .C2(G8), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT62), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n1006), .A2(new_n1012), .A3(new_n1030), .A4(new_n1052), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1044), .A2(new_n1115), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(G8), .B(new_n567), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1006), .A2(new_n1119), .A3(new_n1012), .A4(new_n1030), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1010), .A2(G8), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1005), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1012), .A4(new_n1030), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1029), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1023), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1014), .B(new_n1013), .C1(new_n1130), .C2(KEYINPUT112), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1130), .A2(KEYINPUT112), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1012), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1131), .A2(new_n1132), .B1(new_n1133), .B2(new_n1030), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1117), .A2(new_n1127), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n963), .B1(new_n1110), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n959), .A2(G1986), .A3(G290), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1138));
  XNOR2_X1  g713(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT46), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n758), .B1(new_n1140), .B2(G1996), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n947), .B1(new_n951), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n947), .A2(new_n948), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT125), .A3(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT125), .B1(new_n1143), .B2(new_n1140), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1148));
  AND2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n961), .A2(new_n1139), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n695), .A2(new_n700), .A3(new_n696), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n956), .A2(new_n958), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n815), .A2(new_n1094), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n959), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g732(.A(G319), .B1(new_n637), .B2(new_n638), .ZN(new_n1159));
  AOI211_X1 g733(.A(G227), .B(new_n1159), .C1(new_n676), .C2(new_n677), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n1160), .A2(new_n841), .A3(new_n933), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


