//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(G217), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT92), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n192), .B(new_n198), .C1(new_n194), .C2(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(new_n192), .ZN(new_n200));
  INV_X1    g014(.A(new_n195), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n191), .A2(KEYINPUT91), .A3(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n197), .A2(new_n199), .A3(new_n202), .A4(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G134), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT65), .B(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n210), .A3(new_n200), .ZN(new_n211));
  INV_X1    g025(.A(G122), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G122), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n215), .A3(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(KEYINPUT14), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n223), .A3(G107), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n213), .B(new_n215), .C1(KEYINPUT14), .C2(new_n217), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n207), .A2(new_n200), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n211), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n190), .B1(new_n222), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n220), .B1(G134), .B2(new_n208), .ZN(new_n237));
  INV_X1    g051(.A(new_n190), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n237), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n187), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT93), .ZN(new_n241));
  INV_X1    g055(.A(G478), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT15), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n222), .A2(new_n235), .A3(new_n190), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n238), .B1(new_n237), .B2(new_n234), .ZN(new_n245));
  AOI21_X1  g059(.A(G902), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n250), .C1(new_n243), .C2(new_n240), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G952), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(G234), .B2(G237), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT21), .B(G898), .Z(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT95), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n187), .B(new_n254), .C1(G234), .C2(G237), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G140), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G125), .ZN(new_n265));
  INV_X1    g079(.A(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G140), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT64), .B(G146), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(G237), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n254), .A3(G214), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n204), .ZN(new_n275));
  NOR2_X1   g089(.A1(G237), .A2(G953), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(G143), .A3(G214), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT18), .A3(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT18), .A2(G131), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n275), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n272), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(G113), .B(G122), .Z(new_n283));
  XOR2_X1   g097(.A(KEYINPUT87), .B(G104), .Z(new_n284));
  XOR2_X1   g098(.A(new_n283), .B(new_n284), .Z(new_n285));
  NAND3_X1  g099(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT16), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n266), .A2(KEYINPUT16), .A3(G140), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G146), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(G146), .B1(new_n286), .B2(new_n287), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n276), .A2(G143), .A3(G214), .ZN(new_n292));
  AOI21_X1  g106(.A(G143), .B1(new_n276), .B2(G214), .ZN(new_n293));
  OAI21_X1  g107(.A(G131), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G131), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n275), .A2(new_n295), .A3(new_n277), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n294), .A2(new_n296), .A3(KEYINPUT88), .A4(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n275), .B2(new_n277), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT17), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(new_n297), .A3(new_n296), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n282), .B(new_n285), .C1(new_n301), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT89), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n303), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(new_n291), .A3(new_n298), .A4(new_n300), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n282), .A4(new_n285), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n268), .B(KEYINPUT19), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n289), .B1(new_n312), .B2(new_n269), .ZN(new_n313));
  INV_X1    g127(.A(new_n296), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT86), .B1(new_n314), .B2(new_n299), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n314), .A2(KEYINPUT86), .A3(new_n299), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n282), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n285), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n322));
  NOR2_X1   g136(.A1(G475), .A2(G902), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n306), .A2(new_n310), .B1(new_n319), .B2(new_n318), .ZN(new_n325));
  INV_X1    g139(.A(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n285), .B1(new_n308), .B2(new_n282), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n306), .B2(new_n310), .ZN(new_n330));
  OAI21_X1  g144(.A(G475), .B1(new_n330), .B2(G902), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT96), .B1(new_n263), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n332), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT96), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n262), .A4(new_n253), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G221), .ZN(new_n338));
  INV_X1    g152(.A(new_n188), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n187), .ZN(new_n340));
  INV_X1    g154(.A(G469), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n187), .ZN(new_n342));
  XNOR2_X1  g156(.A(G110), .B(G140), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n254), .A2(G227), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G137), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n229), .A2(new_n231), .A3(new_n347), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(KEYINPUT11), .A3(G134), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G131), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n229), .A2(new_n231), .A3(new_n347), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n295), .A3(new_n350), .A4(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(KEYINPUT66), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT66), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(G131), .C1(new_n348), .C2(new_n351), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT75), .B(G104), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT3), .B1(new_n359), .B2(G107), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n217), .A3(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(new_n361), .A3(new_n217), .A4(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT77), .B(G101), .ZN(new_n367));
  INV_X1    g181(.A(G104), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G104), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n371), .A3(G107), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n360), .A2(new_n366), .A3(new_n367), .A4(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(G107), .B1(new_n369), .B2(new_n371), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n217), .A2(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(G101), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n271), .A2(KEYINPUT64), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT64), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G146), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(G143), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n191), .B1(new_n381), .B2(KEYINPUT1), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n204), .A2(G146), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(new_n380), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n204), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n381), .B(new_n387), .C1(G143), .C2(new_n271), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n271), .A2(G143), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n269), .B2(G143), .ZN(new_n391));
  INV_X1    g205(.A(new_n383), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n191), .B1(new_n392), .B2(KEYINPUT1), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n388), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n373), .A3(new_n376), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n358), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT12), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n388), .B1(new_n382), .B2(new_n385), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n402), .A2(KEYINPUT10), .A3(new_n373), .A4(new_n376), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G101), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n369), .A2(new_n371), .A3(G107), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n369), .A2(new_n371), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n217), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n408), .B2(KEYINPUT3), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n405), .B1(new_n409), .B2(new_n366), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n372), .B1(new_n374), .B2(new_n361), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n363), .A2(new_n365), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n413), .B(G101), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n392), .B1(new_n269), .B2(G143), .ZN(new_n417));
  AND2_X1   g231(.A1(KEYINPUT0), .A2(G128), .ZN(new_n418));
  NOR2_X1   g232(.A1(KEYINPUT0), .A2(G128), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n417), .A2(new_n420), .B1(new_n391), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n412), .A2(KEYINPUT78), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n416), .A2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(G101), .B1(new_n414), .B2(new_n415), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n358), .B(new_n404), .C1(new_n423), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n401), .A2(new_n403), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT78), .B1(new_n412), .B2(new_n422), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(new_n424), .A3(new_n427), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT79), .B1(new_n435), .B2(new_n358), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n399), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n430), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(KEYINPUT79), .A3(new_n358), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n345), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n434), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n358), .B1(new_n441), .B2(new_n404), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n345), .A2(new_n437), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n342), .B1(new_n444), .B2(G469), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n438), .B2(new_n439), .ZN(new_n446));
  INV_X1    g260(.A(new_n345), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n345), .B(new_n398), .C1(new_n438), .C2(new_n439), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n341), .B(new_n187), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n340), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n388), .B(new_n266), .C1(new_n382), .C2(new_n385), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n421), .B2(new_n266), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT84), .B(G224), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G953), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n454), .B(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n373), .A2(new_n376), .ZN(new_n459));
  XNOR2_X1  g273(.A(G116), .B(G119), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT2), .B(G113), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G113), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n214), .A2(G119), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n464), .B1(new_n470), .B2(KEYINPUT81), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n469), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT81), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n471), .A2(new_n478), .A3(new_n473), .A4(new_n475), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n459), .A2(new_n463), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n460), .B(new_n462), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(new_n416), .C1(new_n410), .C2(new_n411), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT6), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n483), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(KEYINPUT6), .A3(new_n488), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n458), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n471), .A2(new_n475), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n461), .A2(new_n466), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n463), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n459), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n484), .B(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n477), .A2(new_n463), .A3(new_n479), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(new_n498), .C1(new_n499), .C2(new_n459), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n454), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n454), .A2(new_n501), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n485), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n187), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n492), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n458), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n485), .A2(KEYINPUT6), .B1(new_n487), .B2(new_n488), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n487), .A2(KEYINPUT6), .A3(new_n488), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n505), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n452), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n337), .A2(new_n451), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n276), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n355), .A2(new_n421), .A3(new_n357), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n295), .B1(G134), .B2(G137), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n232), .B2(G137), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n402), .A2(new_n354), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n525), .A3(new_n481), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT69), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT28), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n522), .A2(new_n525), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n482), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n526), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n481), .B1(new_n522), .B2(new_n525), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n528), .B1(new_n537), .B2(KEYINPUT68), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n521), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n522), .A2(new_n541), .A3(new_n525), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n522), .B2(new_n525), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n482), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n526), .A3(new_n521), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT31), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT67), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n544), .A2(KEYINPUT67), .A3(new_n526), .A4(new_n521), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT31), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(G472), .A2(G902), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n532), .A2(new_n539), .A3(new_n521), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT70), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n521), .B1(new_n544), .B2(new_n526), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT29), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n532), .A2(new_n539), .A3(new_n561), .A4(new_n521), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n531), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n529), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n528), .B1(new_n534), .B2(new_n526), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n521), .A2(KEYINPUT29), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G472), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n552), .A2(KEYINPUT32), .A3(new_n553), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n556), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n574));
  INV_X1    g388(.A(G119), .ZN(new_n575));
  OR3_X1    g389(.A1(new_n575), .A2(KEYINPUT71), .A3(G128), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT71), .B1(new_n575), .B2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT24), .B(G110), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n575), .A2(G128), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n578), .B(new_n582), .C1(new_n583), .C2(KEYINPUT23), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n581), .B1(G110), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n288), .A3(new_n270), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(G110), .ZN(new_n587));
  OAI221_X1 g401(.A(new_n587), .B1(new_n579), .B2(new_n580), .C1(new_n289), .C2(new_n290), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n187), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(KEYINPUT72), .A2(KEYINPUT25), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n189), .B1(G234), .B2(new_n187), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n595), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(KEYINPUT73), .A3(new_n595), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n601), .A2(G902), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n574), .B1(new_n602), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n600), .A2(new_n601), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(KEYINPUT74), .C1(new_n610), .C2(new_n608), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n573), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n517), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n367), .ZN(G3));
  NAND3_X1  g433(.A1(new_n241), .A2(new_n242), .A3(new_n248), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n236), .A2(new_n239), .A3(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n244), .B2(new_n245), .ZN(new_n623));
  OAI211_X1 g437(.A(G478), .B(new_n187), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n332), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n515), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n507), .B1(new_n492), .B2(new_n505), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n512), .A2(new_n513), .A3(new_n506), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(KEYINPUT97), .A3(new_n452), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n261), .B(new_n626), .C1(new_n628), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n547), .B2(new_n551), .ZN(new_n635));
  INV_X1    g449(.A(G472), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n554), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n451), .A2(new_n616), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT34), .B(G104), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n328), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n324), .A2(new_n327), .A3(KEYINPUT98), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n253), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n331), .A2(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n331), .A2(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n647), .A2(new_n262), .A3(new_n648), .A4(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT97), .B1(new_n631), .B2(new_n452), .ZN(new_n654));
  INV_X1    g468(.A(new_n452), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n627), .B(new_n655), .C1(new_n629), .C2(new_n630), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n639), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  XNOR2_X1  g476(.A(new_n589), .B(KEYINPUT100), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n609), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(KEYINPUT101), .A3(new_n613), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n610), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n672), .B1(new_n602), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n333), .B2(new_n336), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n516), .A3(new_n451), .A4(new_n638), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(new_n675), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n451), .A2(new_n573), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n256), .B1(new_n260), .B2(new_n682), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n646), .A2(new_n651), .A3(new_n253), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n628), .A2(new_n632), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n191), .ZN(G30));
  XOR2_X1   g502(.A(new_n683), .B(KEYINPUT39), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n451), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT102), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n690), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n670), .A2(new_n613), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT32), .B1(new_n552), .B2(new_n553), .ZN(new_n698));
  INV_X1    g512(.A(new_n553), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n555), .B(new_n699), .C1(new_n547), .C2(new_n551), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n549), .A2(new_n550), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n521), .B1(new_n534), .B2(new_n526), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n187), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n697), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n631), .B(KEYINPUT38), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n334), .A2(new_n253), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n452), .A2(new_n706), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n693), .A2(new_n696), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NOR2_X1   g525(.A1(new_n626), .A2(new_n683), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n685), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n681), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n271), .ZN(G48));
  AOI21_X1  g529(.A(new_n615), .B1(new_n701), .B2(new_n571), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n443), .B1(new_n431), .B2(new_n436), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n345), .B1(new_n440), .B2(new_n399), .ZN(new_n718));
  OAI21_X1  g532(.A(G469), .B1(new_n718), .B2(G902), .ZN(new_n719));
  INV_X1    g533(.A(new_n340), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n450), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n634), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT41), .B(G113), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NOR2_X1   g540(.A1(new_n723), .A2(new_n659), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n214), .ZN(G18));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n721), .B2(new_n657), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n717), .A2(new_n345), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n447), .B(new_n399), .C1(new_n431), .C2(new_n436), .ZN(new_n732));
  AOI211_X1 g546(.A(G469), .B(G902), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n446), .B2(new_n447), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n341), .B1(new_n734), .B2(new_n187), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n685), .A3(KEYINPUT103), .A4(new_n720), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n676), .A2(new_n573), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NAND2_X1  g555(.A1(new_n685), .A2(new_n708), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n719), .A2(new_n262), .A3(new_n720), .A4(new_n450), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n635), .A2(new_n636), .ZN(new_n745));
  INV_X1    g559(.A(new_n521), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n565), .B2(new_n566), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT105), .B1(new_n551), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n545), .A2(KEYINPUT31), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n551), .A2(KEYINPUT105), .A3(new_n747), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n553), .B(KEYINPUT104), .Z(new_n753));
  AOI21_X1  g567(.A(new_n745), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n602), .A2(new_n611), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT106), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n745), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n751), .A2(new_n750), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n753), .B1(new_n758), .B2(new_n748), .ZN(new_n759));
  AND4_X1   g573(.A1(KEYINPUT106), .A2(new_n757), .A3(new_n759), .A4(new_n755), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n744), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n759), .A3(new_n697), .A4(new_n712), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n730), .B2(new_n737), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n266), .ZN(G27));
  NAND3_X1  g579(.A1(new_n629), .A2(new_n452), .A3(new_n630), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n340), .B(new_n766), .C1(new_n445), .C2(new_n450), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n716), .A2(new_n767), .A3(new_n768), .A4(new_n712), .ZN(new_n769));
  INV_X1    g583(.A(new_n342), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n443), .B(new_n447), .C1(new_n431), .C2(new_n436), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n398), .B1(new_n438), .B2(new_n439), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n771), .B(G469), .C1(new_n447), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n450), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n766), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n774), .A2(new_n712), .A3(new_n720), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT107), .B1(new_n617), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n769), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n776), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n556), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n572), .A4(new_n571), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n780), .A2(KEYINPUT42), .A3(new_n784), .A4(new_n755), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NAND3_X1  g601(.A1(new_n573), .A2(new_n616), .A3(new_n684), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n451), .A2(new_n775), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n228), .ZN(G36));
  AOI21_X1  g605(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n325), .A2(KEYINPUT20), .A3(new_n326), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n625), .B(new_n331), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n637), .A3(KEYINPUT44), .A4(new_n697), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n775), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT109), .A3(new_n775), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n772), .A2(new_n447), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n345), .B(new_n442), .C1(new_n438), .C2(new_n439), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n771), .B(KEYINPUT45), .C1(new_n447), .C2(new_n772), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(G469), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n770), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n733), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(KEYINPUT46), .A3(new_n770), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n340), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n796), .A2(new_n637), .A3(new_n697), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n802), .A2(new_n689), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  NAND3_X1  g632(.A1(new_n712), .A2(new_n615), .A3(new_n775), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n573), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT110), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n811), .A2(new_n812), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT47), .B1(new_n822), .B2(new_n720), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n827), .B(new_n821), .C1(new_n823), .C2(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n716), .B(new_n722), .C1(new_n658), .C2(new_n633), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n740), .A2(new_n761), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n740), .A2(new_n761), .A3(KEYINPUT112), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n626), .B1(new_n332), .B2(new_n253), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n262), .A3(new_n516), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n639), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n677), .C1(new_n617), .C2(new_n517), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n451), .A2(new_n680), .ZN(new_n844));
  INV_X1    g658(.A(new_n686), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n685), .A2(new_n712), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n844), .B(new_n573), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n742), .ZN(new_n848));
  INV_X1    g662(.A(new_n683), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n706), .A3(new_n451), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n738), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n847), .B(new_n850), .C1(new_n851), .C2(new_n763), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n647), .A2(new_n253), .A3(new_n652), .A4(new_n849), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT113), .B1(new_n854), .B2(new_n766), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n648), .A2(new_n651), .A3(new_n683), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n647), .A4(new_n775), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n859), .A2(new_n681), .B1(new_n789), .B2(new_n788), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n754), .A2(new_n697), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT114), .B1(new_n861), .B2(new_n776), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n861), .A2(KEYINPUT114), .A3(new_n776), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n681), .B1(new_n686), .B2(new_n713), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n764), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n850), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n853), .A2(new_n864), .A3(new_n868), .A4(new_n786), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n831), .B1(new_n843), .B2(new_n869), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(KEYINPUT115), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n853), .A2(new_n868), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n864), .A2(new_n786), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n842), .A3(new_n837), .A4(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n870), .B(KEYINPUT115), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT54), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n843), .B2(new_n869), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n833), .A2(new_n841), .A3(new_n831), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n701), .A2(new_n705), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n616), .A2(new_n256), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n721), .A4(new_n766), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n332), .A3(new_n625), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(G952), .A3(new_n254), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n796), .A2(new_n256), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n722), .A3(new_n775), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n784), .A2(new_n755), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT48), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n756), .B2(new_n760), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n889), .B(new_n895), .C1(new_n738), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n823), .A2(new_n824), .ZN(new_n899));
  INV_X1    g713(.A(new_n736), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n720), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n896), .A2(new_n766), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n892), .A2(new_n861), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n332), .A2(new_n625), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n887), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n721), .A2(new_n707), .A3(new_n452), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n897), .A2(KEYINPUT50), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT50), .B1(new_n897), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n903), .B(KEYINPUT51), .C1(new_n904), .C2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n904), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n898), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n903), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n901), .A2(KEYINPUT117), .A3(new_n902), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT51), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n884), .A2(new_n919), .B1(G952), .B2(G953), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n736), .B(KEYINPUT49), .Z(new_n921));
  INV_X1    g735(.A(new_n794), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n755), .A3(new_n452), .A4(new_n720), .ZN(new_n923));
  OR4_X1    g737(.A1(new_n885), .A2(new_n921), .A3(new_n707), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n924), .ZN(G75));
  AOI21_X1  g739(.A(new_n187), .B1(new_n878), .B2(new_n880), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n490), .A2(new_n491), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT119), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n509), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n927), .A2(new_n931), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n254), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G51));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n881), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n342), .B(KEYINPUT57), .Z(new_n938));
  OAI21_X1  g752(.A(new_n734), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n926), .A2(G469), .A3(new_n807), .A4(new_n806), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G54));
  NAND2_X1  g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT120), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n926), .A2(new_n321), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n321), .B1(new_n926), .B2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n934), .ZN(G60));
  OR2_X1    g760(.A1(new_n621), .A2(new_n623), .ZN(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT59), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n884), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n934), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n937), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n950), .A2(new_n953), .ZN(G63));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n881), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n934), .B1(new_n958), .B2(new_n608), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n956), .B1(new_n878), .B2(new_n880), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n960), .A2(KEYINPUT121), .A3(new_n669), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT121), .B1(new_n960), .B2(new_n669), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n959), .B(KEYINPUT61), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n259), .B2(new_n455), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT122), .B1(new_n837), .B2(new_n842), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n970), .B(new_n841), .C1(new_n835), .C2(new_n836), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n972), .B2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n929), .B1(G898), .B2(new_n254), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G69));
  NOR2_X1   g789(.A1(new_n542), .A2(new_n543), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n312), .B(KEYINPUT123), .Z(new_n977));
  XOR2_X1   g791(.A(new_n976), .B(new_n977), .Z(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT124), .Z(new_n979));
  NAND2_X1  g793(.A1(new_n710), .A2(new_n866), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n691), .A2(new_n716), .A3(new_n775), .A4(new_n838), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n829), .A2(new_n817), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n979), .B1(new_n984), .B2(G953), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n865), .A2(new_n764), .A3(new_n790), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n893), .A2(new_n742), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n813), .A3(new_n689), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n817), .A2(new_n986), .A3(new_n786), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n826), .B2(new_n828), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n254), .ZN(new_n991));
  INV_X1    g805(.A(new_n978), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(G953), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n254), .B1(G227), .B2(G900), .ZN(new_n995));
  AOI22_X1  g809(.A1(new_n991), .A2(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n985), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n995), .A2(new_n994), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n984), .B2(new_n972), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n544), .A2(new_n526), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n521), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n871), .A2(new_n876), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n702), .B2(new_n559), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n1003), .A2(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n990), .B1(new_n969), .B2(new_n971), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n1010), .A3(new_n1001), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1004), .A2(new_n521), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n951), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1017), .B(new_n951), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1008), .B1(new_n1016), .B2(new_n1018), .ZN(G57));
endmodule


