//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n461), .A3(G137), .ZN(new_n462));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n468), .B2(G125), .ZN(new_n469));
  AND4_X1   g044(.A1(KEYINPUT68), .A2(new_n459), .A3(new_n461), .A4(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n471), .B2(G2105), .ZN(G160));
  NAND3_X1  g047(.A1(new_n468), .A2(G124), .A3(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n475));
  NOR2_X1   g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n474), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  OAI221_X1 g053(.A(new_n473), .B1(new_n475), .B2(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  NOR2_X1   g055(.A1(new_n458), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G102), .ZN(new_n482));
  NAND2_X1  g057(.A1(G114), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n468), .B2(G126), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(new_n459), .A3(new_n461), .A4(new_n474), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n468), .A2(KEYINPUT4), .A3(new_n474), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n486), .A2(new_n493), .ZN(G164));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(G75), .A2(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT74), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n495), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n511), .A2(G50), .A3(G543), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n505), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n511), .A2(G88), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n516), .B(new_n500), .C1(new_n506), .C2(new_n507), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n509), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n511), .A2(G543), .A3(new_n512), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n522), .A2(new_n525), .A3(new_n526), .A4(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AND3_X1   g107(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(G543), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(new_n500), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(KEYINPUT76), .A3(new_n500), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n511), .A2(G90), .A3(new_n512), .A4(new_n514), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n511), .A2(G52), .A3(G543), .A4(new_n512), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n547), .A2(KEYINPUT77), .A3(new_n540), .A4(new_n541), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  AND2_X1   g124(.A1(new_n521), .A2(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n523), .A2(new_n551), .B1(new_n499), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n535), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n521), .A2(G91), .B1(G651), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n523), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n546), .B2(new_n548), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n546), .A2(new_n548), .A3(new_n571), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G301));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n524), .A2(new_n576), .A3(G49), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n511), .A2(G87), .A3(new_n512), .A4(new_n514), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT80), .B1(new_n523), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n523), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n521), .A2(G86), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n514), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT81), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n500), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n521), .A2(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n524), .A2(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n499), .C2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n535), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n524), .A2(G54), .B1(G651), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n520), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT10), .B1(new_n520), .B2(new_n601), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G301), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(G284));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  XOR2_X1   g185(.A(G299), .B(KEYINPUT82), .Z(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(new_n604), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  INV_X1    g191(.A(new_n554), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n605), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n604), .A2(G559), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT83), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n620), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n468), .A2(new_n481), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n468), .A2(G123), .A3(G2105), .ZN(new_n630));
  NOR2_X1   g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n632));
  INV_X1    g207(.A(G135), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n630), .B1(new_n631), .B2(new_n632), .C1(new_n477), .C2(new_n633), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n634), .A2(G2096), .B1(KEYINPUT85), .B2(new_n626), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n629), .B(new_n635), .C1(G2096), .C2(new_n634), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2435), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2438), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G14), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(KEYINPUT86), .ZN(new_n656));
  OAI21_X1  g231(.A(KEYINPUT17), .B1(new_n656), .B2(new_n651), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(new_n653), .Z(new_n658));
  AND2_X1   g233(.A1(new_n656), .A2(new_n651), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2096), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n626), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n665), .A3(new_n668), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n674), .C1(new_n665), .C2(new_n673), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G1981), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G5), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G171), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G1961), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(KEYINPUT23), .A3(G20), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n689));
  INV_X1    g264(.A(G20), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G299), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n688), .B(new_n691), .C1(new_n692), .C2(new_n683), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT95), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1956), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n683), .A2(G21), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G168), .B2(new_n683), .ZN(new_n697));
  INV_X1    g272(.A(G1966), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G4), .A2(G16), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n614), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT89), .B(G1348), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n685), .A2(G1961), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G35), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G162), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT29), .B(G2090), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G27), .A2(G29), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G164), .B2(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n709), .B1(G2078), .B2(new_n711), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n703), .A2(new_n704), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n695), .A2(new_n699), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT91), .B1(G29), .B2(G33), .ZN(new_n715));
  OR3_X1    g290(.A1(KEYINPUT91), .A2(G29), .A3(G33), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(new_n474), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n481), .A2(G103), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT25), .ZN(new_n720));
  INV_X1    g295(.A(G139), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n477), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n718), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n715), .B(new_n716), .C1(new_n724), .C2(new_n705), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2072), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n705), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G160), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n705), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT30), .B(G28), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n732), .B1(new_n705), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n726), .B(new_n734), .C1(new_n705), .C2(new_n634), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G32), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n481), .A2(G105), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n468), .A2(G2105), .ZN(new_n738));
  INV_X1    g313(.A(G129), .ZN(new_n739));
  INV_X1    g314(.A(G141), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n737), .B1(new_n738), .B2(new_n739), .C1(new_n740), .C2(new_n477), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n736), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G11), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n705), .A2(G26), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n468), .A2(G128), .A3(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n755));
  NOR2_X1   g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT90), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n753), .B1(new_n477), .B2(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(G29), .ZN(new_n759));
  MUX2_X1   g334(.A(new_n752), .B(new_n759), .S(KEYINPUT28), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2067), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n731), .A2(new_n732), .B1(new_n750), .B2(G11), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G2078), .B2(new_n711), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n749), .A2(new_n751), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n714), .A2(new_n735), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n766));
  OR2_X1    g341(.A1(G16), .A2(G23), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G288), .B2(new_n683), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT33), .ZN(new_n769));
  INV_X1    g344(.A(G1976), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(G6), .B(G305), .S(G16), .Z(new_n772));
  XOR2_X1   g347(.A(KEYINPUT32), .B(G1981), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G22), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G166), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT88), .B(G1971), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n771), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT34), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n771), .A2(KEYINPUT34), .A3(new_n774), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n683), .A2(G24), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G290), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1986), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n468), .A2(G119), .A3(G2105), .ZN(new_n789));
  NOR2_X1   g364(.A1(G95), .A2(G2105), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(new_n474), .B2(G107), .ZN(new_n791));
  INV_X1    g366(.A(G131), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n789), .B1(new_n790), .B2(new_n791), .C1(new_n477), .C2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n787), .A2(new_n788), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n766), .B1(new_n783), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n798), .ZN(new_n800));
  AOI211_X1 g375(.A(KEYINPUT36), .B(new_n800), .C1(new_n781), .C2(new_n782), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n687), .B(new_n765), .C1(new_n799), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n683), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n554), .B2(new_n683), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(G311));
  OR2_X1    g381(.A1(new_n799), .A2(new_n801), .ZN(new_n807));
  INV_X1    g382(.A(new_n805), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n807), .A2(new_n687), .A3(new_n765), .A4(new_n808), .ZN(G150));
  XNOR2_X1  g384(.A(KEYINPUT97), .B(G55), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n524), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n520), .A2(new_n812), .B1(new_n499), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NOR2_X1   g393(.A1(new_n604), .A2(new_n615), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT39), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n554), .A2(KEYINPUT98), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n550), .B2(new_n553), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n823), .A3(new_n815), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n617), .A2(new_n816), .A3(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n820), .B(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n818), .B1(new_n829), .B2(G860), .ZN(G145));
  XNOR2_X1  g405(.A(G164), .B(new_n758), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  OR3_X1    g409(.A1(new_n833), .A2(new_n834), .A3(new_n746), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n746), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n723), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n831), .B(new_n745), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n724), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n468), .A2(G130), .A3(G2105), .ZN(new_n841));
  NOR2_X1   g416(.A1(G106), .A2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n843));
  INV_X1    g418(.A(G142), .ZN(new_n844));
  OAI221_X1 g419(.A(new_n841), .B1(new_n842), .B2(new_n843), .C1(new_n477), .C2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n624), .B(new_n845), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n793), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n837), .A2(new_n839), .A3(new_n847), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(KEYINPUT100), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n837), .A2(new_n852), .A3(new_n839), .A4(new_n847), .ZN(new_n853));
  XNOR2_X1  g428(.A(G160), .B(new_n634), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(G37), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n849), .A2(new_n850), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g436(.A1(new_n816), .A2(G868), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n620), .A2(new_n826), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n826), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n614), .A2(new_n692), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n604), .A2(G299), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n863), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n869), .A2(KEYINPUT102), .A3(KEYINPUT41), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(KEYINPUT41), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(KEYINPUT102), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(new_n871), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n869), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n864), .A2(KEYINPUT101), .A3(new_n877), .A4(new_n865), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n870), .A2(new_n876), .A3(new_n881), .A4(new_n878), .ZN(new_n882));
  XOR2_X1   g457(.A(G290), .B(G305), .Z(new_n883));
  XNOR2_X1  g458(.A(G288), .B(G166), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n883), .B(new_n884), .Z(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT42), .Z(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n882), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n862), .B1(new_n889), .B2(G868), .ZN(G295));
  AOI21_X1  g465(.A(new_n862), .B1(new_n889), .B2(G868), .ZN(G331));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  INV_X1    g467(.A(new_n574), .ZN(new_n893));
  OAI21_X1  g468(.A(G168), .B1(new_n893), .B2(new_n572), .ZN(new_n894));
  NAND2_X1  g469(.A1(G171), .A2(G286), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n826), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n826), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n871), .B(new_n875), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n885), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n877), .A3(new_n896), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n900), .B1(new_n899), .B2(new_n902), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n892), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n874), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(new_n872), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n874), .A2(new_n908), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n901), .A2(new_n896), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n902), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n885), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n904), .A3(new_n903), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n907), .B1(new_n915), .B2(new_n892), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT44), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n905), .B2(new_n906), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n903), .A3(new_n892), .A4(new_n904), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(G397));
  XNOR2_X1  g498(.A(KEYINPUT105), .B(G1384), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n486), .B2(new_n493), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n459), .A2(new_n461), .A3(G126), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n483), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G2105), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n482), .A3(new_n491), .A4(new_n492), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n924), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(new_n927), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G40), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n936), .B(new_n464), .C1(new_n471), .C2(G2105), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n939), .A3(new_n745), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n746), .A2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(G2067), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n758), .B(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n938), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n793), .B(new_n796), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n938), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n938), .ZN(new_n951));
  XNOR2_X1  g526(.A(G290), .B(G1986), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n491), .A2(new_n492), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n929), .A2(G2105), .B1(G102), .B2(new_n481), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n937), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(KEYINPUT115), .A3(G8), .ZN(new_n958));
  INV_X1    g533(.A(new_n464), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT68), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n459), .A2(new_n461), .ZN(new_n961));
  INV_X1    g536(.A(G125), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n468), .A2(KEYINPUT68), .A3(G125), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n466), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(G40), .B(new_n959), .C1(new_n965), .C2(new_n474), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n486), .B2(new_n493), .ZN(new_n968));
  OAI21_X1  g543(.A(G8), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n958), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n586), .A2(new_n587), .A3(new_n973), .A4(new_n591), .ZN(new_n974));
  INV_X1    g549(.A(G86), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n591), .B1(new_n520), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(G1981), .B1(new_n976), .B2(new_n585), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT49), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n981), .B1(new_n958), .B2(new_n971), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n982), .A2(G1976), .A3(G288), .ZN(new_n983));
  INV_X1    g558(.A(new_n974), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n972), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n577), .A2(new_n582), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(KEYINPUT116), .A3(G1976), .A4(new_n580), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(G288), .B2(new_n770), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(G288), .B2(new_n770), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n990), .A2(new_n972), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n990), .B2(new_n972), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n992), .A2(new_n994), .A3(new_n982), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n956), .B2(KEYINPUT45), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n968), .A2(KEYINPUT108), .A3(new_n927), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT45), .B(new_n924), .C1(new_n486), .C2(new_n493), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT109), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n931), .A2(new_n1003), .A3(KEYINPUT45), .A4(new_n924), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n999), .A2(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1971), .B1(new_n1005), .B2(new_n937), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n931), .B2(new_n967), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n967), .B(new_n1010), .C1(new_n486), .C2(new_n493), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n937), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT111), .B(G2090), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n997), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n999), .A2(new_n1000), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n937), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1971), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1014), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(KEYINPUT112), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT114), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G303), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(new_n1024), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1030), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1034));
  AOI211_X1 g609(.A(KEYINPUT113), .B(KEYINPUT114), .C1(G303), .C2(G8), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1015), .A2(new_n1022), .A3(new_n1037), .A4(G8), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n985), .B1(new_n996), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n956), .A2(new_n1041), .A3(new_n1007), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT117), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1010), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n968), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n937), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n1013), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1006), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1038), .A2(new_n995), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1011), .A2(G40), .A3(G160), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1052), .A2(G2084), .A3(new_n1008), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n931), .B2(new_n967), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n966), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n968), .A2(new_n927), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n937), .A3(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1053), .B1(new_n1060), .B2(new_n698), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1062), .A3(G286), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1040), .B1(new_n1051), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1015), .A2(new_n1022), .A3(G8), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1040), .B1(new_n1066), .B2(new_n1049), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(new_n1038), .A3(new_n995), .A4(new_n1063), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1039), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G299), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n565), .A2(KEYINPUT57), .A3(new_n568), .A4(new_n569), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1016), .A2(new_n937), .A3(new_n1017), .A4(new_n1074), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT119), .B(G1956), .Z(new_n1076));
  NAND2_X1  g651(.A1(new_n1046), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n702), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1012), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n957), .A2(G2067), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n604), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(new_n1077), .A3(new_n1073), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1016), .A2(new_n939), .A3(new_n937), .A4(new_n1017), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n957), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n554), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT120), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1093), .A3(new_n554), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(KEYINPUT59), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1090), .B2(new_n554), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT120), .B(new_n617), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(KEYINPUT61), .A3(new_n1085), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1075), .A2(new_n1077), .A3(new_n1073), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1078), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1083), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1080), .B(KEYINPUT60), .C1(G2067), .C2(new_n957), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n614), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1086), .B1(new_n1100), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n471), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n467), .B(KEYINPUT122), .C1(new_n469), .C2(new_n470), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(G2105), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(G40), .A4(new_n959), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(new_n934), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G2078), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(G40), .A3(new_n959), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1120), .A2(new_n1017), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G2078), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1016), .A2(new_n1126), .A3(new_n937), .A4(new_n1017), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1121), .ZN(new_n1128));
  INV_X1    g703(.A(G1961), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1012), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .A4(new_n1122), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1135), .A2(G301), .A3(new_n1128), .A4(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1132), .A2(KEYINPUT54), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n1051), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1060), .A2(new_n698), .ZN(new_n1141));
  OAI21_X1  g716(.A(G286), .B1(new_n1141), .B2(new_n1053), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1062), .B1(new_n1061), .B2(G168), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT51), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  AOI211_X1 g720(.A(G286), .B(new_n1053), .C1(new_n1060), .C2(new_n698), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n1062), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1113), .A2(new_n1140), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  AND4_X1   g726(.A1(G301), .A2(new_n1125), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1135), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n607), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1154), .B2(KEYINPUT54), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n607), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT124), .B(new_n1156), .C1(new_n1158), .C2(new_n1152), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1069), .B1(new_n1150), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1148), .A2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1038), .A2(new_n995), .A3(new_n1050), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1144), .A2(KEYINPUT62), .A3(new_n1147), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1158), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1157), .B1(new_n1148), .B2(new_n1162), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1169), .A2(KEYINPUT125), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n953), .B1(new_n1161), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n938), .A2(G1986), .A3(G290), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1174));
  XNOR2_X1  g749(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n793), .A2(new_n795), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n1177), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n758), .A2(G2067), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n938), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n938), .B1(new_n745), .B2(new_n946), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n938), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT46), .B1(new_n938), .B2(G1996), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT47), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1176), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g762(.A(new_n662), .B1(new_n648), .B2(new_n649), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n857), .B2(new_n859), .ZN(new_n1190));
  AND4_X1   g764(.A1(G319), .A2(new_n920), .A3(new_n681), .A4(new_n1190), .ZN(G308));
  NAND4_X1  g765(.A1(new_n920), .A2(new_n1190), .A3(G319), .A4(new_n681), .ZN(G225));
endmodule


