//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT71), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT71), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT72), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n473), .A2(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT73), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n464), .A2(new_n466), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n462), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT74), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n477), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n492), .B2(G136), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n467), .B2(new_n468), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n476), .A2(KEYINPUT75), .A3(G126), .A4(G2105), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT76), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT7), .Z(new_n530));
  INV_X1    g105(.A(new_n519), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n516), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n519), .A2(new_n537), .B1(new_n521), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n516), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n519), .A2(new_n543), .B1(new_n521), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n521), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n521), .B2(new_n554), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(new_n556), .B1(G91), .B2(new_n531), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n511), .A2(new_n513), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n516), .B1(new_n561), .B2(KEYINPUT78), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(KEYINPUT78), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n557), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  XNOR2_X1  g140(.A(G166), .B(KEYINPUT79), .ZN(G303));
  INV_X1    g141(.A(G74), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n516), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT80), .ZN(new_n569));
  INV_X1    g144(.A(new_n521), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n531), .A2(G87), .B1(G49), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G288));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT81), .B1(new_n559), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G73), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n510), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n559), .A2(KEYINPUT81), .A3(new_n573), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n531), .A2(G86), .B1(G48), .B2(new_n570), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n516), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n519), .A2(new_n583), .B1(new_n521), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n582), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n531), .A2(G92), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT84), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(KEYINPUT86), .B(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n559), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n588), .A2(new_n590), .B1(G651), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n521), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n521), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n591), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n587), .B1(new_n601), .B2(G868), .ZN(new_n602));
  MUX2_X1   g177(.A(new_n587), .B(new_n602), .S(KEYINPUT82), .Z(G284));
  MUX2_X1   g178(.A(new_n587), .B(new_n602), .S(KEYINPUT82), .Z(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n601), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n465), .A2(G2104), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT71), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT72), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n472), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n484), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n462), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G135), .B2(new_n492), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT88), .Z(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT89), .B(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n635), .ZN(G156));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT16), .B(G1341), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n642), .A2(new_n648), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(KEYINPUT17), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n658), .B(new_n660), .C1(new_n661), .C2(new_n657), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n660), .A2(KEYINPUT18), .A3(new_n656), .ZN(new_n663));
  OAI21_X1  g238(.A(KEYINPUT18), .B1(new_n660), .B2(new_n656), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n670), .A2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n674), .B(new_n676), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1991), .ZN(new_n682));
  INV_X1    g257(.A(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G4), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n601), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT93), .B(G1348), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  NOR2_X1   g268(.A1(G29), .A2(G32), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n622), .A2(G105), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT26), .Z(new_n699));
  INV_X1    g274(.A(G129), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n485), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n492), .A2(G141), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n694), .B1(new_n707), .B2(G29), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT27), .B(G1996), .Z(new_n709));
  AOI21_X1  g284(.A(new_n693), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(G164), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G27), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G2078), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n689), .A2(G19), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n546), .B2(new_n689), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT94), .B(G1341), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G5), .A2(G16), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G301), .B2(new_n689), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n720), .B1(G1961), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n711), .A2(new_n716), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n710), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n712), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n712), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2090), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n689), .A2(G20), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G299), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1956), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT103), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n712), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n484), .A2(G128), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n743), .A2(G104), .A3(G2105), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(G104), .B2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n742), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n492), .B2(G140), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(new_n712), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n715), .B2(new_n714), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n712), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n492), .A2(G139), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n620), .A2(G127), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n462), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(new_n712), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n730), .A2(G2090), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT101), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n751), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  OR2_X1    g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NAND2_X1  g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G160), .B2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n727), .A2(new_n738), .A3(new_n767), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n633), .A2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n712), .B1(new_n778), .B2(G28), .ZN(new_n780));
  INV_X1    g355(.A(G1961), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n777), .B1(new_n779), .B2(new_n780), .C1(new_n723), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n689), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n689), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n782), .B1(G1966), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n776), .B(new_n785), .C1(G1966), .C2(new_n784), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT100), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n774), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT92), .B1(new_n689), .B2(G22), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n689), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n689), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n796), .B1(new_n798), .B2(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n794), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT32), .B(G1981), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n799), .A2(new_n795), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n809));
  INV_X1    g384(.A(G119), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n485), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n484), .A2(KEYINPUT91), .A3(G119), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n462), .A2(G107), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n492), .A2(G131), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G25), .B(new_n817), .S(G29), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G24), .B(G290), .S(G16), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1986), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n808), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n808), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n789), .A2(new_n829), .ZN(G311));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n789), .B2(new_n829), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n788), .A2(new_n828), .A3(KEYINPUT104), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(G150));
  NOR2_X1   g409(.A1(new_n600), .A2(new_n609), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n531), .A2(G93), .B1(G55), .B2(new_n570), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n516), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n546), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(new_n841), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n817), .B(new_n748), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n624), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n706), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n760), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n706), .B(new_n624), .ZN(new_n854));
  INV_X1    g429(.A(new_n760), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n492), .A2(G142), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n484), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n462), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n495), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n618), .B2(new_n619), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT105), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n496), .B2(new_n498), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n507), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n861), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n853), .A2(new_n856), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n853), .B2(new_n856), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n850), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n854), .A2(new_n855), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n852), .A2(new_n760), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(new_n849), .A3(new_n871), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n633), .B(G160), .Z(new_n880));
  INV_X1    g455(.A(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT106), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  AOI211_X1 g460(.A(new_n885), .B(new_n882), .C1(new_n874), .C2(new_n878), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n848), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n874), .A2(new_n878), .A3(new_n882), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n874), .A2(new_n878), .A3(KEYINPUT107), .A4(new_n882), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT40), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n872), .A2(new_n850), .A3(new_n873), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n849), .B1(new_n877), .B2(new_n871), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n883), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n885), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n879), .A2(KEYINPUT106), .A3(new_n883), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n900), .A2(new_n892), .A3(new_n901), .A4(new_n848), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n894), .A2(new_n902), .ZN(G395));
  NAND2_X1  g478(.A1(new_n840), .A2(new_n605), .ZN(new_n904));
  XNOR2_X1  g479(.A(G290), .B(G288), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n905), .A2(KEYINPUT110), .ZN(new_n906));
  XOR2_X1   g481(.A(G305), .B(G166), .Z(new_n907));
  OR2_X1    g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(KEYINPUT110), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT111), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT42), .Z(new_n914));
  OR2_X1    g489(.A1(G299), .A2(KEYINPUT108), .ZN(new_n915));
  NAND2_X1  g490(.A1(G299), .A2(KEYINPUT108), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n601), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n600), .A2(G299), .A3(KEYINPUT108), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT109), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n919), .B2(KEYINPUT41), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n611), .B(new_n841), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n919), .B(new_n926), .S(new_n927), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n914), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n904), .B1(new_n929), .B2(new_n605), .ZN(G295));
  OAI21_X1  g505(.A(new_n904), .B1(new_n929), .B2(new_n605), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  NOR2_X1   g507(.A1(G286), .A2(G171), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n841), .ZN(new_n935));
  NAND2_X1  g510(.A1(G286), .A2(G171), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n841), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n919), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n920), .A2(new_n922), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n848), .B1(new_n944), .B2(new_n911), .ZN(new_n945));
  INV_X1    g520(.A(new_n940), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n923), .B2(new_n925), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n947), .A2(new_n912), .A3(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT112), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n941), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n911), .B(new_n950), .C1(new_n926), .C2(new_n946), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n942), .B2(new_n946), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n952), .B2(new_n912), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n932), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n912), .B1(new_n947), .B2(new_n941), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n848), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n958), .A2(new_n932), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT44), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n953), .A3(new_n932), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n505), .A2(new_n506), .ZN(new_n968));
  INV_X1    g543(.A(new_n502), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n863), .B2(new_n864), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n496), .A2(new_n866), .A3(new_n498), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n973), .B2(G1384), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n471), .A2(new_n976), .A3(new_n478), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT115), .ZN(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n748), .B(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(G1996), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n707), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n979), .A2(new_n981), .B1(new_n983), .B2(KEYINPUT114), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n706), .ZN(new_n985));
  OAI221_X1 g560(.A(new_n984), .B1(KEYINPUT114), .B2(new_n983), .C1(new_n683), .C2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n817), .B(new_n819), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n979), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n990));
  INV_X1    g565(.A(new_n978), .ZN(new_n991));
  AND2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT113), .Z(new_n994));
  NOR2_X1   g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G303), .A2(G8), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT55), .Z(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n973), .A2(new_n967), .A3(G1384), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n499), .B2(new_n507), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n977), .B1(KEYINPUT45), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT116), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n868), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(G101), .A2(new_n622), .B1(new_n488), .B2(G137), .ZN(new_n1005));
  INV_X1    g580(.A(new_n470), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n620), .B2(G125), .ZN(new_n1007));
  OAI211_X1 g582(.A(G40), .B(new_n1005), .C1(new_n1007), .C2(new_n462), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n508), .A2(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n967), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1971), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT50), .B1(new_n973), .B2(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n508), .A2(new_n1015), .A3(new_n1003), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1000), .A2(KEYINPUT119), .A3(new_n1015), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1014), .A2(new_n1018), .A3(new_n977), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT120), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G2090), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1013), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n998), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n868), .A2(new_n977), .A3(new_n1003), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1027), .B2(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n578), .A2(new_n1034), .A3(new_n579), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n1030), .A2(new_n1031), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1031), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1029), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n791), .B2(G1976), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1041), .B(new_n1046), .C1(new_n1042), .C2(new_n1029), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1012), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1011), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n795), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1008), .B1(new_n1009), .B2(KEYINPUT50), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n868), .A2(new_n1003), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(KEYINPUT50), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G2090), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n1013), .B2(new_n1056), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(G8), .A4(new_n997), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1002), .A2(new_n1012), .A3(new_n715), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1061), .A2(new_n1062), .B1(new_n781), .B2(new_n1055), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1000), .A2(KEYINPUT45), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(G2078), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n974), .A2(new_n1064), .A3(new_n977), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G301), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  AND4_X1   g642(.A1(new_n1026), .A2(new_n1048), .A3(new_n1060), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n974), .A2(new_n1064), .A3(new_n977), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1053), .B(new_n772), .C1(new_n1054), .C2(KEYINPUT50), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(G8), .A3(G286), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(G168), .A3(new_n1073), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT126), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT126), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1069), .B(new_n1075), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1068), .A2(new_n1083), .A3(KEYINPUT127), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT127), .B1(new_n1068), .B2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1086), .A2(KEYINPUT62), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1039), .A2(new_n1040), .A3(new_n791), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1035), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1060), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1058), .A2(new_n1059), .A3(G8), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n998), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1074), .A2(G8), .A3(G168), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT121), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1095), .A2(new_n1097), .A3(new_n1060), .A4(new_n1048), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(KEYINPUT63), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(G171), .B(KEYINPUT54), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1004), .A2(new_n974), .A3(new_n977), .A4(new_n1065), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1063), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1055), .A2(new_n781), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1066), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n973), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n479), .B(G40), .C1(new_n1000), .C2(new_n1015), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n692), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n977), .A3(new_n1003), .A4(new_n980), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT123), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n973), .A2(G1384), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n980), .A4(new_n977), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1111), .A2(new_n601), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1004), .A2(new_n1010), .A3(new_n683), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1027), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n546), .A2(KEYINPUT125), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT59), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n1123), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1118), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  INV_X1    g704(.A(G1956), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1020), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(G299), .B(KEYINPUT57), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(new_n762), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1004), .A2(new_n1010), .A3(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1131), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1133), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1129), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1132), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1131), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1111), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n600), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1117), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1128), .A2(new_n1139), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n601), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1144), .A2(KEYINPUT124), .A3(new_n601), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1141), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1142), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1108), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1101), .B1(new_n1154), .B2(new_n1086), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1026), .A2(new_n1048), .A3(new_n1060), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1099), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n995), .B1(new_n1088), .B2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n982), .B(KEYINPUT46), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n979), .A2(new_n981), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n985), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT47), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n990), .B(KEYINPUT48), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n989), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n748), .A2(new_n980), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n817), .A2(new_n819), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n986), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1164), .B1(new_n979), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g744(.A1(new_n900), .A2(new_n848), .A3(new_n892), .ZN(new_n1171));
  OAI211_X1 g745(.A(G319), .B(new_n667), .C1(new_n650), .C2(new_n649), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G229), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1171), .A2(new_n963), .A3(new_n1173), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n963), .A3(new_n1173), .ZN(G225));
endmodule


