//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT69), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(new_n187), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT69), .B(G128), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT95), .B1(new_n196), .B2(G143), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n188), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n188), .C1(new_n195), .C2(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n203));
  INV_X1    g017(.A(G122), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G116), .ZN(new_n205));
  INV_X1    g019(.A(G116), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT94), .A3(G122), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n205), .A2(new_n207), .B1(G116), .B2(new_n204), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G116), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(KEYINPUT14), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n208), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n202), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT9), .B(G234), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(G217), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT96), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT13), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n188), .B(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n194), .B1(new_n193), .B2(new_n187), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n196), .A2(KEYINPUT95), .A3(G143), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n219), .B1(new_n224), .B2(new_n200), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n195), .A2(new_n197), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT96), .B(G134), .C1(new_n226), .C2(new_n221), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n208), .B(new_n209), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n201), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n213), .B(new_n218), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n225), .B2(new_n227), .ZN(new_n232));
  INV_X1    g046(.A(new_n212), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n199), .B2(new_n201), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n217), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G478), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(G902), .B1(new_n231), .B2(new_n235), .ZN(new_n242));
  INV_X1    g056(.A(new_n240), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G234), .ZN(new_n246));
  INV_X1    g060(.A(G237), .ZN(new_n247));
  OAI211_X1 g061(.A(G952), .B(new_n216), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(new_n248), .B(KEYINPUT97), .Z(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT71), .A2(G953), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT71), .A2(G953), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI211_X1 g067(.A(new_n237), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT21), .B(G898), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT98), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n250), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n245), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n216), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT71), .A2(G953), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(G214), .A3(new_n247), .A4(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(new_n187), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n187), .ZN(new_n265));
  OAI21_X1  g079(.A(G131), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n187), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n253), .A2(G143), .A3(G214), .A4(new_n247), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT92), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n266), .A2(new_n274), .A3(new_n267), .A4(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(G140), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G125), .ZN(new_n277));
  INV_X1    g091(.A(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G140), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT79), .A4(KEYINPUT16), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT16), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n277), .B2(KEYINPUT16), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G146), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT16), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n278), .A2(KEYINPUT16), .A3(G140), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n282), .ZN(new_n288));
  INV_X1    g102(.A(G146), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n280), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n267), .B(new_n270), .C1(new_n268), .C2(new_n269), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n273), .A2(new_n275), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(G113), .B(G122), .ZN(new_n295));
  INV_X1    g109(.A(G104), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n268), .A2(new_n269), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT87), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT87), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n268), .A2(new_n269), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(KEYINPUT18), .A2(G131), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n268), .A2(new_n269), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n302), .B(KEYINPUT89), .Z(new_n306));
  AOI21_X1  g120(.A(new_n289), .B1(new_n277), .B2(new_n279), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT88), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n277), .A2(new_n279), .A3(new_n289), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT88), .B1(new_n312), .B2(new_n307), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n305), .A2(new_n306), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n294), .A2(new_n297), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n266), .A2(new_n271), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n289), .B1(new_n288), .B2(new_n280), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT90), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n277), .A2(new_n279), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT19), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n277), .A2(new_n279), .A3(new_n319), .A4(KEYINPUT19), .ZN(new_n323));
  AOI21_X1  g137(.A(G146), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n304), .A2(new_n314), .B1(new_n317), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n324), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n329), .B(new_n285), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n268), .A2(new_n269), .A3(new_n300), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n300), .B1(new_n268), .B2(new_n269), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n333), .A2(new_n334), .A3(new_n302), .ZN(new_n335));
  INV_X1    g149(.A(new_n311), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n337));
  INV_X1    g151(.A(new_n306), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n336), .A2(new_n337), .B1(new_n298), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n327), .B(new_n332), .C1(new_n335), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n297), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n316), .B1(new_n328), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n344));
  NOR2_X1   g158(.A1(G475), .A2(G902), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT93), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n343), .A2(new_n348), .A3(new_n344), .A4(new_n345), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n335), .A2(new_n339), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT17), .B(G131), .C1(new_n264), .C2(new_n265), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n290), .A3(new_n285), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(KEYINPUT92), .B2(new_n272), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n353), .B2(new_n275), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n297), .B1(new_n326), .B2(new_n327), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n315), .A2(new_n332), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT91), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n297), .A2(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n345), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n349), .A3(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n354), .A2(new_n297), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n316), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n237), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G475), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n259), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT99), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT99), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n259), .A2(new_n361), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  INV_X1    g185(.A(G119), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G116), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n206), .A2(G119), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT2), .B(G113), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT11), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n200), .B2(G137), .ZN(new_n383));
  INV_X1    g197(.A(G137), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT11), .A3(G134), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n200), .A2(G137), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G131), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT65), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(new_n385), .A3(new_n270), .A4(new_n386), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(KEYINPUT65), .A3(G131), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT64), .B1(new_n187), .B2(G146), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT64), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n289), .A3(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n187), .A2(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(KEYINPUT0), .A2(G128), .ZN(new_n398));
  NOR2_X1   g212(.A1(KEYINPUT0), .A2(G128), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G143), .B(G146), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n397), .A2(new_n400), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n391), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G134), .B(G137), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT66), .B1(new_n404), .B2(new_n270), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n200), .A2(G137), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n384), .A2(G134), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n406), .B(G131), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n390), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n289), .A2(G143), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n396), .A3(G128), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT67), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT67), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT1), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n411), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n401), .A2(new_n420), .A3(KEYINPUT68), .A4(G128), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n412), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n193), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n397), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n410), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n403), .A2(new_n426), .A3(KEYINPUT30), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n425), .ZN(new_n429));
  INV_X1    g243(.A(new_n410), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n391), .A2(new_n392), .A3(new_n402), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n381), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n253), .A2(G210), .A3(new_n247), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT27), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT26), .B(G101), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT70), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n381), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n379), .A2(KEYINPUT70), .A3(new_n380), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n431), .A3(new_n432), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n434), .A2(new_n438), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n381), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT30), .B1(new_n403), .B2(new_n426), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n431), .A2(new_n428), .A3(new_n432), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n438), .ZN(new_n450));
  INV_X1    g264(.A(new_n443), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT31), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n445), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n419), .A2(new_n421), .B1(new_n424), .B2(new_n397), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n432), .B1(new_n455), .B2(new_n410), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT73), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n431), .A2(new_n458), .A3(new_n432), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n442), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT28), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n381), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n443), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT28), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n438), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT32), .B(new_n371), .C1(new_n454), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT75), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n441), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT70), .B1(new_n379), .B2(new_n380), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n456), .B2(KEYINPUT73), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT28), .B1(new_n473), .B2(new_n459), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n461), .B1(new_n463), .B2(new_n443), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n450), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n476), .B(new_n445), .C1(new_n453), .C2(new_n452), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n371), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n371), .B1(new_n454), .B2(new_n466), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT74), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n462), .A2(new_n438), .A3(new_n465), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n472), .B1(new_n403), .B2(new_n426), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n461), .B1(new_n488), .B2(new_n443), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n461), .B2(new_n460), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n450), .A2(new_n485), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G472), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT74), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n495), .A3(new_n481), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n479), .A2(new_n483), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n372), .A2(G128), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n372), .A2(G128), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n196), .A2(G119), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT23), .ZN(new_n502));
  OAI221_X1 g316(.A(new_n498), .B1(new_n499), .B2(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(G110), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT77), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n501), .A2(new_n505), .A3(new_n498), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n501), .B2(new_n498), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  NOR3_X1   g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n285), .B(new_n310), .C1(new_n504), .C2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n506), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n503), .A2(G110), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n291), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n513), .A3(new_n517), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n237), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G217), .B1(new_n246), .B2(G902), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT76), .ZN(new_n525));
  INV_X1    g339(.A(new_n520), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n517), .B1(new_n510), .B2(new_n513), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n525), .A2(G902), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n523), .A2(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G221), .B1(new_n214), .B2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G469), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n237), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT10), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n401), .A2(G128), .B1(new_n414), .B2(new_n396), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n419), .B2(new_n421), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n296), .A2(G107), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n296), .A2(G107), .ZN(new_n540));
  OAI21_X1  g354(.A(G101), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT3), .B1(new_n296), .B2(G107), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT3), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n209), .A3(G104), .ZN(new_n544));
  INV_X1    g358(.A(G101), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n538), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n535), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n535), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n429), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n542), .A2(new_n544), .A3(new_n538), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G101), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT4), .A3(new_n546), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT4), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n554), .A3(G101), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n402), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n391), .A2(new_n392), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n548), .A2(new_n550), .A3(new_n558), .A4(new_n556), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n253), .A2(G227), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT80), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G140), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n422), .A2(new_n425), .A3(new_n547), .ZN(new_n569));
  INV_X1    g383(.A(new_n536), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n547), .B1(new_n422), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n559), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n559), .B(new_n575), .C1(new_n569), .C2(new_n571), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n574), .A2(new_n561), .A3(new_n566), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n534), .B1(new_n578), .B2(new_n533), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n561), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n567), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(G469), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n532), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n402), .A2(new_n278), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n422), .A2(new_n278), .A3(new_n425), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G224), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT84), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n587), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(G110), .B(G122), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n553), .A2(new_n381), .A3(new_n555), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT5), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n372), .A3(G116), .ZN(new_n595));
  OAI211_X1 g409(.A(G113), .B(new_n595), .C1(new_n375), .C2(new_n594), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n379), .A2(new_n596), .A3(new_n546), .A4(new_n541), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n592), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n593), .A2(new_n592), .A3(new_n597), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT6), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT6), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n598), .A2(KEYINPUT83), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT83), .B1(new_n598), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n591), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n402), .A2(new_n278), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n455), .B2(new_n278), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT85), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT85), .ZN(new_n611));
  INV_X1    g425(.A(new_n609), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n587), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT86), .B1(new_n587), .B2(new_n612), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT86), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n607), .A2(new_n616), .A3(new_n609), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n592), .B(KEYINPUT8), .ZN(new_n619));
  INV_X1    g433(.A(new_n597), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n379), .A2(new_n596), .B1(new_n546), .B2(new_n541), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n600), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n614), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n605), .A2(new_n237), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G210), .B1(G237), .B2(G902), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n623), .B1(new_n610), .B2(new_n613), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n630), .B2(new_n618), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n627), .A3(new_n605), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(G214), .B1(G237), .B2(G902), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT82), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n584), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n370), .A2(new_n497), .A3(new_n530), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  NAND2_X1  g453(.A1(new_n477), .A2(new_n237), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n530), .A2(new_n480), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n579), .A2(new_n583), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n531), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n361), .A2(new_n365), .ZN(new_n646));
  INV_X1    g460(.A(new_n634), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n258), .B(new_n647), .C1(new_n629), .C2(new_n632), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n235), .A2(KEYINPUT100), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n236), .A2(new_n649), .A3(KEYINPUT33), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n231), .B(new_n235), .C1(KEYINPUT100), .C2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(G478), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n239), .A2(new_n237), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n242), .B2(new_n239), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n646), .A2(new_n648), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n645), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n360), .A2(KEYINPUT101), .A3(new_n346), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n365), .A2(new_n648), .A3(new_n668), .A4(new_n245), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n645), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NAND2_X1  g487(.A1(new_n641), .A2(new_n480), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n518), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n514), .B(new_n675), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n523), .A2(new_n525), .B1(new_n529), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n370), .A2(new_n637), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n250), .B1(new_n254), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n365), .A2(new_n668), .A3(new_n245), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n632), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n627), .B1(new_n631), .B2(new_n605), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n634), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n644), .A2(new_n677), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n497), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XOR2_X1   g505(.A(new_n683), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n584), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT40), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n633), .B(KEYINPUT38), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n634), .A3(new_n677), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n646), .A2(new_n245), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n450), .B1(new_n434), .B2(new_n443), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n488), .A2(new_n443), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n237), .B1(new_n700), .B2(new_n438), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n479), .A2(new_n483), .A3(new_n496), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n694), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  AOI211_X1 g519(.A(new_n683), .B(new_n656), .C1(new_n361), .C2(new_n365), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n497), .A2(new_n689), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  OR2_X1    g522(.A1(new_n578), .A2(new_n533), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n578), .A2(new_n533), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n531), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n497), .A2(new_n658), .A3(new_n530), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n669), .A2(new_n497), .A3(new_n530), .A4(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AOI21_X1  g531(.A(KEYINPUT25), .B1(new_n528), .B2(new_n237), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n521), .A2(new_n522), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n525), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n676), .A2(new_n529), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n711), .B2(new_n688), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n578), .B(G469), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n647), .B1(new_n629), .B2(new_n632), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT102), .A4(new_n531), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n370), .A2(new_n497), .A3(new_n722), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n646), .B2(new_n245), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n241), .A2(new_n244), .ZN(new_n733));
  AOI211_X1 g547(.A(KEYINPUT103), .B(new_n733), .C1(new_n361), .C2(new_n365), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n490), .A2(new_n438), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n371), .B1(new_n454), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n530), .A2(new_n641), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n258), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n726), .A3(new_n739), .A4(new_n531), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  AND3_X1   g557(.A1(new_n722), .A2(new_n641), .A3(new_n737), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n728), .A2(new_n744), .A3(new_n706), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NAND2_X1  g560(.A1(new_n581), .A2(new_n582), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT104), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n582), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(G469), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n532), .B1(new_n751), .B2(new_n579), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT105), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n629), .A2(new_n755), .A3(new_n632), .A4(new_n634), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n528), .ZN(new_n758));
  INV_X1    g572(.A(new_n529), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n720), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n481), .A2(new_n480), .B1(new_n493), .B2(G472), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n467), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n762), .A3(new_n706), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT42), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n766), .A2(new_n646), .A3(new_n657), .A4(new_n684), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n497), .A3(new_n530), .A4(new_n757), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n764), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n764), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND4_X1  g586(.A1(new_n685), .A2(new_n497), .A3(new_n530), .A4(new_n757), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NAND3_X1  g588(.A1(new_n748), .A2(KEYINPUT45), .A3(new_n750), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n533), .B1(new_n747), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n534), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n534), .B1(new_n775), .B2(new_n777), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n710), .A4(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(new_n531), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n692), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n657), .A2(new_n361), .A3(new_n365), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n789), .B2(new_n792), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n674), .A3(new_n722), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n788), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n754), .A2(new_n756), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n795), .B2(new_n796), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(KEYINPUT109), .B(G137), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(G39));
  NAND3_X1  g618(.A1(new_n706), .A2(new_n799), .A3(new_n760), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n497), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n738), .A2(new_n249), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n794), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n808), .A2(new_n809), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n725), .A2(new_n532), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n800), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n799), .A2(new_n712), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n249), .B1(new_n818), .B2(KEYINPUT115), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n703), .A2(new_n760), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n646), .A2(new_n657), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n744), .A3(new_n794), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n647), .B1(KEYINPUT114), .B2(KEYINPUT50), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n695), .A2(new_n711), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n794), .A2(new_n813), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT114), .B1(KEYINPUT113), .B2(KEYINPUT50), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n824), .A2(new_n825), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n812), .B1(new_n817), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n812), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n815), .A2(KEYINPUT116), .A3(new_n816), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n814), .A2(new_n800), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n815), .B2(new_n816), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n821), .A2(new_n762), .A3(new_n794), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT48), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n216), .A2(G952), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n814), .B1(new_n724), .B2(new_n727), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n821), .A2(new_n822), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n646), .A2(new_n657), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n834), .A2(new_n840), .A3(new_n842), .A4(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n690), .A2(new_n745), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n752), .A2(new_n677), .A3(new_n684), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n735), .A2(new_n726), .A3(new_n703), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n707), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n690), .A2(new_n745), .A3(new_n707), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n646), .A2(new_n731), .A3(new_n245), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n726), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n703), .A2(new_n851), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n854), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n757), .A2(new_n706), .A3(new_n744), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n241), .A2(new_n244), .A3(new_n684), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n664), .A2(new_n665), .A3(new_n663), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT101), .B1(new_n360), .B2(new_n346), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n365), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n668), .A2(KEYINPUT110), .A3(new_n365), .A4(new_n865), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n754), .A2(new_n584), .A3(new_n756), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n497), .A2(new_n722), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n863), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n773), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT111), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n754), .A2(new_n584), .A3(new_n756), .ZN(new_n878));
  INV_X1    g692(.A(G475), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n363), .B2(new_n237), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n864), .B(new_n880), .C1(new_n666), .C2(new_n667), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n881), .B2(KEYINPUT110), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n497), .A3(new_n722), .A4(new_n870), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT111), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n773), .A4(new_n863), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n642), .A2(new_n636), .A3(new_n258), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n846), .B1(new_n646), .B2(new_n733), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n638), .A2(new_n742), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n729), .A2(new_n679), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n716), .A2(new_n713), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n862), .A2(new_n886), .A3(new_n771), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT53), .ZN(new_n895));
  INV_X1    g709(.A(new_n892), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n497), .A2(new_n722), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n367), .A2(new_n369), .B1(new_n724), .B2(new_n727), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n636), .B1(new_n367), .B2(new_n369), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n897), .A2(new_n898), .B1(new_n899), .B2(new_n678), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n735), .A2(new_n741), .B1(new_n887), .B2(new_n888), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n896), .A2(new_n900), .A3(new_n638), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n877), .B2(new_n885), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n771), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n853), .A2(new_n861), .A3(KEYINPUT112), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT112), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n907), .B(new_n854), .C1(new_n855), .C2(new_n860), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n895), .B(KEYINPUT54), .C1(new_n905), .C2(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n768), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n903), .A2(new_n908), .A3(new_n906), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n894), .A2(new_n904), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n910), .B1(KEYINPUT54), .B2(new_n914), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n849), .A2(new_n915), .B1(G952), .B2(G953), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n530), .A2(new_n531), .A3(new_n635), .ZN(new_n917));
  INV_X1    g731(.A(new_n725), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT49), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n657), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(KEYINPUT49), .ZN(new_n921));
  OR4_X1    g735(.A1(new_n646), .A2(new_n920), .A3(new_n695), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n916), .B1(new_n703), .B2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n253), .A2(G952), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT118), .Z(new_n925));
  AOI21_X1  g739(.A(new_n237), .B1(new_n912), .B2(new_n913), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n591), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n925), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n906), .A2(new_n908), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n886), .A2(new_n893), .A3(new_n911), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n932), .A2(new_n933), .B1(new_n894), .B2(new_n904), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT117), .B1(new_n934), .B2(new_n237), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n894), .A2(new_n904), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n886), .A2(new_n893), .A3(new_n911), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n909), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n936), .B(G902), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n935), .A2(new_n940), .A3(new_n628), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n930), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n931), .B1(new_n941), .B2(new_n943), .ZN(G51));
  XNOR2_X1  g758(.A(new_n534), .B(KEYINPUT57), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n934), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n568), .A2(new_n577), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n778), .B(KEYINPUT119), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n935), .A2(new_n940), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n924), .B1(new_n951), .B2(new_n953), .ZN(G54));
  AND3_X1   g768(.A1(new_n343), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n935), .A2(new_n940), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n924), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n935), .A2(new_n940), .A3(KEYINPUT58), .A4(G475), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n358), .B2(new_n959), .ZN(G60));
  NOR2_X1   g774(.A1(new_n946), .A2(new_n948), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n650), .A2(new_n652), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n654), .B(KEYINPUT121), .ZN(new_n963));
  XOR2_X1   g777(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n925), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n962), .B1(new_n915), .B2(new_n965), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(G63));
  INV_X1    g783(.A(new_n925), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n914), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n974), .B2(new_n758), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n676), .B(KEYINPUT122), .Z(new_n976));
  OAI211_X1 g790(.A(new_n975), .B(KEYINPUT61), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n934), .A2(new_n972), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n925), .B1(new_n979), .B2(new_n528), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n974), .A2(new_n976), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n977), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n257), .B2(new_n588), .ZN(new_n984));
  INV_X1    g798(.A(new_n253), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n893), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n928), .B1(G898), .B2(new_n253), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NOR2_X1   g802(.A1(new_n427), .A2(new_n433), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n322), .A2(new_n323), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n855), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n704), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n800), .A2(new_n693), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(new_n497), .A3(new_n530), .A4(new_n888), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n810), .A2(new_n802), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n998), .A2(KEYINPUT123), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(KEYINPUT123), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n991), .B1(new_n1001), .B2(new_n985), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n991), .B1(G900), .B2(new_n985), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n810), .A2(new_n992), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n735), .A2(new_n726), .A3(new_n762), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n773), .B1(new_n788), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n798), .B2(new_n801), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1004), .A2(new_n771), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1003), .B1(new_n1008), .B2(new_n985), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n991), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT125), .Z(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1002), .A2(new_n1009), .A3(new_n1014), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G72));
  XNOR2_X1  g832(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1022), .B1(new_n1008), .B2(new_n902), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n449), .A2(new_n438), .A3(new_n451), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n924), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n699), .A2(new_n1024), .A3(new_n1021), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n895), .B(new_n1026), .C1(new_n905), .C2(new_n909), .ZN(new_n1027));
  NOR4_X1   g841(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n902), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n699), .B1(new_n1028), .B2(new_n1021), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .ZN(G57));
endmodule


