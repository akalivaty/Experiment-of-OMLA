//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT12), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT64), .A3(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n201), .B2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G104), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n202), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n201), .A2(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n204), .A2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(G101), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n198), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT67), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n194), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n197), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n200), .B(new_n212), .C1(new_n215), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n193), .A2(new_n195), .B1(G143), .B2(new_n192), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n200), .B1(new_n224), .B2(new_n213), .ZN(new_n225));
  INV_X1    g039(.A(new_n212), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT76), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n223), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(new_n233), .C1(new_n234), .C2(G137), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT66), .A2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT66), .A2(G137), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n235), .A2(new_n238), .A3(new_n242), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n189), .B(new_n190), .C1(new_n231), .C2(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n225), .A2(new_n229), .A3(new_n226), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n229), .B1(new_n225), .B2(new_n226), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n222), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT12), .A3(new_n244), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n244), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n189), .B1(new_n252), .B2(new_n190), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n200), .B1(new_n215), .B2(new_n221), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT10), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n212), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT0), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n198), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  OR3_X1    g075(.A1(new_n214), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n224), .A2(new_n260), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G101), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n267), .A2(KEYINPUT4), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n258), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n228), .A2(new_n230), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n256), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n273), .B(new_n256), .C1(new_n247), .C2(new_n248), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n245), .B(new_n272), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  INV_X1    g093(.A(G227), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n279), .B(new_n281), .Z(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n254), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n272), .B1(new_n275), .B2(new_n277), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n244), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n282), .B1(new_n286), .B2(new_n278), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n188), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n278), .B1(new_n251), .B2(new_n253), .ZN(new_n290));
  INV_X1    g104(.A(new_n282), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n256), .B1(new_n247), .B2(new_n248), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT77), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n271), .B1(new_n293), .B2(new_n276), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n294), .B2(new_n245), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n290), .A2(new_n291), .B1(new_n295), .B2(new_n286), .ZN(new_n296));
  OAI21_X1  g110(.A(G469), .B1(new_n296), .B2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT79), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(G469), .C1(new_n296), .C2(G902), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n289), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT69), .A2(G116), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(G122), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT90), .B1(new_n303), .B2(G122), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n309));
  INV_X1    g123(.A(G122), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G107), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n306), .A3(new_n204), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n198), .A2(G143), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n194), .A2(G128), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(new_n234), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n198), .B2(G143), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT91), .B1(new_n324), .B2(new_n317), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n194), .A2(G128), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(new_n318), .C2(new_n323), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G134), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(KEYINPUT92), .A3(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n312), .A2(new_n306), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G107), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n337), .A2(new_n316), .B1(new_n234), .B2(new_n319), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n322), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n330), .A2(KEYINPUT92), .A3(G134), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT92), .B1(new_n330), .B2(G134), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n322), .B(new_n338), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n321), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT9), .B(G234), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n345), .A2(new_n346), .A3(G953), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n321), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT93), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n349), .B1(new_n351), .B2(new_n342), .ZN(new_n352));
  INV_X1    g166(.A(new_n347), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n188), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT94), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT94), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n348), .A2(new_n354), .A3(new_n357), .A4(new_n188), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT15), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G478), .ZN(new_n361));
  INV_X1    g175(.A(G478), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n355), .B1(KEYINPUT15), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G952), .ZN(new_n365));
  AOI211_X1 g179(.A(G953), .B(new_n365), .C1(G234), .C2(G237), .ZN(new_n366));
  INV_X1    g180(.A(G953), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n188), .B(new_n367), .C1(G234), .C2(G237), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT21), .B(G898), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n372));
  XNOR2_X1  g186(.A(G125), .B(G140), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n373), .A2(new_n192), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n373), .B(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n377), .B2(new_n192), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n367), .A3(G214), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n194), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT18), .B(G131), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n380), .B(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT88), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n377), .B2(KEYINPUT19), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n381), .A2(G131), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n242), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n394));
  INV_X1    g208(.A(G125), .ZN(new_n395));
  OR3_X1    g209(.A1(new_n395), .A2(KEYINPUT16), .A3(G140), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(G146), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n387), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n201), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT89), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(KEYINPUT89), .A3(new_n402), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n396), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n192), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(new_n397), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n381), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(new_n409), .C1(KEYINPUT17), .C2(new_n393), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n387), .A3(new_n401), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n372), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n411), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n372), .B(new_n413), .C1(new_n415), .C2(new_n403), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n410), .A2(new_n387), .A3(new_n401), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n401), .B1(new_n410), .B2(new_n387), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n188), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n421), .A2(G475), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n364), .A2(new_n371), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G221), .B1(new_n345), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n301), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n264), .A2(G125), .ZN(new_n429));
  INV_X1    g243(.A(new_n255), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(G125), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n367), .A2(G224), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n433), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G119), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G116), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT2), .B(G113), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(KEYINPUT69), .A2(G116), .ZN(new_n443));
  NOR2_X1   g257(.A1(KEYINPUT69), .A2(G116), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT70), .B1(new_n445), .B2(G119), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n447));
  NOR4_X1   g261(.A1(new_n443), .A2(new_n444), .A3(new_n447), .A4(new_n439), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n440), .B(new_n442), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(KEYINPUT71), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n451));
  INV_X1    g265(.A(new_n440), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n304), .A2(G119), .A3(new_n305), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n447), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n304), .A2(KEYINPUT70), .A3(G119), .A4(new_n305), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n451), .B1(new_n456), .B2(new_n442), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n441), .A2(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(KEYINPUT68), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI22_X1  g274(.A1(new_n450), .A2(new_n457), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n270), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(KEYINPUT80), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n454), .A2(new_n455), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n465), .A2(new_n440), .B1(new_n458), .B2(new_n459), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n449), .A2(KEYINPUT71), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n451), .A3(new_n442), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n464), .B1(new_n469), .B2(new_n270), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n468), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g286(.A(G113), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n452), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n226), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n463), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT81), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n463), .A2(new_n470), .A3(new_n480), .A4(new_n477), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT82), .Z(new_n483));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT6), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(new_n481), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n482), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n478), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT6), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n483), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n478), .B2(KEYINPUT81), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n486), .B1(new_n493), .B2(new_n481), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n438), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n436), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT85), .B(KEYINPUT7), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n432), .B1(new_n434), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n482), .B(KEYINPUT8), .Z(new_n503));
  OR2_X1    g317(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n475), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n471), .A3(new_n226), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n471), .A2(new_n476), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n212), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n436), .A2(new_n497), .A3(new_n498), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n502), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n489), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n495), .A2(new_n496), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n496), .B1(new_n495), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n428), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n427), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n244), .A2(new_n264), .ZN(new_n520));
  AOI21_X1  g334(.A(G134), .B1(new_n236), .B2(new_n237), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n234), .A2(G137), .ZN(new_n522));
  OAI21_X1  g336(.A(G131), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n255), .A2(new_n243), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT72), .B(KEYINPUT30), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n520), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT72), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT30), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n520), .B2(new_n524), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n461), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n379), .A2(new_n367), .A3(G210), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT27), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND3_X1  g348(.A1(new_n469), .A2(new_n520), .A3(new_n524), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT31), .ZN(new_n537));
  INV_X1    g351(.A(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n520), .A2(new_n524), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n461), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT28), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n461), .A2(new_n539), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n535), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n538), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n530), .A2(new_n546), .A3(new_n534), .A4(new_n535), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n537), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G472), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n188), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT74), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  OR3_X1    g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n541), .A2(new_n544), .A3(new_n538), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n556), .B2(KEYINPUT29), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n556), .A2(KEYINPUT29), .ZN(new_n558));
  INV_X1    g372(.A(new_n528), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n539), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n520), .A2(new_n524), .A3(new_n525), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n469), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n538), .B1(new_n562), .B2(new_n540), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT73), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n538), .C1(new_n562), .C2(new_n540), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n557), .B1(new_n558), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G472), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n407), .A2(new_n397), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n439), .B2(G128), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n573), .B(new_n574), .C1(G119), .C2(new_n198), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G110), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n439), .A2(KEYINPUT75), .A3(G128), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT75), .B1(new_n439), .B2(G128), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(G119), .C2(new_n198), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT24), .B(G110), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n571), .B(new_n576), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(G110), .B2(new_n575), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(new_n397), .A3(new_n375), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT22), .B(G137), .Z(new_n586));
  NAND3_X1  g400(.A1(new_n367), .A2(G221), .A3(G234), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n585), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n188), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n346), .B1(G234), .B2(new_n188), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n590), .B2(new_n188), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n593), .A2(G902), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n590), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n570), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n519), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT96), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT95), .B(G101), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  NAND2_X1  g418(.A1(new_n517), .A2(KEYINPUT97), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n428), .C1(new_n515), .C2(new_n516), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n370), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n598), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n548), .A2(new_n188), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n550), .ZN(new_n612));
  NOR4_X1   g426(.A1(new_n301), .A2(new_n609), .A3(new_n426), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n356), .A2(new_n362), .A3(new_n358), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n356), .A2(KEYINPUT100), .A3(new_n362), .A4(new_n358), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n353), .A2(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n352), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT33), .B1(new_n352), .B2(new_n620), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n344), .A2(KEYINPUT98), .A3(new_n353), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n625), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n621), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n348), .A2(new_n627), .A3(new_n354), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n362), .A2(G902), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n423), .B1(new_n618), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n608), .A2(new_n613), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT101), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT34), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G104), .ZN(G6));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n416), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n414), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n421), .A2(KEYINPUT103), .A3(G475), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT103), .B1(new_n421), .B2(G475), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n412), .A2(new_n413), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n364), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n608), .A2(new_n613), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n585), .B(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n596), .B1(new_n597), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n612), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n519), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NOR2_X1   g470(.A1(new_n645), .A2(new_n639), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n368), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n366), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n657), .A2(new_n363), .A3(new_n361), .A4(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n301), .A2(new_n426), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n652), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n570), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n495), .A2(new_n514), .ZN(new_n669));
  INV_X1    g483(.A(new_n496), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n495), .A2(new_n496), .A3(new_n514), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n606), .B1(new_n673), .B2(new_n428), .ZN(new_n674));
  INV_X1    g488(.A(new_n607), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n668), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT105), .B(G128), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G30));
  XNOR2_X1  g493(.A(new_n661), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n665), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT40), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n673), .B(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n536), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n534), .B1(new_n543), .B2(new_n535), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n188), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G472), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n364), .A2(new_n423), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n428), .A3(new_n652), .A4(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n682), .A2(new_n684), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT107), .B(G143), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G45));
  NAND2_X1  g508(.A1(new_n618), .A2(new_n631), .ZN(new_n695));
  INV_X1    g509(.A(new_n423), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n661), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT108), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n632), .A2(new_n699), .A3(new_n661), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n665), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n676), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n192), .ZN(G48));
  INV_X1    g517(.A(new_n278), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n294), .A2(new_n245), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n291), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n254), .B2(new_n283), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n188), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n425), .A3(new_n288), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n599), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n608), .A2(new_n632), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT109), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND3_X1  g529(.A1(new_n608), .A2(new_n646), .A3(new_n711), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND2_X1  g531(.A1(new_n570), .A2(new_n667), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n424), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n605), .A2(new_n607), .ZN(new_n721));
  INV_X1    g535(.A(new_n710), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI211_X1 g537(.A(KEYINPUT110), .B(new_n710), .C1(new_n605), .C2(new_n607), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT111), .B(new_n719), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AND2_X1   g544(.A1(new_n721), .A2(new_n690), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n550), .A2(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n550), .A2(KEYINPUT112), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n611), .A3(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(new_n609), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n370), .A3(new_n710), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  AOI21_X1  g552(.A(new_n699), .B1(new_n632), .B2(new_n661), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n616), .A2(new_n617), .B1(new_n629), .B2(new_n630), .ZN(new_n740));
  INV_X1    g554(.A(new_n661), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n423), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n734), .A2(new_n652), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n723), .B2(new_n724), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NAND4_X1  g561(.A1(new_n671), .A2(new_n428), .A3(new_n672), .A4(new_n425), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n297), .A2(new_n749), .A3(new_n288), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n749), .B1(new_n297), .B2(new_n288), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n569), .A2(new_n554), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n550), .A2(new_n552), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n609), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n698), .A3(new_n700), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n743), .A2(new_n760), .A3(new_n600), .A4(new_n753), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n759), .B1(new_n758), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND3_X1  g579(.A1(new_n664), .A2(new_n600), .A3(new_n753), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  XOR2_X1   g581(.A(new_n296), .B(KEYINPUT45), .Z(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n768), .B2(G902), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n289), .B1(new_n769), .B2(KEYINPUT46), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n426), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(new_n680), .ZN(new_n773));
  INV_X1    g587(.A(new_n428), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n673), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n740), .A2(new_n696), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT43), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n612), .A3(new_n667), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n773), .B(new_n781), .C1(new_n780), .C2(new_n779), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  XNOR2_X1  g597(.A(new_n772), .B(KEYINPUT47), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n776), .A2(new_n570), .A3(new_n598), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n743), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  NAND2_X1  g601(.A1(new_n709), .A2(new_n288), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n598), .A2(new_n366), .ZN(new_n789));
  OR4_X1    g603(.A1(new_n689), .A2(new_n748), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n632), .ZN(new_n791));
  OAI211_X1 g605(.A(G952), .B(new_n367), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n722), .B1(new_n674), .B2(new_n675), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n721), .A2(new_n720), .A3(new_n722), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n778), .A2(new_n366), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n735), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n792), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n797), .A2(new_n788), .A3(new_n748), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n756), .ZN(new_n802));
  NOR2_X1   g616(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n802), .B(new_n803), .Z(new_n804));
  NAND3_X1  g618(.A1(new_n684), .A2(new_n774), .A3(new_n722), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT116), .Z(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n798), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT50), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n790), .A2(new_n696), .A3(new_n695), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n801), .B2(new_n744), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n788), .A2(new_n425), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n775), .B(new_n798), .C1(new_n784), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  OAI221_X1 g630(.A(new_n799), .B1(new_n800), .B2(new_n804), .C1(new_n808), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n808), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n814), .A2(new_n810), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n737), .A2(new_n712), .A3(new_n716), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n727), .B2(new_n728), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n743), .A2(new_n744), .A3(new_n753), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n364), .A2(new_n667), .A3(new_n657), .A4(new_n661), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n775), .A3(new_n570), .A4(new_n665), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n826), .A3(new_n766), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n762), .A2(new_n763), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n427), .B(new_n518), .C1(new_n600), .C2(new_n653), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n791), .B1(new_n364), .B2(new_n696), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n613), .A2(new_n830), .A3(new_n518), .A4(new_n371), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n823), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n676), .B1(new_n666), .B2(new_n701), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n796), .B2(new_n745), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n752), .A2(new_n426), .A3(new_n667), .A4(new_n741), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n731), .A2(new_n689), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n718), .B1(new_n605), .B2(new_n607), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n665), .C1(new_n743), .C2(new_n664), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n746), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT53), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n823), .A2(new_n833), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n828), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n837), .B1(new_n836), .B2(new_n839), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n837), .A2(new_n746), .A3(new_n839), .A4(new_n842), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT115), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n840), .A2(new_n844), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(KEYINPUT54), .B(new_n846), .C1(new_n850), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n758), .A2(new_n761), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT53), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n827), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n822), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n729), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n853), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n849), .B1(new_n834), .B2(new_n845), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n821), .A2(new_n857), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(G952), .B2(G953), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n788), .B(KEYINPUT49), .ZN(new_n869));
  INV_X1    g683(.A(new_n777), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n598), .A2(new_n428), .A3(new_n425), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n869), .A2(new_n689), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n684), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n367), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n188), .B1(new_n863), .B2(new_n864), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT56), .B1(new_n877), .B2(G210), .ZN(new_n878));
  OR3_X1    g692(.A1(new_n491), .A2(new_n438), .A3(new_n494), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n495), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT55), .Z(new_n881));
  OAI21_X1  g695(.A(new_n876), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n878), .B2(new_n881), .ZN(G51));
  XNOR2_X1  g697(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g698(.A1(G469), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n866), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n707), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n877), .A2(G469), .A3(new_n768), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n875), .B1(new_n893), .B2(new_n894), .ZN(G54));
  AND3_X1   g709(.A1(new_n877), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n876), .B1(new_n896), .B2(new_n412), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n412), .B2(new_n896), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n866), .B2(new_n857), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n876), .B1(new_n901), .B2(new_n629), .ZN(new_n902));
  INV_X1    g716(.A(new_n900), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n629), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n890), .B2(new_n891), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT121), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n907), .B(new_n904), .C1(new_n890), .C2(new_n891), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n902), .B1(new_n906), .B2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT60), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n865), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n589), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n865), .A2(new_n651), .A3(new_n911), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(KEYINPUT61), .A3(new_n876), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n865), .A2(new_n917), .A3(new_n651), .A4(new_n911), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(new_n913), .A3(new_n876), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(G66));
  NAND2_X1  g738(.A1(G224), .A2(G953), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n847), .A2(G953), .B1(new_n369), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n367), .A2(G898), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n491), .A2(new_n494), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  NOR2_X1   g743(.A1(new_n526), .A2(new_n529), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n389), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n280), .ZN(new_n933));
  OAI21_X1  g747(.A(G900), .B1(new_n931), .B2(G227), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n773), .A2(new_n731), .A3(new_n756), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n786), .A2(new_n936), .A3(new_n766), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n782), .A2(KEYINPUT125), .A3(new_n836), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT125), .B1(new_n782), .B2(new_n836), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n937), .B(new_n764), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n746), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n941), .A2(new_n692), .A3(new_n835), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT62), .ZN(new_n943));
  INV_X1    g757(.A(new_n681), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n600), .A3(new_n775), .A4(new_n830), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n943), .A2(new_n782), .A3(new_n786), .A4(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  MUX2_X1   g762(.A(new_n940), .B(new_n948), .S(new_n932), .Z(new_n949));
  OAI21_X1  g763(.A(new_n935), .B1(new_n949), .B2(G953), .ZN(G72));
  XNOR2_X1  g764(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n549), .A2(new_n188), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT127), .Z(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n940), .B2(new_n847), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n562), .A2(new_n534), .A3(new_n540), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n875), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n846), .B1(new_n850), .B2(new_n856), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n953), .B1(new_n567), .B2(new_n685), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n948), .A2(new_n848), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n954), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n538), .B1(new_n530), .B2(new_n535), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G57));
endmodule


