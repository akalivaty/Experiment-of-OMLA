

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U557 ( .A1(n767), .A2(n769), .ZN(n724) );
  INV_X1 U558 ( .A(n724), .ZN(n710) );
  NAND2_X1 U559 ( .A1(G8), .A2(n724), .ZN(n763) );
  NAND2_X1 U560 ( .A1(n706), .A2(n705), .ZN(n708) );
  NOR2_X1 U561 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U562 ( .A(n717), .B(n716), .Z(n522) );
  NAND2_X1 U563 ( .A1(n763), .A2(n757), .ZN(n523) );
  XOR2_X1 U564 ( .A(n771), .B(KEYINPUT89), .Z(n524) );
  XNOR2_X1 U565 ( .A(KEYINPUT30), .B(KEYINPUT95), .ZN(n716) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n707) );
  NAND2_X1 U567 ( .A1(n723), .A2(n722), .ZN(n734) );
  AND2_X1 U568 ( .A1(n734), .A2(n733), .ZN(n737) );
  XNOR2_X1 U569 ( .A(n738), .B(KEYINPUT96), .ZN(n739) );
  NOR2_X1 U570 ( .A1(G164), .A2(G1384), .ZN(n769) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n530), .Z(n647) );
  AND2_X1 U572 ( .A1(n550), .A2(G2104), .ZN(n889) );
  XNOR2_X1 U573 ( .A(n583), .B(KEYINPUT15), .ZN(n1022) );
  NOR2_X1 U574 ( .A1(G651), .A2(n622), .ZN(n646) );
  AND2_X1 U575 ( .A1(G138), .A2(n890), .ZN(n556) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n644) );
  NAND2_X1 U577 ( .A1(n644), .A2(G89), .ZN(n525) );
  XNOR2_X1 U578 ( .A(n525), .B(KEYINPUT4), .ZN(n527) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  INV_X1 U580 ( .A(G651), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n622), .A2(n529), .ZN(n651) );
  NAND2_X1 U582 ( .A1(G76), .A2(n651), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n528), .B(KEYINPUT5), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G51), .A2(n646), .ZN(n532) );
  NOR2_X1 U586 ( .A1(G543), .A2(n529), .ZN(n530) );
  NAND2_X1 U587 ( .A1(G63), .A2(n647), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U589 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U591 ( .A(n536), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(n537) );
  XNOR2_X1 U593 ( .A(KEYINPUT74), .B(n537), .ZN(G286) );
  NAND2_X1 U594 ( .A1(G64), .A2(n647), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n538), .B(KEYINPUT66), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G52), .A2(n646), .ZN(n539) );
  XOR2_X1 U597 ( .A(KEYINPUT67), .B(n539), .Z(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n651), .A2(G77), .ZN(n542) );
  XNOR2_X1 U600 ( .A(KEYINPUT69), .B(n542), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n644), .A2(G90), .ZN(n543) );
  XOR2_X1 U602 ( .A(KEYINPUT68), .B(n543), .Z(n544) );
  NOR2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT9), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U607 ( .A1(G2104), .A2(G2105), .ZN(n549) );
  XOR2_X2 U608 ( .A(KEYINPUT17), .B(n549), .Z(n890) );
  INV_X1 U609 ( .A(G2105), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G102), .A2(n889), .ZN(n554) );
  AND2_X1 U611 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U612 ( .A1(G114), .A2(n893), .ZN(n552) );
  INV_X1 U613 ( .A(G2104), .ZN(n558) );
  AND2_X1 U614 ( .A1(n558), .A2(G2105), .ZN(n894) );
  NAND2_X1 U615 ( .A1(G126), .A2(n894), .ZN(n551) );
  AND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U619 ( .A1(G101), .A2(n889), .ZN(n557) );
  XNOR2_X1 U620 ( .A(KEYINPUT23), .B(n557), .ZN(n563) );
  AND2_X1 U621 ( .A1(n558), .A2(G125), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G2105), .A2(n559), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G113), .A2(n893), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n683) );
  NAND2_X1 U626 ( .A1(n890), .A2(G137), .ZN(n685) );
  AND2_X1 U627 ( .A1(n683), .A2(n685), .ZN(G160) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT10), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT72), .B(n565), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n832) );
  NAND2_X1 U635 ( .A1(n832), .A2(G567), .ZN(n566) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  XNOR2_X1 U637 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n644), .A2(G81), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U640 ( .A1(G68), .A2(n651), .ZN(n568) );
  NAND2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U642 ( .A(n571), .B(n570), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n647), .A2(G56), .ZN(n572) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n646), .A2(G43), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n1003) );
  INV_X1 U648 ( .A(G860), .ZN(n839) );
  OR2_X1 U649 ( .A1(n1003), .A2(n839), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G54), .A2(n646), .ZN(n578) );
  NAND2_X1 U653 ( .A1(G66), .A2(n647), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G92), .A2(n644), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G79), .A2(n651), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U659 ( .A(G868), .ZN(n665) );
  NAND2_X1 U660 ( .A1(n1022), .A2(n665), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U662 ( .A1(n644), .A2(G91), .ZN(n586) );
  XNOR2_X1 U663 ( .A(n586), .B(KEYINPUT70), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G65), .A2(n647), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G78), .A2(n651), .ZN(n590) );
  NAND2_X1 U667 ( .A1(G53), .A2(n646), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n1025) );
  XNOR2_X1 U670 ( .A(n1025), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G299), .A2(n665), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n839), .A2(G559), .ZN(n595) );
  INV_X1 U675 ( .A(n1022), .ZN(n641) );
  NAND2_X1 U676 ( .A1(n595), .A2(n641), .ZN(n596) );
  XNOR2_X1 U677 ( .A(n596), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(n1022), .A2(n665), .ZN(n597) );
  XNOR2_X1 U679 ( .A(n597), .B(KEYINPUT75), .ZN(n598) );
  NOR2_X1 U680 ( .A1(G559), .A2(n598), .ZN(n600) );
  NOR2_X1 U681 ( .A1(G868), .A2(n1003), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G123), .A2(n894), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n601), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G111), .A2(n893), .ZN(n602) );
  XNOR2_X1 U686 ( .A(n602), .B(KEYINPUT76), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G99), .A2(n889), .ZN(n606) );
  NAND2_X1 U689 ( .A1(G135), .A2(n890), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n981) );
  XNOR2_X1 U692 ( .A(G2096), .B(n981), .ZN(n610) );
  INV_X1 U693 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G88), .A2(n644), .ZN(n612) );
  NAND2_X1 U696 ( .A1(G75), .A2(n651), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n647), .A2(G62), .ZN(n613) );
  XOR2_X1 U699 ( .A(KEYINPUT84), .B(n613), .Z(n614) );
  NOR2_X1 U700 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n646), .A2(G50), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(G303) );
  NAND2_X1 U703 ( .A1(G49), .A2(n646), .ZN(n619) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n618) );
  NAND2_X1 U705 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U706 ( .A1(n647), .A2(n620), .ZN(n621) );
  XNOR2_X1 U707 ( .A(n621), .B(KEYINPUT82), .ZN(n624) );
  NAND2_X1 U708 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U710 ( .A1(n647), .A2(G60), .ZN(n625) );
  XNOR2_X1 U711 ( .A(n625), .B(KEYINPUT64), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G85), .A2(n644), .ZN(n627) );
  NAND2_X1 U713 ( .A1(G72), .A2(n651), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G47), .A2(n646), .ZN(n628) );
  XNOR2_X1 U716 ( .A(KEYINPUT65), .B(n628), .ZN(n629) );
  NOR2_X1 U717 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G73), .A2(n651), .ZN(n633) );
  XNOR2_X1 U720 ( .A(n633), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G86), .A2(n644), .ZN(n635) );
  NAND2_X1 U722 ( .A1(G48), .A2(n646), .ZN(n634) );
  NAND2_X1 U723 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U724 ( .A1(G61), .A2(n647), .ZN(n636) );
  XNOR2_X1 U725 ( .A(KEYINPUT83), .B(n636), .ZN(n637) );
  NOR2_X1 U726 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U727 ( .A1(n640), .A2(n639), .ZN(G305) );
  XNOR2_X1 U728 ( .A(n1003), .B(KEYINPUT77), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n641), .A2(G559), .ZN(n642) );
  XNOR2_X1 U730 ( .A(n643), .B(n642), .ZN(n838) );
  XOR2_X1 U731 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n659) );
  NAND2_X1 U732 ( .A1(G93), .A2(n644), .ZN(n645) );
  XNOR2_X1 U733 ( .A(n645), .B(KEYINPUT78), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G55), .A2(n646), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G67), .A2(n647), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U737 ( .A(KEYINPUT80), .B(n650), .ZN(n654) );
  NAND2_X1 U738 ( .A1(G80), .A2(n651), .ZN(n652) );
  XNOR2_X1 U739 ( .A(KEYINPUT79), .B(n652), .ZN(n653) );
  NOR2_X1 U740 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U741 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U742 ( .A(KEYINPUT81), .B(n657), .Z(n840) );
  XNOR2_X1 U743 ( .A(G303), .B(n840), .ZN(n658) );
  XNOR2_X1 U744 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n661), .B(G299), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n662), .B(G290), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(G305), .ZN(n905) );
  XNOR2_X1 U749 ( .A(n838), .B(n905), .ZN(n664) );
  NAND2_X1 U750 ( .A1(n664), .A2(G868), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n665), .A2(n840), .ZN(n666) );
  NAND2_X1 U752 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U755 ( .A1(n669), .A2(G2090), .ZN(n670) );
  XNOR2_X1 U756 ( .A(n670), .B(KEYINPUT86), .ZN(n671) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U758 ( .A1(G2072), .A2(n672), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U762 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U763 ( .A1(G96), .A2(n675), .ZN(n836) );
  NAND2_X1 U764 ( .A1(n836), .A2(G2106), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G120), .A2(G108), .ZN(n676) );
  NOR2_X1 U766 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U767 ( .A1(G69), .A2(n677), .ZN(n837) );
  NAND2_X1 U768 ( .A1(n837), .A2(G567), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n842) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U771 ( .A1(n842), .A2(n680), .ZN(n681) );
  XOR2_X1 U772 ( .A(KEYINPUT87), .B(n681), .Z(n835) );
  NAND2_X1 U773 ( .A1(G36), .A2(n835), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n682), .B(KEYINPUT88), .ZN(G176) );
  AND2_X1 U775 ( .A1(n683), .A2(G40), .ZN(n684) );
  AND2_X1 U776 ( .A1(n685), .A2(n684), .ZN(n767) );
  NAND2_X1 U777 ( .A1(n710), .A2(G2072), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n687), .B(KEYINPUT27), .ZN(n689) );
  AND2_X1 U779 ( .A1(G1956), .A2(n724), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U781 ( .A1(n1025), .A2(n691), .ZN(n690) );
  XOR2_X1 U782 ( .A(n690), .B(KEYINPUT28), .Z(n706) );
  NAND2_X1 U783 ( .A1(n1025), .A2(n691), .ZN(n704) );
  NAND2_X1 U784 ( .A1(G1348), .A2(n724), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n710), .A2(G2067), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n700) );
  NOR2_X1 U787 ( .A1(n1022), .A2(n700), .ZN(n699) );
  INV_X1 U788 ( .A(G1996), .ZN(n917) );
  NOR2_X1 U789 ( .A1(n724), .A2(n917), .ZN(n694) );
  XOR2_X1 U790 ( .A(n694), .B(KEYINPUT26), .Z(n696) );
  NAND2_X1 U791 ( .A1(n724), .A2(G1341), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U793 ( .A1(n1003), .A2(n697), .ZN(n698) );
  OR2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n1022), .A2(n700), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n708), .B(n707), .ZN(n714) );
  INV_X1 U799 ( .A(G1961), .ZN(n937) );
  NAND2_X1 U800 ( .A1(n724), .A2(n937), .ZN(n712) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n709) );
  XNOR2_X1 U802 ( .A(n709), .B(KEYINPUT94), .ZN(n918) );
  NAND2_X1 U803 ( .A1(n710), .A2(n918), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U805 ( .A1(G171), .A2(n718), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n723) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n763), .ZN(n732) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n724), .ZN(n735) );
  NOR2_X1 U809 ( .A1(n732), .A2(n735), .ZN(n715) );
  NAND2_X1 U810 ( .A1(G8), .A2(n715), .ZN(n717) );
  NOR2_X1 U811 ( .A1(G168), .A2(n522), .ZN(n720) );
  NOR2_X1 U812 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U814 ( .A(n721), .B(KEYINPUT31), .Z(n722) );
  NAND2_X1 U815 ( .A1(n734), .A2(G286), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n763), .ZN(n726) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n727), .A2(G303), .ZN(n728) );
  NAND2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U822 ( .A(n731), .B(KEYINPUT32), .ZN(n740) );
  INV_X1 U823 ( .A(n732), .ZN(n733) );
  NAND2_X1 U824 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n756) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n1027) );
  NOR2_X1 U829 ( .A1(n1005), .A2(n1027), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n756), .A2(n741), .ZN(n742) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n1020) );
  NAND2_X1 U832 ( .A1(n742), .A2(n1020), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n1005), .A2(KEYINPUT33), .ZN(n743) );
  NOR2_X1 U834 ( .A1(n743), .A2(n763), .ZN(n745) );
  XOR2_X1 U835 ( .A(G1981), .B(G305), .Z(n1014) );
  INV_X1 U836 ( .A(n1014), .ZN(n744) );
  NOR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n749) );
  INV_X1 U838 ( .A(n749), .ZN(n746) );
  OR2_X1 U839 ( .A1(n763), .A2(n746), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n751) );
  AND2_X1 U841 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U843 ( .A(n752), .B(KEYINPUT97), .ZN(n753) );
  INV_X1 U844 ( .A(n753), .ZN(n758) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U846 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n523), .ZN(n759) );
  XNOR2_X1 U849 ( .A(n759), .B(KEYINPUT98), .ZN(n765) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XNOR2_X1 U851 ( .A(n760), .B(KEYINPUT93), .ZN(n761) );
  XNOR2_X1 U852 ( .A(n761), .B(KEYINPUT24), .ZN(n762) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U854 ( .A(n766), .B(KEYINPUT99), .ZN(n772) );
  NOR2_X1 U855 ( .A1(G1986), .A2(G290), .ZN(n806) );
  INV_X1 U856 ( .A(n806), .ZN(n1010) );
  NAND2_X1 U857 ( .A1(G1986), .A2(G290), .ZN(n1021) );
  NAND2_X1 U858 ( .A1(n1010), .A2(n1021), .ZN(n770) );
  INV_X1 U859 ( .A(n767), .ZN(n768) );
  NOR2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n813) );
  NAND2_X1 U861 ( .A1(n770), .A2(n813), .ZN(n771) );
  AND2_X1 U862 ( .A1(n772), .A2(n524), .ZN(n802) );
  NAND2_X1 U863 ( .A1(G107), .A2(n893), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G119), .A2(n894), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G95), .A2(n889), .ZN(n776) );
  NAND2_X1 U867 ( .A1(G131), .A2(n890), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n871) );
  NAND2_X1 U870 ( .A1(G1991), .A2(n871), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT91), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G129), .A2(n894), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G141), .A2(n890), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G105), .A2(n889), .ZN(n782) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n782), .Z(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n893), .A2(G117), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n882) );
  AND2_X1 U880 ( .A1(G1996), .A2(n882), .ZN(n787) );
  NOR2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n983) );
  XOR2_X1 U882 ( .A(KEYINPUT92), .B(n813), .Z(n789) );
  NOR2_X1 U883 ( .A1(n983), .A2(n789), .ZN(n809) );
  INV_X1 U884 ( .A(n809), .ZN(n800) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n803) );
  NAND2_X1 U886 ( .A1(G116), .A2(n893), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G128), .A2(n894), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U889 ( .A(KEYINPUT35), .B(n792), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G104), .A2(n889), .ZN(n794) );
  NAND2_X1 U891 ( .A1(G140), .A2(n890), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n796) );
  XOR2_X1 U893 ( .A(KEYINPUT90), .B(KEYINPUT34), .Z(n795) );
  XNOR2_X1 U894 ( .A(n796), .B(n795), .ZN(n797) );
  NAND2_X1 U895 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U896 ( .A(KEYINPUT36), .B(n799), .Z(n902) );
  NOR2_X1 U897 ( .A1(n803), .A2(n902), .ZN(n986) );
  NAND2_X1 U898 ( .A1(n986), .A2(n813), .ZN(n804) );
  AND2_X1 U899 ( .A1(n800), .A2(n804), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n820) );
  AND2_X1 U901 ( .A1(n803), .A2(n902), .ZN(n993) );
  NAND2_X1 U902 ( .A1(n993), .A2(n813), .ZN(n818) );
  INV_X1 U903 ( .A(n804), .ZN(n816) );
  XNOR2_X1 U904 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n805) );
  XNOR2_X1 U905 ( .A(n805), .B(KEYINPUT39), .ZN(n812) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n882), .ZN(n978) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n871), .ZN(n982) );
  NOR2_X1 U908 ( .A1(n806), .A2(n982), .ZN(n807) );
  XNOR2_X1 U909 ( .A(n807), .B(KEYINPUT100), .ZN(n808) );
  NOR2_X1 U910 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U911 ( .A1(n978), .A2(n810), .ZN(n811) );
  XOR2_X1 U912 ( .A(n812), .B(n811), .Z(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  AND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U918 ( .A(G2454), .B(G2435), .Z(n823) );
  XNOR2_X1 U919 ( .A(G2438), .B(G2427), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n830) );
  XOR2_X1 U921 ( .A(KEYINPUT103), .B(G2446), .Z(n825) );
  XNOR2_X1 U922 ( .A(G2443), .B(G2430), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U924 ( .A(n826), .B(G2451), .Z(n828) );
  XNOR2_X1 U925 ( .A(G1341), .B(G1348), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n831), .A2(G14), .ZN(n911) );
  XOR2_X1 U929 ( .A(KEYINPUT104), .B(n911), .Z(G401) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U932 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U935 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  NOR2_X1 U939 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  NAND2_X1 U941 ( .A1(n839), .A2(n838), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(G145) );
  INV_X1 U943 ( .A(n842), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n845), .B(G2096), .Z(n847) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2678), .Z(n849) );
  XNOR2_X1 U951 ( .A(KEYINPUT105), .B(G2100), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(G227) );
  XOR2_X1 U954 ( .A(G1976), .B(G1966), .Z(n853) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1981), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U958 ( .A(G1961), .B(G1956), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT41), .B(G1971), .Z(n858) );
  XNOR2_X1 U961 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G100), .A2(n889), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G112), .A2(n893), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G124), .A2(n894), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n863), .B(KEYINPUT44), .ZN(n864) );
  XNOR2_X1 U969 ( .A(n864), .B(KEYINPUT106), .ZN(n866) );
  NAND2_X1 U970 ( .A1(G136), .A2(n890), .ZN(n865) );
  NAND2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U972 ( .A(KEYINPUT107), .B(n867), .Z(n868) );
  NOR2_X1 U973 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U974 ( .A(G160), .B(n981), .Z(n870) );
  XNOR2_X1 U975 ( .A(n871), .B(n870), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G106), .A2(n889), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G142), .A2(n890), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n874), .B(KEYINPUT45), .ZN(n876) );
  NAND2_X1 U980 ( .A1(G118), .A2(n893), .ZN(n875) );
  NAND2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n894), .A2(G130), .ZN(n877) );
  XOR2_X1 U983 ( .A(KEYINPUT108), .B(n877), .Z(n878) );
  NOR2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U985 ( .A(n881), .B(n880), .Z(n884) );
  XOR2_X1 U986 ( .A(n882), .B(G162), .Z(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n886) );
  XNOR2_X1 U989 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U991 ( .A(n888), .B(n887), .Z(n901) );
  NAND2_X1 U992 ( .A1(G103), .A2(n889), .ZN(n892) );
  NAND2_X1 U993 ( .A1(G139), .A2(n890), .ZN(n891) );
  NAND2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U995 ( .A1(G115), .A2(n893), .ZN(n896) );
  NAND2_X1 U996 ( .A1(G127), .A2(n894), .ZN(n895) );
  NAND2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n973) );
  XNOR2_X1 U1000 ( .A(G164), .B(n973), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n905), .B(n1003), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(n1022), .ZN(n908) );
  XOR2_X1 U1006 ( .A(G286), .B(G171), .Z(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n909), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT111), .B(n910), .Z(G397) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n911), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G303), .ZN(G166) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1019 ( .A(G32), .B(n917), .ZN(n922) );
  XOR2_X1 U1020 ( .A(n918), .B(G27), .Z(n920) );
  XNOR2_X1 U1021 ( .A(G26), .B(G2067), .ZN(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(KEYINPUT116), .B(n925), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n926), .A2(G28), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G25), .B(G1991), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1030 ( .A(KEYINPUT53), .B(n929), .Z(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(G34), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(G2084), .B(n931), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n966) );
  NAND2_X1 U1037 ( .A1(KEYINPUT55), .A2(n966), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(G11), .A2(n936), .ZN(n972) );
  XNOR2_X1 U1039 ( .A(n937), .B(G5), .ZN(n961) );
  XOR2_X1 U1040 ( .A(G1966), .B(G21), .Z(n949) );
  XOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .Z(n938) );
  XNOR2_X1 U1042 ( .A(G4), .B(n938), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G1341), .B(G19), .ZN(n939) );
  XNOR2_X1 U1044 ( .A(n939), .B(KEYINPUT122), .ZN(n943) );
  XOR2_X1 U1045 ( .A(G1981), .B(G6), .Z(n941) );
  XOR2_X1 U1046 ( .A(G1956), .B(G20), .Z(n940) );
  NAND2_X1 U1047 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1048 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1049 ( .A(n944), .B(KEYINPUT123), .ZN(n945) );
  NOR2_X1 U1050 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1051 ( .A(n947), .B(KEYINPUT60), .ZN(n948) );
  NAND2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G1986), .B(G24), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n950) );
  XNOR2_X1 U1055 ( .A(n950), .B(KEYINPUT124), .ZN(n952) );
  XNOR2_X1 U1056 ( .A(G23), .B(G1976), .ZN(n951) );
  NOR2_X1 U1057 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1058 ( .A(KEYINPUT125), .B(n953), .ZN(n954) );
  NOR2_X1 U1059 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1060 ( .A(KEYINPUT58), .B(n956), .Z(n957) );
  XNOR2_X1 U1061 ( .A(KEYINPUT126), .B(n957), .ZN(n958) );
  NOR2_X1 U1062 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1064 ( .A(n962), .B(KEYINPUT127), .ZN(n963) );
  XNOR2_X1 U1065 ( .A(n963), .B(KEYINPUT61), .ZN(n965) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT121), .ZN(n964) );
  NAND2_X1 U1067 ( .A1(n965), .A2(n964), .ZN(n970) );
  INV_X1 U1068 ( .A(n966), .ZN(n968) );
  NOR2_X1 U1069 ( .A1(G29), .A2(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1070 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1071 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n1002) );
  XOR2_X1 U1073 ( .A(G2072), .B(n973), .Z(n975) );
  XOR2_X1 U1074 ( .A(G164), .B(G2078), .Z(n974) );
  NOR2_X1 U1075 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1076 ( .A(KEYINPUT50), .B(n976), .Z(n996) );
  XOR2_X1 U1077 ( .A(G2090), .B(G162), .Z(n977) );
  NOR2_X1 U1078 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1079 ( .A(KEYINPUT114), .B(n979), .Z(n980) );
  XNOR2_X1 U1080 ( .A(KEYINPUT51), .B(n980), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n982), .A2(n981), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G160), .B(G2084), .ZN(n984) );
  NAND2_X1 U1083 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(KEYINPUT113), .B(n989), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(KEYINPUT115), .B(n994), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT52), .B(n997), .ZN(n999) );
  INV_X1 U1092 ( .A(KEYINPUT55), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(G29), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1035) );
  XOR2_X1 U1096 ( .A(G16), .B(KEYINPUT56), .Z(n1033) );
  XNOR2_X1 U1097 ( .A(G171), .B(G1961), .ZN(n1019) );
  XNOR2_X1 U1098 ( .A(G1341), .B(KEYINPUT120), .ZN(n1004) );
  XNOR2_X1 U1099 ( .A(n1004), .B(n1003), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT119), .B(n1005), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  NAND2_X1 U1102 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1103 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1104 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G168), .ZN(n1012) );
  XNOR2_X1 U1106 ( .A(n1012), .B(KEYINPUT118), .ZN(n1013) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1108 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1031) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(G1348), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(n1025), .B(G1956), .Z(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(n1036), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

