//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n189), .A3(G125), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n193), .B2(new_n194), .ZN(new_n196));
  MUX2_X1   g010(.A(new_n193), .B(new_n196), .S(G146), .Z(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(new_n198), .B2(G119), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G128), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT67), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT67), .A2(G128), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .A4(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G110), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n206), .A2(KEYINPUT75), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n201), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n198), .A2(G119), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT67), .B(G128), .Z(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G119), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT24), .B(G110), .Z(new_n213));
  OAI21_X1  g027(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n197), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n190), .A2(new_n192), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT16), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G146), .A3(new_n195), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n196), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n201), .A2(new_n204), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G110), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(new_n213), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n216), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT22), .B(G137), .Z(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n228), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n216), .B1(new_n215), .B2(new_n226), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI211_X1 g049(.A(new_n216), .B(new_n232), .C1(new_n215), .C2(new_n226), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n187), .B(new_n188), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G234), .ZN(new_n238));
  OAI21_X1  g052(.A(G217), .B1(new_n238), .B2(G902), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n239), .B(KEYINPUT74), .Z(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n234), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n232), .A3(new_n227), .ZN(new_n243));
  INV_X1    g057(.A(new_n236), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n187), .B1(new_n245), .B2(new_n188), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n188), .ZN(new_n248));
  XOR2_X1   g062(.A(new_n248), .B(KEYINPUT77), .Z(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n255), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n253), .B2(new_n252), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(KEYINPUT0), .B2(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n220), .A2(G143), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT0), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT64), .B1(new_n271), .B2(new_n198), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n261), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT65), .A2(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT11), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(G137), .A3(new_n279), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(KEYINPUT11), .A3(G134), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n282), .A2(new_n285), .A3(G131), .ZN(new_n286));
  INV_X1    g100(.A(G131), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n281), .A2(KEYINPUT11), .A3(G134), .ZN(new_n288));
  AND2_X1   g102(.A1(KEYINPUT65), .A2(G134), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT65), .A2(G134), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n288), .B1(new_n291), .B2(G137), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n281), .B1(new_n289), .B2(new_n290), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT11), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n287), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n275), .B1(new_n286), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n263), .A3(G128), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n302), .A2(new_n267), .B1(new_n202), .B2(new_n203), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n263), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(new_n295), .A3(new_n287), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n293), .B1(G134), .B2(new_n281), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n297), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT70), .B1(new_n297), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n260), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n282), .B2(new_n285), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n274), .B1(new_n315), .B2(new_n305), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n314), .A2(new_n316), .A3(new_n259), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n260), .B1(new_n297), .B2(new_n308), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT28), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n317), .C2(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G210), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT27), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT30), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n297), .B2(new_n308), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n259), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n317), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n328), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT30), .B1(new_n314), .B2(new_n316), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n297), .A2(new_n332), .A3(new_n308), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n317), .B1(new_n341), .B2(new_n259), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT31), .A3(new_n328), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G472), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n330), .A2(new_n344), .A3(KEYINPUT71), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n188), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n349), .A2(new_n188), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n348), .A4(new_n347), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n313), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n335), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(KEYINPUT72), .B2(new_n335), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n359), .B2(KEYINPUT28), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT29), .A3(new_n328), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n342), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n329), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n365), .B(new_n366), .C1(new_n323), .C2(new_n329), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n360), .A2(KEYINPUT73), .A3(KEYINPUT29), .A4(new_n328), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n188), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G472), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n251), .B1(new_n355), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT9), .B(G234), .ZN(new_n372));
  OAI21_X1  g186(.A(G221), .B1(new_n372), .B2(G902), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT78), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n315), .A2(new_n305), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G107), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n377), .A2(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n267), .B1(new_n298), .B2(new_n299), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n202), .A2(new_n203), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n263), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n394), .B2(new_n301), .ZN(new_n395));
  INV_X1    g209(.A(new_n269), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n270), .A2(new_n198), .B1(new_n396), .B2(KEYINPUT1), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n301), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n389), .A2(new_n395), .B1(new_n399), .B2(new_n390), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(G101), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n274), .B1(new_n384), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n401), .A3(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT79), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n402), .A2(new_n407), .A3(new_n401), .A4(G101), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT80), .B1(new_n404), .B2(new_n409), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n376), .B(new_n400), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G140), .ZN(new_n413));
  INV_X1    g227(.A(G227), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G953), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n413), .B(new_n415), .Z(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n388), .B1(new_n301), .B2(new_n397), .ZN(new_n418));
  INV_X1    g232(.A(new_n301), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT10), .B1(new_n419), .B2(new_n393), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n418), .A2(KEYINPUT10), .B1(new_n420), .B2(new_n388), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n404), .A2(new_n409), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n404), .A2(new_n409), .A3(KEYINPUT80), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n417), .A2(KEYINPUT81), .B1(new_n376), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n417), .A2(KEYINPUT81), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n304), .A2(new_n389), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n375), .B1(new_n429), .B2(new_n418), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n432), .A2(new_n412), .ZN(new_n433));
  OAI22_X1  g247(.A1(new_n427), .A2(new_n428), .B1(new_n416), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n188), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G469), .ZN(new_n436));
  INV_X1    g250(.A(new_n416), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n424), .A2(new_n425), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n376), .B1(new_n438), .B2(new_n400), .ZN(new_n439));
  INV_X1    g253(.A(new_n412), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT83), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n417), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n412), .A2(KEYINPUT82), .A3(new_n416), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n432), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(new_n437), .C1(new_n439), .C2(new_n440), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n188), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n374), .B1(new_n436), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G113), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n377), .ZN(new_n454));
  INV_X1    g268(.A(G237), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n229), .A3(G214), .ZN(new_n456));
  NOR2_X1   g270(.A1(KEYINPUT90), .A2(G143), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n324), .B(G214), .C1(KEYINPUT90), .C2(G143), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n287), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT17), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n219), .A3(new_n221), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n458), .A2(new_n459), .A3(new_n287), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n463), .A2(new_n460), .A3(KEYINPUT17), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT18), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n287), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n193), .B(G146), .ZN(new_n469));
  INV_X1    g283(.A(new_n460), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n468), .B(new_n469), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n454), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n471), .B(new_n454), .C1(new_n464), .C2(new_n462), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT91), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n465), .A2(KEYINPUT91), .A3(new_n454), .A4(new_n471), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G475), .B1(new_n477), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n476), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n217), .B(KEYINPUT19), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI221_X1 g296(.A(new_n219), .B1(new_n463), .B2(new_n460), .C1(new_n482), .C2(G146), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n471), .ZN(new_n484));
  INV_X1    g298(.A(new_n454), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n479), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n475), .A2(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n490));
  INV_X1    g304(.A(new_n488), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n478), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G116), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(G122), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n380), .B1(new_n495), .B2(KEYINPUT14), .ZN(new_n496));
  XNOR2_X1  g310(.A(G116), .B(G122), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n498), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n202), .A2(G143), .A3(new_n203), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n268), .A2(G128), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n291), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n291), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n499), .B(new_n500), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(KEYINPUT13), .A3(new_n502), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(G134), .C1(KEYINPUT13), .C2(new_n502), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n497), .B(new_n380), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n503), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G217), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n372), .A2(new_n511), .A3(G953), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT92), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n506), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n506), .B2(new_n510), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n188), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  OAI211_X1 g334(.A(KEYINPUT93), .B(new_n188), .C1(new_n514), .C2(new_n515), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT94), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n518), .A2(new_n524), .A3(new_n520), .A4(new_n521), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n516), .A2(new_n520), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n188), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n229), .A2(G952), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n238), .B2(new_n455), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n493), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G214), .B1(G237), .B2(G902), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n419), .A2(new_n393), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n191), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT84), .B1(new_n304), .B2(G125), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n275), .A2(new_n191), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT7), .ZN(new_n543));
  INV_X1    g357(.A(G224), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G953), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n545), .A2(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(KEYINPUT89), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n403), .A2(new_n384), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n409), .A2(new_n259), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n257), .A2(new_n252), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n553));
  OR3_X1    g367(.A1(new_n494), .A2(KEYINPUT5), .A3(G119), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(G113), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n389), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G122), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n545), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n540), .A2(new_n542), .B1(KEYINPUT7), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n557), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n555), .A2(new_n552), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n384), .A2(new_n387), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n384), .A2(new_n387), .A3(new_n567), .ZN(new_n568));
  AND4_X1   g382(.A1(KEYINPUT87), .A2(new_n564), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n564), .A2(new_n566), .B1(KEYINPUT87), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n563), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT88), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT88), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(new_n563), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n562), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(KEYINPUT85), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT85), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n579), .B(new_n541), .C1(new_n538), .C2(new_n539), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n545), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n540), .A2(new_n542), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(KEYINPUT85), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n560), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n551), .A2(new_n556), .ZN(new_n586));
  INV_X1    g400(.A(new_n557), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT6), .A3(new_n558), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT6), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(new_n585), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n576), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n576), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n535), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n452), .A2(new_n534), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n371), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  INV_X1    g415(.A(new_n251), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n349), .A2(new_n188), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT71), .B1(new_n330), .B2(new_n344), .ZN(new_n604));
  OAI21_X1  g418(.A(G472), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n452), .A2(new_n602), .A3(new_n605), .A4(new_n350), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n596), .A2(new_n533), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n514), .A2(new_n515), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT33), .Z(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(G478), .A3(new_n188), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n493), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n606), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n607), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n487), .A2(new_n479), .A3(new_n488), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT20), .B1(new_n490), .B2(new_n491), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n490), .C2(new_n491), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n487), .A2(KEYINPUT96), .A3(new_n479), .A4(new_n488), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n622), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n478), .B(KEYINPUT97), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n527), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n606), .A2(new_n619), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NAND2_X1  g447(.A1(new_n215), .A2(new_n226), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n249), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n241), .B2(new_n246), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(KEYINPUT98), .B(new_n637), .C1(new_n241), .C2(new_n246), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n605), .A2(new_n642), .A3(new_n350), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n598), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT37), .B(G110), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  NAND2_X1  g460(.A1(new_n452), .A2(new_n642), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n355), .B2(new_n370), .ZN(new_n648));
  INV_X1    g462(.A(new_n528), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n532), .B1(new_n649), .B2(G900), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT99), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n628), .A2(new_n629), .A3(new_n527), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT100), .B1(new_n654), .B2(new_n597), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n653), .A2(new_n656), .A3(new_n596), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT101), .B(G128), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G30));
  INV_X1    g475(.A(new_n452), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n651), .B(KEYINPUT39), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT40), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n359), .A2(new_n329), .ZN(new_n666));
  INV_X1    g480(.A(new_n336), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n188), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n355), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n576), .A2(new_n592), .ZN(new_n671));
  INV_X1    g485(.A(new_n593), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n576), .A2(new_n592), .A3(new_n593), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n535), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n493), .A2(new_n527), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n677), .A2(new_n678), .A3(new_n642), .A4(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n665), .A2(new_n670), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  NAND2_X1  g496(.A1(new_n642), .A2(new_n597), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n355), .B2(new_n370), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n613), .A2(new_n651), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n452), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NAND2_X1  g502(.A1(new_n449), .A2(new_n188), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G469), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n451), .A3(new_n373), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n690), .A2(KEYINPUT102), .A3(new_n451), .A4(new_n373), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n371), .ZN(new_n698));
  INV_X1    g512(.A(new_n615), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NOR2_X1   g516(.A1(new_n619), .A2(new_n630), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND3_X1   g519(.A1(new_n693), .A2(new_n534), .A3(new_n695), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n684), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  OAI21_X1  g522(.A(new_n344), .B1(new_n360), .B2(new_n328), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(G472), .B2(G902), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n348), .A2(new_n188), .A3(KEYINPUT103), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n605), .A2(new_n602), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n596), .A2(new_n679), .A3(new_n533), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n693), .A2(new_n714), .A3(new_n695), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT104), .B(G122), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G24));
  AND3_X1   g532(.A1(new_n693), .A2(new_n597), .A3(new_n695), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n605), .A2(new_n642), .A3(new_n713), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n605), .A2(new_n642), .A3(KEYINPUT105), .A4(new_n713), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n685), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NAND2_X1  g542(.A1(new_n436), .A2(new_n451), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n675), .A2(new_n678), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n729), .A2(new_n730), .A3(new_n373), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n371), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n371), .A2(KEYINPUT42), .A3(new_n726), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  NAND3_X1  g551(.A1(new_n371), .A2(new_n654), .A3(new_n731), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  INV_X1    g553(.A(new_n493), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n612), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT43), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n605), .A2(new_n350), .B1(new_n640), .B2(new_n641), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n742), .B1(new_n743), .B2(KEYINPUT107), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT44), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n730), .B(KEYINPUT108), .Z(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n663), .ZN(new_n749));
  INV_X1    g563(.A(new_n373), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n434), .B(KEYINPUT45), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n751), .B2(G902), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n753));
  INV_X1    g567(.A(new_n451), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n750), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT44), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n748), .A2(new_n749), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  AND3_X1   g573(.A1(new_n685), .A2(new_n251), .A3(new_n730), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(new_n370), .A3(new_n355), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n753), .A2(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n373), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n766), .B1(new_n763), .B2(new_n765), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n761), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NOR2_X1   g584(.A1(new_n596), .A2(new_n679), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n651), .B(KEYINPUT114), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n638), .A2(new_n750), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n670), .A2(new_n729), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n727), .A2(new_n659), .A3(new_n687), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT115), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n648), .A2(new_n658), .B1(new_n684), .B2(new_n686), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n727), .A4(new_n774), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n775), .A2(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n628), .A2(new_n629), .A3(new_n652), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n527), .A2(KEYINPUT110), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n523), .A2(new_n786), .A3(new_n525), .A4(new_n526), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n789), .A3(new_n730), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n648), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n648), .A2(new_n791), .A3(KEYINPUT113), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n724), .A2(new_n726), .A3(new_n731), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n738), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n736), .A3(new_n800), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n606), .A2(new_n615), .B1(new_n598), .B2(new_n643), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n788), .B2(new_n740), .ZN(new_n804));
  AOI211_X1 g618(.A(KEYINPUT111), .B(new_n493), .C1(new_n785), .C2(new_n787), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n607), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n606), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n716), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n684), .A2(new_n706), .B1(new_n371), .B2(new_n599), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n697), .B(new_n371), .C1(new_n699), .C2(new_n703), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n783), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n799), .B1(new_n795), .B2(new_n796), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n736), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n776), .A2(new_n780), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n818), .B2(new_n781), .ZN(new_n819));
  MUX2_X1   g633(.A(new_n813), .B(new_n819), .S(KEYINPUT53), .Z(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT54), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n819), .B2(KEYINPUT53), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n777), .B1(new_n776), .B2(new_n780), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n812), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(KEYINPUT117), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n812), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n823), .B(new_n824), .C1(KEYINPUT54), .C2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n690), .A2(new_n451), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n768), .B(new_n767), .C1(new_n374), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n742), .A2(new_n532), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n714), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n838), .A2(new_n747), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n697), .A2(new_n678), .A3(new_n677), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n840), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT50), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n697), .A2(new_n730), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n724), .A3(new_n839), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n670), .A2(new_n251), .A3(new_n532), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n740), .A3(new_n611), .A4(new_n610), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n841), .A2(new_n844), .A3(new_n846), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n614), .ZN(new_n854));
  INV_X1    g668(.A(new_n719), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n531), .C1(new_n855), .C2(new_n840), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT118), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n845), .A2(new_n371), .A3(new_n839), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT48), .Z(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(KEYINPUT118), .B2(new_n856), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n852), .A2(new_n853), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n836), .A2(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n837), .B(KEYINPUT49), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n741), .A2(new_n374), .A3(new_n678), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n602), .A3(new_n677), .A4(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n670), .B2(new_n865), .ZN(G75));
  NAND2_X1  g680(.A1(new_n581), .A2(new_n585), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n589), .A2(new_n591), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n592), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n833), .B1(new_n826), .B2(new_n831), .ZN(new_n872));
  INV_X1    g686(.A(G210), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n188), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT119), .B(new_n871), .C1(new_n874), .C2(KEYINPUT56), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n229), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n874), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n871), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT119), .B1(new_n874), .B2(KEYINPUT56), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(G51));
  NAND2_X1  g699(.A1(G469), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT57), .Z(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n832), .B2(new_n834), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT54), .B(new_n833), .C1(new_n826), .C2(new_n831), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(KEYINPUT120), .B(new_n887), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n449), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n872), .A2(new_n188), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(G469), .A3(new_n751), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n876), .B1(new_n895), .B2(new_n897), .ZN(G54));
  AND2_X1   g712(.A1(KEYINPUT58), .A2(G475), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n896), .A2(new_n487), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n487), .B1(new_n896), .B2(new_n899), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n876), .ZN(G60));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT59), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n609), .B1(new_n836), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n609), .B(new_n904), .C1(new_n889), .C2(new_n890), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n877), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(G63));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT121), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n835), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n245), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n835), .A2(new_n636), .A3(new_n911), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n877), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G66));
  NAND2_X1  g732(.A1(new_n811), .A2(new_n229), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n529), .B2(new_n544), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n868), .B1(G898), .B2(new_n229), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G69));
  XNOR2_X1  g739(.A(new_n341), .B(new_n482), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n681), .A2(new_n727), .A3(new_n778), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n804), .A2(new_n805), .A3(new_n614), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n371), .A2(new_n929), .A3(new_n664), .A4(new_n730), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n769), .A2(new_n758), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n926), .B1(new_n932), .B2(G953), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n229), .A2(G900), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n756), .A2(new_n371), .A3(new_n749), .A4(new_n771), .ZN(new_n935));
  AND4_X1   g749(.A1(new_n727), .A2(new_n935), .A3(new_n738), .A4(new_n778), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n769), .A2(new_n936), .A3(new_n758), .A4(new_n736), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n937), .B2(new_n229), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n926), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n938), .A2(new_n939), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(G900), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n944), .B(G953), .C1(new_n414), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n414), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n933), .B(new_n947), .C1(new_n942), .C2(new_n943), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(KEYINPUT124), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(KEYINPUT124), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT125), .B(new_n946), .C1(new_n949), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n365), .A2(new_n336), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n820), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n937), .B2(new_n811), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n364), .A2(new_n328), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n876), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n932), .A2(new_n814), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n957), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n328), .A3(new_n364), .A4(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(KEYINPUT127), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(G57));
endmodule


