//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G1gat), .B(G29gat), .Z(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G57gat), .B(G85gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G127gat), .A2(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n213));
  AND2_X1   g012(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n215));
  OAI21_X1  g014(.A(G134gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT68), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G120gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(G120gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n216), .A4(new_n211), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n219), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(G127gat), .A2(G134gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(new_n210), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G148gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(G141gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT76), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(G141gat), .ZN(new_n238));
  INV_X1    g037(.A(G141gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G148gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT76), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244));
  OR2_X1    g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT2), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT75), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n239), .A2(G148gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n236), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G155gat), .B(G162gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT2), .B1(new_n240), .B2(new_n238), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n255), .A2(KEYINPUT75), .A3(new_n252), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n247), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(new_n253), .A3(new_n248), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT75), .B1(new_n255), .B2(new_n252), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n259), .A2(new_n260), .B1(new_n246), .B2(new_n243), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n216), .B(new_n211), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n262), .A2(KEYINPUT68), .B1(new_n231), .B2(new_n232), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n263), .A3(new_n226), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n234), .B2(new_n257), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n261), .A2(new_n263), .A3(new_n274), .A4(new_n226), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n279), .B(new_n247), .C1(new_n254), .C2(new_n256), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n234), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n266), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n270), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n257), .A2(KEYINPUT3), .B1(new_n263), .B2(new_n226), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n267), .B1(new_n284), .B2(new_n280), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT78), .A3(new_n276), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n269), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n288));
  INV_X1    g087(.A(new_n234), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(new_n261), .A3(new_n272), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n264), .A2(new_n274), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n204), .B(new_n209), .C1(new_n287), .C2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n209), .B1(new_n287), .B2(new_n294), .ZN(new_n296));
  INV_X1    g095(.A(new_n269), .ZN(new_n297));
  AND4_X1   g096(.A1(KEYINPUT78), .A2(new_n276), .A3(new_n266), .A4(new_n281), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT78), .B1(new_n285), .B2(new_n276), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n209), .B1(new_n288), .B2(new_n292), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n204), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI211_X1 g103(.A(KEYINPUT81), .B(new_n204), .C1(new_n300), .C2(new_n301), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n307), .B1(new_n312), .B2(KEYINPUT22), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n308), .A2(G211gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n308), .A2(G211gat), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT74), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n311), .ZN(new_n322));
  OAI21_X1  g121(.A(G218gat), .B1(new_n322), .B2(new_n309), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n325), .A2(new_n307), .A3(new_n316), .A4(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G226gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT27), .B(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(KEYINPUT28), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT27), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(G190gat), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n333), .B1(new_n339), .B2(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(KEYINPUT26), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n340), .A2(new_n341), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(KEYINPUT24), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(G183gat), .A3(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT64), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n342), .B2(KEYINPUT23), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n342), .A2(KEYINPUT23), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .A4(new_n345), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n352), .A2(KEYINPUT64), .A3(new_n353), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT25), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n334), .A2(new_n335), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n332), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n366), .B2(new_n352), .ZN(new_n367));
  INV_X1    g166(.A(new_n360), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n348), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n330), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n346), .A2(new_n341), .A3(new_n347), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT66), .B(G183gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n337), .B1(new_n376), .B2(KEYINPUT27), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n377), .B2(G190gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n374), .B1(new_n378), .B2(new_n333), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n352), .A2(new_n353), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n368), .A2(new_n382), .A3(new_n362), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n364), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n384), .B2(new_n369), .ZN(new_n385));
  INV_X1    g184(.A(new_n330), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n327), .B1(new_n373), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n385), .B2(KEYINPUT29), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n327), .B1(new_n371), .B2(new_n330), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT30), .A4(new_n394), .ZN(new_n398));
  INV_X1    g197(.A(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n327), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n330), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n389), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n385), .B2(new_n386), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n373), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(new_n398), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n306), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G78gat), .B(G106gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n321), .A2(new_n372), .A3(new_n326), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n279), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n257), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n280), .A2(new_n372), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n327), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n417), .A2(new_n419), .A3(G228gat), .A4(G233gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n421), .B(KEYINPUT83), .Z(new_n422));
  AOI21_X1  g221(.A(new_n261), .B1(new_n415), .B2(new_n279), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n280), .A2(new_n372), .B1(new_n326), .B2(new_n321), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT84), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n414), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AND4_X1   g229(.A1(new_n414), .A2(new_n429), .A3(new_n420), .A4(new_n425), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n413), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n414), .A3(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(new_n429), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n420), .A2(new_n425), .ZN(new_n435));
  OAI21_X1  g234(.A(G22gat), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(new_n412), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n383), .A2(new_n364), .B1(new_n368), .B2(new_n367), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n289), .B1(new_n440), .B2(new_n379), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n348), .B(new_n234), .C1(new_n363), .C2(new_n370), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  AOI211_X1 g245(.A(KEYINPUT34), .B(new_n446), .C1(new_n441), .C2(new_n442), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT70), .B(G71gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(G99gat), .ZN(new_n450));
  XOR2_X1   g249(.A(G15gat), .B(G43gat), .Z(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n441), .A2(new_n446), .A3(new_n442), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n453), .B(KEYINPUT32), .C1(new_n454), .C2(new_n452), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n448), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT72), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n458), .ZN(new_n462));
  INV_X1    g261(.A(new_n448), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n448), .A2(new_n457), .A3(KEYINPUT72), .A4(new_n458), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n463), .B1(new_n462), .B2(KEYINPUT71), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT36), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n408), .A2(new_n438), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n403), .B2(new_n373), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n399), .B1(new_n475), .B2(new_n402), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n388), .B2(new_n391), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT37), .B1(new_n402), .B2(new_n404), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT37), .B1(new_n389), .B2(new_n390), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n388), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n394), .A2(KEYINPUT38), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n478), .A2(new_n295), .A3(new_n483), .A4(new_n395), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n300), .A2(new_n293), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT86), .B1(new_n485), .B2(new_n209), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  INV_X1    g286(.A(new_n209), .ZN(new_n488));
  AOI211_X1 g287(.A(new_n487), .B(new_n488), .C1(new_n300), .C2(new_n293), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n490), .B2(new_n302), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n296), .A2(new_n487), .ZN(new_n492));
  OAI211_X1 g291(.A(KEYINPUT86), .B(new_n209), .C1(new_n287), .C2(new_n294), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n281), .A2(new_n290), .A3(new_n291), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n267), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n258), .A2(new_n264), .A3(new_n266), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT39), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n494), .B2(new_n267), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT40), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n494), .A2(new_n267), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT39), .A3(new_n498), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n488), .A4(new_n496), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n492), .A2(new_n406), .A3(new_n493), .A4(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n432), .A2(new_n437), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n491), .A2(new_n509), .A3(KEYINPUT87), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n405), .A2(new_n398), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n512), .A2(new_n397), .B1(new_n501), .B2(new_n505), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n438), .B1(new_n490), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n302), .A3(new_n493), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n295), .A2(new_n483), .A3(new_n395), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n478), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n511), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n473), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT71), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n438), .A2(new_n520), .A3(new_n469), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n306), .A3(new_n407), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n523));
  NOR4_X1   g322(.A1(new_n466), .A2(new_n438), .A3(KEYINPUT35), .A4(new_n406), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n515), .A2(new_n295), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G197gat), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT11), .B(G169gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT12), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT88), .Z(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT95), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n539), .A2(new_n540), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n539), .B(KEYINPUT91), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n540), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(G29gat), .B2(G36gat), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n548), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(G1gat), .ZN(new_n556));
  INV_X1    g355(.A(G1gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT16), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT93), .ZN(new_n560));
  INV_X1    g359(.A(G8gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT94), .B(G8gat), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n554), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n546), .A2(new_n553), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT92), .B1(new_n570), .B2(KEYINPUT17), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n570), .B2(KEYINPUT17), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n569), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n536), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n572), .B1(new_n554), .B2(new_n573), .ZN(new_n580));
  AOI211_X1 g379(.A(KEYINPUT92), .B(KEYINPUT17), .C1(new_n546), .C2(new_n553), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n576), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n536), .A3(new_n578), .A4(new_n568), .ZN(new_n583));
  OR3_X1    g382(.A1(new_n554), .A2(new_n567), .A3(KEYINPUT96), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT96), .B1(new_n554), .B2(new_n567), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n568), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n578), .B(KEYINPUT13), .Z(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n534), .B1(new_n579), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n578), .A3(new_n568), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT95), .A3(new_n535), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n592), .A2(new_n533), .A3(new_n588), .A4(new_n583), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n202), .B1(new_n528), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  AOI211_X1 g395(.A(KEYINPUT97), .B(new_n596), .C1(new_n519), .C2(new_n527), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  AND2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(KEYINPUT9), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(KEYINPUT100), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(KEYINPUT100), .B2(new_n602), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n601), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n606), .B2(new_n601), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n567), .B1(new_n612), .B2(KEYINPUT21), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G127gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(G127gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  INV_X1    g420(.A(new_n613), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n617), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g424(.A(G155gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n620), .A2(new_n623), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT7), .ZN(new_n634));
  INV_X1    g433(.A(G85gat), .ZN(new_n635));
  OAI21_X1  g434(.A(G92gat), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G92gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n636), .A2(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT8), .ZN(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(KEYINPUT101), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(KEYINPUT101), .B2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G99gat), .B(G106gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI221_X1 g446(.A(new_n647), .B1(new_n573), .B2(new_n554), .C1(new_n580), .C2(new_n581), .ZN(new_n648));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT102), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n554), .A2(new_n646), .B1(KEYINPUT41), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n648), .B2(new_n653), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n655), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n648), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n650), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n663), .B2(new_n654), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n611), .A2(new_n647), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n606), .A2(new_n601), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n608), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n604), .A3(new_n646), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n668), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT10), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n669), .A2(new_n680), .A3(new_n673), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n672), .A2(KEYINPUT10), .A3(new_n604), .A4(new_n646), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n681), .A2(new_n682), .B1(G230gat), .B2(G233gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n667), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n668), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n674), .A2(new_n678), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n677), .B(KEYINPUT104), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n668), .B(KEYINPUT105), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n681), .B2(new_n682), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n692), .B2(new_n674), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n633), .A2(new_n666), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n598), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n306), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g499(.A1(new_n598), .A2(new_n407), .A3(new_n696), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n701), .A2(new_n702), .A3(new_n561), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n701), .B2(new_n561), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n701), .A2(new_n705), .A3(new_n706), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n703), .B(new_n704), .C1(new_n707), .C2(new_n708), .ZN(G1325gat));
  INV_X1    g508(.A(G15gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n466), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n697), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n468), .A2(new_n472), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n468), .B2(new_n472), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n598), .A2(new_n696), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n712), .B1(new_n717), .B2(new_n710), .ZN(G1326gat));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n697), .A2(new_n721), .A3(new_n438), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n697), .B2(new_n438), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n724), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n722), .A3(new_n719), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1327gat));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n528), .B2(new_n665), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n665), .A2(new_n729), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n508), .B1(new_n306), .B2(new_n407), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT87), .B1(new_n491), .B2(new_n509), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n514), .A2(new_n511), .A3(new_n517), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n716), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n731), .B1(new_n736), .B2(new_n527), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n633), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n695), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n596), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G29gat), .B1(new_n742), .B2(new_n306), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n522), .A2(KEYINPUT35), .B1(new_n524), .B2(new_n525), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n734), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n473), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT97), .B1(new_n746), .B2(new_n596), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n528), .A2(new_n202), .A3(new_n594), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n740), .A2(new_n666), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n306), .A2(G29gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n749), .A2(new_n755), .A3(new_n750), .A4(new_n751), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n753), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n743), .B1(new_n757), .B2(new_n758), .ZN(G1328gat));
  NAND2_X1  g558(.A1(new_n749), .A2(new_n750), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n406), .A2(new_n538), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G36gat), .B1(new_n742), .B2(new_n407), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT46), .B1(new_n760), .B2(new_n761), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(G1329gat));
  NAND2_X1  g564(.A1(new_n468), .A2(new_n472), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n468), .A2(new_n472), .A3(new_n713), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(new_n741), .C1(new_n730), .C2(new_n737), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G43gat), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n740), .A2(G43gat), .A3(new_n466), .A4(new_n666), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n595), .B2(new_n597), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n749), .A2(KEYINPUT110), .A3(new_n772), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n771), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n774), .B1(new_n781), .B2(new_n782), .ZN(G1330gat));
  OAI211_X1 g582(.A(new_n438), .B(new_n741), .C1(new_n730), .C2(new_n737), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G50gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n508), .A2(G50gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n749), .A2(new_n750), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n788), .B(new_n791), .ZN(G1331gat));
  AOI21_X1  g591(.A(new_n744), .B1(new_n735), .B2(new_n716), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n633), .A2(new_n666), .A3(new_n694), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n594), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n698), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n406), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT49), .B(G64gat), .Z(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(G1333gat));
  NAND2_X1  g600(.A1(new_n795), .A2(new_n769), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n466), .A2(G71gat), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n802), .A2(G71gat), .B1(new_n795), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n795), .A2(new_n438), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g606(.A1(new_n739), .A2(new_n596), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n695), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n738), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810), .B2(new_n306), .ZN(new_n811));
  INV_X1    g610(.A(new_n732), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n510), .B2(new_n518), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n527), .B1(new_n813), .B2(new_n769), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n739), .A2(new_n596), .A3(new_n665), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(KEYINPUT51), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n793), .B2(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n698), .A2(new_n635), .A3(new_n694), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n811), .B1(new_n821), .B2(new_n822), .ZN(G1336gat));
  OAI21_X1  g622(.A(G92gat), .B1(new_n810), .B2(new_n407), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n695), .A2(G92gat), .A3(new_n407), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n820), .A2(new_n827), .B1(new_n825), .B2(KEYINPUT52), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n824), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n810), .B2(new_n716), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n695), .A2(new_n466), .A3(G99gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n821), .B2(new_n833), .ZN(G1338gat));
  OAI211_X1 g633(.A(new_n438), .B(new_n809), .C1(new_n730), .C2(new_n737), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G106gat), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n695), .A2(new_n508), .A3(G106gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(KEYINPUT115), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n836), .A2(KEYINPUT114), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n835), .A2(G106gat), .B1(new_n820), .B2(new_n837), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT114), .B1(new_n845), .B2(KEYINPUT115), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n842), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(G1339gat));
  NAND3_X1  g647(.A1(new_n681), .A2(new_n682), .A3(new_n691), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n686), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n677), .B1(new_n692), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n850), .A2(new_n852), .A3(new_n853), .A4(KEYINPUT55), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n689), .ZN(new_n855));
  INV_X1    g654(.A(new_n691), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n685), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n857), .B(new_n678), .C1(new_n858), .C2(new_n683), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n855), .A2(new_n594), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT117), .B1(new_n577), .B2(new_n578), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n586), .A2(new_n587), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n577), .A2(KEYINPUT117), .A3(new_n578), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n532), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n593), .A3(new_n694), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n665), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n665), .A2(new_n869), .A3(new_n593), .A4(new_n861), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n863), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n739), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n633), .A2(new_n596), .A3(new_n666), .A4(new_n695), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n306), .A2(new_n406), .A3(new_n466), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n508), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n220), .A3(new_n596), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n306), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n521), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n407), .A3(new_n594), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(new_n220), .ZN(G1340gat));
  INV_X1    g685(.A(G120gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n879), .A2(new_n887), .A3(new_n695), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n884), .A2(new_n407), .A3(new_n694), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n887), .ZN(G1341gat));
  OAI22_X1  g689(.A1(new_n879), .A2(new_n739), .B1(new_n215), .B2(new_n214), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n884), .A2(new_n407), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n739), .A2(new_n215), .A3(new_n214), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(G1342gat));
  NOR2_X1   g693(.A1(new_n666), .A2(G134gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n884), .A2(new_n407), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  OAI21_X1  g696(.A(G134gat), .B1(new_n879), .B2(new_n666), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n769), .A2(new_n508), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n881), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n594), .A2(new_n239), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n902), .A2(new_n406), .A3(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n769), .A2(new_n306), .A3(new_n406), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n874), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n850), .A2(new_n852), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n860), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n855), .A2(new_n911), .A3(new_n594), .A4(new_n863), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n870), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n666), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n912), .B2(new_n870), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n739), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n876), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n508), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n877), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n923), .B2(new_n508), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n906), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n594), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n904), .B1(new_n926), .B2(G141gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n406), .B1(new_n902), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n929), .B2(new_n902), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n903), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n239), .B1(new_n925), .B2(new_n594), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n927), .A2(new_n928), .B1(new_n932), .B2(new_n933), .ZN(G1344gat));
  OAI21_X1  g733(.A(KEYINPUT59), .B1(new_n931), .B2(new_n695), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n235), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n922), .A2(new_n924), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n905), .A2(new_n694), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n937), .A2(KEYINPUT59), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n919), .B2(new_n438), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n877), .A2(new_n921), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(KEYINPUT59), .B(G148gat), .C1(new_n943), .C2(new_n938), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n936), .A2(new_n939), .A3(new_n944), .ZN(G1345gat));
  OR2_X1    g744(.A1(new_n931), .A2(new_n739), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n633), .A2(G155gat), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT122), .Z(new_n948));
  AOI22_X1  g747(.A1(new_n946), .A2(new_n626), .B1(new_n925), .B2(new_n948), .ZN(G1346gat));
  NAND2_X1  g748(.A1(new_n925), .A2(new_n665), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G162gat), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n666), .A2(G162gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n931), .B2(new_n952), .ZN(G1347gat));
  AOI21_X1  g752(.A(new_n698), .B1(new_n875), .B2(new_n876), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n521), .A2(new_n406), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT123), .Z(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n594), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n306), .A2(new_n406), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n466), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n877), .A2(new_n508), .A3(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n877), .A2(KEYINPUT124), .A3(new_n508), .A4(new_n961), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n594), .A2(G169gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n959), .B1(new_n966), .B2(new_n967), .ZN(G1348gat));
  INV_X1    g767(.A(G176gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n958), .A2(new_n969), .A3(new_n694), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n966), .A2(new_n694), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n969), .ZN(G1349gat));
  AOI21_X1  g771(.A(new_n365), .B1(new_n966), .B2(new_n633), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n958), .A2(new_n331), .A3(new_n633), .ZN(new_n974));
  OR3_X1    g773(.A1(new_n973), .A2(KEYINPUT60), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT60), .B1(new_n973), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n964), .A2(new_n665), .A3(new_n965), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G190gat), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n978), .A2(new_n981), .A3(G190gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(KEYINPUT61), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n958), .A2(new_n332), .A3(new_n665), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n983), .B(new_n984), .C1(KEYINPUT61), .C2(new_n980), .ZN(G1351gat));
  NOR3_X1   g784(.A1(new_n769), .A2(new_n407), .A3(new_n508), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n877), .A2(new_n306), .A3(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n594), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n769), .A2(new_n960), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n876), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n992), .B1(new_n917), .B2(new_n739), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n920), .B1(new_n993), .B2(new_n508), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n991), .B1(new_n994), .B2(new_n941), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n594), .A2(G197gat), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(G1352gat));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  INV_X1    g797(.A(G204gat), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n999), .B1(new_n995), .B2(new_n694), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n695), .A2(G204gat), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT126), .B1(new_n987), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n954), .A2(new_n1004), .A3(new_n986), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1003), .A2(KEYINPUT62), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n998), .B1(new_n1000), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n694), .B(new_n990), .C1(new_n940), .C2(new_n942), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(G204gat), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1003), .A2(KEYINPUT62), .A3(new_n1005), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT62), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1013), .A2(KEYINPUT127), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1011), .A2(new_n1017), .ZN(G1353gat));
  NAND4_X1  g817(.A1(new_n988), .A2(new_n310), .A3(new_n311), .A4(new_n633), .ZN(new_n1019));
  OAI211_X1 g818(.A(new_n633), .B(new_n990), .C1(new_n940), .C2(new_n942), .ZN(new_n1020));
  AND3_X1   g819(.A1(new_n1020), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1021));
  AOI21_X1  g820(.A(KEYINPUT63), .B1(new_n1020), .B2(G211gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(G1354gat));
  NAND3_X1  g822(.A1(new_n988), .A2(new_n308), .A3(new_n665), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n995), .A2(new_n665), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1024), .B1(new_n1025), .B2(new_n308), .ZN(G1355gat));
endmodule


